// application_selector.v


`timescale 1 ps / 1 ps
module application_selector (
		output wire        local_wdata_req_from_the_ddr2_sdram,          //            ddr2_sdram_external_connection.local_wdata_req
		output wire        local_init_done_from_the_ddr2_sdram,          //                                          .local_init_done
		output wire        local_refresh_ack_from_the_ddr2_sdram,        //                                          .local_refresh_ack
		output wire        reset_phy_clk_n_from_the_ddr2_sdram,          //                                          .reset_phy_clk_n
		output wire        MOSI_from_the_touch_panel_spi,                //                  touch_panel_spi_external.MOSI
		input  wire        MISO_to_the_touch_panel_spi,                  //                                          .MISO
		output wire        SCLK_from_the_touch_panel_spi,                //                                          .SCLK
		output wire        SS_n_from_the_touch_panel_spi,                //                                          .SS_n
		output wire        out_port_from_the_lcd_i2c_en,                 //            lcd_i2c_en_external_connection.export
		output wire        local_wdata_req_from_the_ddr2_sdram_1,        //          ddr2_sdram_1_external_connection.local_wdata_req
		output wire        local_refresh_ack_from_the_ddr2_sdram_1,      //                                          .local_refresh_ack
		output wire        reset_phy_clk_n_from_the_ddr2_sdram_1,        //                                          .reset_phy_clk_n
		output wire        local_init_done_from_the_ddr2_sdram_1,        //                                          .local_init_done
		output wire        pll_c2_out,                                   //                                c2_out_clk.clk
		input  wire        reset_n,                                      //                    merged_resets_in_reset.reset_n
		inout  wire        bidir_port_to_and_from_the_lcd_i2c_sdat,      //          lcd_i2c_sdat_external_connection.export
		output wire        HD_from_the_lcd_sync_generator,               //                   lcd_sync_generator_sync.HD
		output wire [7:0]  RGB_OUT_from_the_lcd_sync_generator,          //                                          .RGB_OUT
		output wire        VD_from_the_lcd_sync_generator,               //                                          .VD
		output wire        DEN_from_the_lcd_sync_generator,              //                                          .DEN
		output wire        ddr2_sdram_1_phy_clk_out,                     //                        sysclk_001_out_clk.clk
		output wire        pll_c0_out,                                   //                                c0_out_clk.clk
		input  wire        in_port_to_the_touch_panel_pen_irq_n,         // touch_panel_pen_irq_n_external_connection.export
		input  wire        ddr2_sdram_reset_n,                           //                 ddr2_sdram_global_reset_n.reset_n
		output wire        ddr2_sdram_phy_clk_out,                       //                            sysclk_out_clk.clk
		output wire        ddr2_sdram_aux_half_rate_clk_out,             //                        ddr2_sdram_auxhalf.clk
		input  wire        clk,                                          //                                clk_clk_in.clk
		output wire        mdio_out_from_the_tse_mac,                    //                tse_mac_conduit_connection.mdio_out
		output wire        ena_10_from_the_tse_mac,                      //                                          .ena_10
		input  wire        rx_clk_to_the_tse_mac,                        //                                          .rx_clk
		output wire        mdio_oen_from_the_tse_mac,                    //                                          .mdio_oen
		input  wire        set_1000_to_the_tse_mac,                      //                                          .set_1000
		output wire        gm_tx_err_from_the_tse_mac,                   //                                          .gm_tx_err
		output wire [3:0]  m_tx_d_from_the_tse_mac,                      //                                          .m_tx_d
		output wire        eth_mode_from_the_tse_mac,                    //                                          .eth_mode
		input  wire        m_rx_en_to_the_tse_mac,                       //                                          .m_rx_en
		input  wire [7:0]  gm_rx_d_to_the_tse_mac,                       //                                          .gm_rx_d
		input  wire        m_rx_col_to_the_tse_mac,                      //                                          .m_rx_col
		output wire [7:0]  gm_tx_d_from_the_tse_mac,                     //                                          .gm_tx_d
		input  wire        tx_clk_to_the_tse_mac,                        //                                          .tx_clk
		output wire        m_tx_en_from_the_tse_mac,                     //                                          .m_tx_en
		output wire        gm_tx_en_from_the_tse_mac,                    //                                          .gm_tx_en
		input  wire        set_10_to_the_tse_mac,                        //                                          .set_10
		input  wire        gm_rx_err_to_the_tse_mac,                     //                                          .gm_rx_err
		input  wire        mdio_in_to_the_tse_mac,                       //                                          .mdio_in
		input  wire        gm_rx_dv_to_the_tse_mac,                      //                                          .gm_rx_dv
		output wire        m_tx_err_from_the_tse_mac,                    //                                          .m_tx_err
		input  wire        m_rx_crs_to_the_tse_mac,                      //                                          .m_rx_crs
		output wire        mdc_from_the_tse_mac,                         //                                          .mdc
		input  wire [3:0]  m_rx_d_to_the_tse_mac,                        //                                          .m_rx_d
		input  wire        m_rx_err_to_the_tse_mac,                      //                                          .m_rx_err
		input  wire        rxd_to_the_uart1,                             //                 uart1_external_connection.rxd
		output wire        txd_from_the_uart1,                           //                                          .txd
		output wire        out_port_from_the_lcd_i2c_scl,                //           lcd_i2c_scl_external_connection.export
		input  wire        ddr2_sdram_1_reset_n,                         //               ddr2_sdram_1_global_reset_n.reset_n
		output wire        ddr2_sdram_aux_full_rate_clk_out,             //                        ddr2_sdram_auxfull.clk
		output wire        mem_odt_from_the_ddr2_sdram,                  //                         ddr2_sdram_memory.mem_odt
		output wire        mem_cas_n_from_the_ddr2_sdram,                //                                          .mem_cas_n
		inout  wire [1:0]  mem_dqs_to_and_from_the_ddr2_sdram,           //                                          .mem_dqs
		output wire        mem_cs_n_from_the_ddr2_sdram,                 //                                          .mem_cs_n
		output wire        mem_we_n_from_the_ddr2_sdram,                 //                                          .mem_we_n
		output wire [1:0]  mem_ba_from_the_ddr2_sdram,                   //                                          .mem_ba
		inout  wire        mem_clk_to_and_from_the_ddr2_sdram,           //                                          .mem_clk
		output wire        mem_cke_from_the_ddr2_sdram,                  //                                          .mem_cke
		inout  wire        mem_clk_n_to_and_from_the_ddr2_sdram,         //                                          .mem_clk_n
		output wire        mem_ras_n_from_the_ddr2_sdram,                //                                          .mem_ras_n
		output wire [1:0]  mem_dm_from_the_ddr2_sdram,                   //                                          .mem_dm
		output wire [12:0] mem_addr_from_the_ddr2_sdram,                 //                                          .mem_addr
		inout  wire [15:0] mem_dq_to_and_from_the_ddr2_sdram,            //                                          .mem_dq
		inout  wire        bidir_port_to_and_from_the_pio_id_eeprom_dat, //     pio_id_eeprom_dat_external_connection.export
		inout  wire [31:0] flash_tristate_bridge_data,                   //        flash_tristate_bridge_bridge_0_out.flash_tristate_bridge_data
		inout  wire        we_n_to_the_max2,                             //                                          .we_n_to_the_max2
		inout  wire        read_n_to_the_ext_flash,                      //                                          .read_n_to_the_ext_flash
		inout  wire [25:0] flash_tristate_bridge_address,                //                                          .flash_tristate_bridge_address
		inout  wire        cs_n_to_the_max2,                             //                                          .cs_n_to_the_max2
		inout  wire        oe_n_to_the_max2,                             //                                          .oe_n_to_the_max2
		inout  wire        select_n_to_the_ext_flash,                    //                                          .select_n_to_the_ext_flash
		inout  wire        write_n_to_the_ext_flash,                     //                                          .write_n_to_the_ext_flash
		output wire        mem_cke_from_the_ddr2_sdram_1,                //                       ddr2_sdram_1_memory.mem_cke
		inout  wire        mem_clk_to_and_from_the_ddr2_sdram_1,         //                                          .mem_clk
		inout  wire [15:0] mem_dq_to_and_from_the_ddr2_sdram_1,          //                                          .mem_dq
		output wire        mem_cas_n_from_the_ddr2_sdram_1,              //                                          .mem_cas_n
		inout  wire        mem_clk_n_to_and_from_the_ddr2_sdram_1,       //                                          .mem_clk_n
		output wire        mem_cs_n_from_the_ddr2_sdram_1,               //                                          .mem_cs_n
		output wire [12:0] mem_addr_from_the_ddr2_sdram_1,               //                                          .mem_addr
		output wire        mem_ras_n_from_the_ddr2_sdram_1,              //                                          .mem_ras_n
		output wire [1:0]  mem_dm_from_the_ddr2_sdram_1,                 //                                          .mem_dm
		output wire        mem_we_n_from_the_ddr2_sdram_1,               //                                          .mem_we_n
		inout  wire [1:0]  mem_dqs_to_and_from_the_ddr2_sdram_1,         //                                          .mem_dqs
		output wire [1:0]  mem_ba_from_the_ddr2_sdram_1,                 //                                          .mem_ba
		output wire        mem_odt_from_the_ddr2_sdram_1,                //                                          .mem_odt
		output wire [7:0]  out_port_from_the_led_pio,                    //               led_pio_external_connection.export
		input  wire [3:0]  in_port_to_the_button_pio,                    //            button_pio_external_connection.export
		input  wire        clk_125,                                      //                            clk_125_clk_in.clk
		output wire        ddr2_sdram_1_aux_full_rate_clk_out,           //                      ddr2_sdram_1_auxfull.clk
		inout  wire        SD_DAT2_to_and_from_the_sls_sdhc,             //                      sls_sdhc_conduit_end.DAT2
		inout  wire        SD_DAT3_to_and_from_the_sls_sdhc,             //                                          .DAT3
		output wire        SD_Busy_from_the_sls_sdhc,                    //                                          .Busy
		input  wire        SD_In_to_the_sls_sdhc,                        //                                          .In
		inout  wire        SD_DAT1_to_and_from_the_sls_sdhc,             //                                          .DAT1
		inout  wire        SD_CMD_to_and_from_the_sls_sdhc,              //                                          .CMD
		inout  wire        SD_DAT0_to_and_from_the_sls_sdhc,             //                                          .DAT0
		input  wire        SD_Wp_to_the_sls_sdhc,                        //                                          .Wp
		output wire        SD_CLK_from_the_sls_sdhc,                     //                                          .CLK
		output wire        out_port_from_the_pio_id_eeprom_scl,          //     pio_id_eeprom_scl_external_connection.export
		output wire        ddr2_sdram_1_aux_half_rate_clk_out            //                      ddr2_sdram_1_auxhalf.clk
	);

	wire          sgdma_tx_out_endofpacket;                                                                                       // sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	wire          sgdma_tx_out_valid;                                                                                             // sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	wire          sgdma_tx_out_startofpacket;                                                                                     // sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	wire          sgdma_tx_out_error;                                                                                             // sgdma_tx:out_error -> tse_mac:ff_tx_err
	wire    [1:0] sgdma_tx_out_empty;                                                                                             // sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	wire   [31:0] sgdma_tx_out_data;                                                                                              // sgdma_tx:out_data -> tse_mac:ff_tx_data
	wire          sgdma_tx_out_ready;                                                                                             // tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	wire          tse_mac_receive_endofpacket;                                                                                    // tse_mac:ff_rx_eop -> sgdma_rx:in_endofpacket
	wire          tse_mac_receive_valid;                                                                                          // tse_mac:ff_rx_dval -> sgdma_rx:in_valid
	wire          tse_mac_receive_startofpacket;                                                                                  // tse_mac:ff_rx_sop -> sgdma_rx:in_startofpacket
	wire    [5:0] tse_mac_receive_error;                                                                                          // tse_mac:rx_err -> sgdma_rx:in_error
	wire    [1:0] tse_mac_receive_empty;                                                                                          // tse_mac:ff_rx_mod -> sgdma_rx:in_empty
	wire   [31:0] tse_mac_receive_data;                                                                                           // tse_mac:ff_rx_data -> sgdma_rx:in_data
	wire          tse_mac_receive_ready;                                                                                          // sgdma_rx:in_ready -> tse_mac:ff_rx_rdy
	wire          lcd_32_to_8_bits_dfa_out_endofpacket;                                                                           // lcd_32_to_8_bits_dfa:out_endofpacket -> lcd_sync_generator:eop
	wire          lcd_32_to_8_bits_dfa_out_valid;                                                                                 // lcd_32_to_8_bits_dfa:out_valid -> lcd_sync_generator:valid
	wire          lcd_32_to_8_bits_dfa_out_startofpacket;                                                                         // lcd_32_to_8_bits_dfa:out_startofpacket -> lcd_sync_generator:sop
	wire          lcd_32_to_8_bits_dfa_out_empty;                                                                                 // lcd_32_to_8_bits_dfa:out_empty -> lcd_sync_generator:empty
	wire    [7:0] lcd_32_to_8_bits_dfa_out_data;                                                                                  // lcd_32_to_8_bits_dfa:out_data -> lcd_sync_generator:data
	wire          lcd_32_to_8_bits_dfa_out_ready;                                                                                 // lcd_sync_generator:ready -> lcd_32_to_8_bits_dfa:out_ready
	wire          lcd_64_to_32_bits_dfa_out_endofpacket;                                                                          // lcd_64_to_32_bits_dfa:out_endofpacket -> lcd_pixel_converter:eop_in
	wire          lcd_64_to_32_bits_dfa_out_valid;                                                                                // lcd_64_to_32_bits_dfa:out_valid -> lcd_pixel_converter:valid_in
	wire          lcd_64_to_32_bits_dfa_out_startofpacket;                                                                        // lcd_64_to_32_bits_dfa:out_startofpacket -> lcd_pixel_converter:sop_in
	wire    [1:0] lcd_64_to_32_bits_dfa_out_empty;                                                                                // lcd_64_to_32_bits_dfa:out_empty -> lcd_pixel_converter:empty_in
	wire   [31:0] lcd_64_to_32_bits_dfa_out_data;                                                                                 // lcd_64_to_32_bits_dfa:out_data -> lcd_pixel_converter:data_in
	wire          lcd_64_to_32_bits_dfa_out_ready;                                                                                // lcd_pixel_converter:ready_out -> lcd_64_to_32_bits_dfa:out_ready
	wire          lcd_pixel_converter_out_endofpacket;                                                                            // lcd_pixel_converter:eop_out -> lcd_32_to_8_bits_dfa:in_endofpacket
	wire          lcd_pixel_converter_out_valid;                                                                                  // lcd_pixel_converter:valid_out -> lcd_32_to_8_bits_dfa:in_valid
	wire          lcd_pixel_converter_out_startofpacket;                                                                          // lcd_pixel_converter:sop_out -> lcd_32_to_8_bits_dfa:in_startofpacket
	wire    [1:0] lcd_pixel_converter_out_empty;                                                                                  // lcd_pixel_converter:empty_out -> lcd_32_to_8_bits_dfa:in_empty
	wire   [23:0] lcd_pixel_converter_out_data;                                                                                   // lcd_pixel_converter:data_out -> lcd_32_to_8_bits_dfa:in_data
	wire          lcd_pixel_converter_out_ready;                                                                                  // lcd_32_to_8_bits_dfa:in_ready -> lcd_pixel_converter:ready_in
	wire          lcd_pixel_fifo_out_endofpacket;                                                                                 // lcd_pixel_fifo:avalonst_source_endofpacket -> lcd_ta_fifo_to_dfa:in_endofpacket
	wire          lcd_pixel_fifo_out_valid;                                                                                       // lcd_pixel_fifo:avalonst_source_valid -> lcd_ta_fifo_to_dfa:in_valid
	wire          lcd_pixel_fifo_out_startofpacket;                                                                               // lcd_pixel_fifo:avalonst_source_startofpacket -> lcd_ta_fifo_to_dfa:in_startofpacket
	wire    [2:0] lcd_pixel_fifo_out_empty;                                                                                       // lcd_pixel_fifo:avalonst_source_empty -> lcd_ta_fifo_to_dfa:in_empty
	wire   [63:0] lcd_pixel_fifo_out_data;                                                                                        // lcd_pixel_fifo:avalonst_source_data -> lcd_ta_fifo_to_dfa:in_data
	wire          lcd_pixel_fifo_out_ready;                                                                                       // lcd_ta_fifo_to_dfa:in_ready -> lcd_pixel_fifo:avalonst_source_ready
	wire          lcd_sgdma_out_endofpacket;                                                                                      // lcd_sgdma:out_endofpacket -> lcd_ta_sgdma_to_fifo:in_endofpacket
	wire          lcd_sgdma_out_valid;                                                                                            // lcd_sgdma:out_valid -> lcd_ta_sgdma_to_fifo:in_valid
	wire          lcd_sgdma_out_startofpacket;                                                                                    // lcd_sgdma:out_startofpacket -> lcd_ta_sgdma_to_fifo:in_startofpacket
	wire    [2:0] lcd_sgdma_out_empty;                                                                                            // lcd_sgdma:out_empty -> lcd_ta_sgdma_to_fifo:in_empty
	wire   [63:0] lcd_sgdma_out_data;                                                                                             // lcd_sgdma:out_data -> lcd_ta_sgdma_to_fifo:in_data
	wire          lcd_sgdma_out_ready;                                                                                            // lcd_ta_sgdma_to_fifo:in_ready -> lcd_sgdma:out_ready
	wire          lcd_ta_fifo_to_dfa_out_endofpacket;                                                                             // lcd_ta_fifo_to_dfa:out_endofpacket -> lcd_64_to_32_bits_dfa:in_endofpacket
	wire          lcd_ta_fifo_to_dfa_out_valid;                                                                                   // lcd_ta_fifo_to_dfa:out_valid -> lcd_64_to_32_bits_dfa:in_valid
	wire          lcd_ta_fifo_to_dfa_out_startofpacket;                                                                           // lcd_ta_fifo_to_dfa:out_startofpacket -> lcd_64_to_32_bits_dfa:in_startofpacket
	wire    [2:0] lcd_ta_fifo_to_dfa_out_empty;                                                                                   // lcd_ta_fifo_to_dfa:out_empty -> lcd_64_to_32_bits_dfa:in_empty
	wire   [63:0] lcd_ta_fifo_to_dfa_out_data;                                                                                    // lcd_ta_fifo_to_dfa:out_data -> lcd_64_to_32_bits_dfa:in_data
	wire          lcd_ta_fifo_to_dfa_out_ready;                                                                                   // lcd_64_to_32_bits_dfa:in_ready -> lcd_ta_fifo_to_dfa:out_ready
	wire          lcd_ta_sgdma_to_fifo_out_endofpacket;                                                                           // lcd_ta_sgdma_to_fifo:out_endofpacket -> lcd_pixel_fifo:avalonst_sink_endofpacket
	wire          lcd_ta_sgdma_to_fifo_out_valid;                                                                                 // lcd_ta_sgdma_to_fifo:out_valid -> lcd_pixel_fifo:avalonst_sink_valid
	wire          lcd_ta_sgdma_to_fifo_out_startofpacket;                                                                         // lcd_ta_sgdma_to_fifo:out_startofpacket -> lcd_pixel_fifo:avalonst_sink_startofpacket
	wire    [2:0] lcd_ta_sgdma_to_fifo_out_empty;                                                                                 // lcd_ta_sgdma_to_fifo:out_empty -> lcd_pixel_fifo:avalonst_sink_empty
	wire   [63:0] lcd_ta_sgdma_to_fifo_out_data;                                                                                  // lcd_ta_sgdma_to_fifo:out_data -> lcd_pixel_fifo:avalonst_sink_data
	wire          lcd_ta_sgdma_to_fifo_out_ready;                                                                                 // lcd_pixel_fifo:avalonst_sink_ready -> lcd_ta_sgdma_to_fifo:out_ready
	wire    [0:0] flash_tristate_bridge_pinsharer_0_tcm_cs_n_to_the_max2_out;                                                     // flash_tristate_bridge_pinSharer_0:cs_n_to_the_max2 -> flash_tristate_bridge_bridge_0:tcs_cs_n_to_the_max2
	wire    [0:0] flash_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out;                                            // flash_tristate_bridge_pinSharer_0:select_n_to_the_ext_flash -> flash_tristate_bridge_bridge_0:tcs_select_n_to_the_ext_flash
	wire          flash_tristate_bridge_pinsharer_0_tcm_grant;                                                                    // flash_tristate_bridge_bridge_0:grant -> flash_tristate_bridge_pinSharer_0:grant
	wire   [31:0] flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_out;                                           // flash_tristate_bridge_pinSharer_0:flash_tristate_bridge_data -> flash_tristate_bridge_bridge_0:tcs_flash_tristate_bridge_data
	wire          flash_tristate_bridge_pinsharer_0_tcm_request;                                                                  // flash_tristate_bridge_pinSharer_0:request -> flash_tristate_bridge_bridge_0:request
	wire    [0:0] flash_tristate_bridge_pinsharer_0_tcm_read_n_to_the_ext_flash_out;                                              // flash_tristate_bridge_pinSharer_0:read_n_to_the_ext_flash -> flash_tristate_bridge_bridge_0:tcs_read_n_to_the_ext_flash
	wire    [0:0] flash_tristate_bridge_pinsharer_0_tcm_we_n_to_the_max2_out;                                                     // flash_tristate_bridge_pinSharer_0:we_n_to_the_max2 -> flash_tristate_bridge_bridge_0:tcs_we_n_to_the_max2
	wire          flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_outen;                                         // flash_tristate_bridge_pinSharer_0:flash_tristate_bridge_data_outen -> flash_tristate_bridge_bridge_0:tcs_flash_tristate_bridge_data_outen
	wire    [0:0] flash_tristate_bridge_pinsharer_0_tcm_oe_n_to_the_max2_out;                                                     // flash_tristate_bridge_pinSharer_0:oe_n_to_the_max2 -> flash_tristate_bridge_bridge_0:tcs_oe_n_to_the_max2
	wire    [0:0] flash_tristate_bridge_pinsharer_0_tcm_write_n_to_the_ext_flash_out;                                             // flash_tristate_bridge_pinSharer_0:write_n_to_the_ext_flash -> flash_tristate_bridge_bridge_0:tcs_write_n_to_the_ext_flash
	wire   [31:0] flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_in;                                            // flash_tristate_bridge_bridge_0:tcs_flash_tristate_bridge_data_in -> flash_tristate_bridge_pinSharer_0:flash_tristate_bridge_data_in
	wire   [25:0] flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_address_out;                                        // flash_tristate_bridge_pinSharer_0:flash_tristate_bridge_address -> flash_tristate_bridge_bridge_0:tcs_flash_tristate_bridge_address
	wire          ext_flash_tcm_chipselect_n_out;                                                                                 // ext_flash:tcm_chipselect_n_out -> flash_tristate_bridge_pinSharer_0:tcs0_chipselect_n_out
	wire          ext_flash_tcm_grant;                                                                                            // flash_tristate_bridge_pinSharer_0:tcs0_grant -> ext_flash:tcm_grant
	wire          ext_flash_tcm_data_outen;                                                                                       // ext_flash:tcm_data_outen -> flash_tristate_bridge_pinSharer_0:tcs0_data_outen
	wire          ext_flash_tcm_request;                                                                                          // ext_flash:tcm_request -> flash_tristate_bridge_pinSharer_0:tcs0_request
	wire   [15:0] ext_flash_tcm_data_out;                                                                                         // ext_flash:tcm_data_out -> flash_tristate_bridge_pinSharer_0:tcs0_data_out
	wire          ext_flash_tcm_write_n_out;                                                                                      // ext_flash:tcm_write_n_out -> flash_tristate_bridge_pinSharer_0:tcs0_write_n_out
	wire   [25:0] ext_flash_tcm_address_out;                                                                                      // ext_flash:tcm_address_out -> flash_tristate_bridge_pinSharer_0:tcs0_address_out
	wire   [15:0] ext_flash_tcm_data_in;                                                                                          // flash_tristate_bridge_pinSharer_0:tcs0_data_in -> ext_flash:tcm_data_in
	wire          ext_flash_tcm_read_n_out;                                                                                       // ext_flash:tcm_read_n_out -> flash_tristate_bridge_pinSharer_0:tcs0_read_n_out
	wire          max2_tcm_chipselect_n_out;                                                                                      // max2:tcm_chipselect_n_out -> flash_tristate_bridge_pinSharer_0:tcs1_chipselect_n_out
	wire          max2_tcm_grant;                                                                                                 // flash_tristate_bridge_pinSharer_0:tcs1_grant -> max2:tcm_grant
	wire          max2_tcm_data_outen;                                                                                            // max2:tcm_data_outen -> flash_tristate_bridge_pinSharer_0:tcs1_data_outen
	wire          max2_tcm_request;                                                                                               // max2:tcm_request -> flash_tristate_bridge_pinSharer_0:tcs1_request
	wire   [31:0] max2_tcm_data_out;                                                                                              // max2:tcm_data_out -> flash_tristate_bridge_pinSharer_0:tcs1_data_out
	wire          max2_tcm_write_n_out;                                                                                           // max2:tcm_write_n_out -> flash_tristate_bridge_pinSharer_0:tcs1_write_n_out
	wire    [4:0] max2_tcm_address_out;                                                                                           // max2:tcm_address_out -> flash_tristate_bridge_pinSharer_0:tcs1_address_out
	wire   [31:0] max2_tcm_data_in;                                                                                               // flash_tristate_bridge_pinSharer_0:tcs1_data_in -> max2:tcm_data_in
	wire          max2_tcm_read_n_out;                                                                                            // max2:tcm_read_n_out -> flash_tristate_bridge_pinSharer_0:tcs1_read_n_out
	wire          cpu_data_master_waitrequest;                                                                                    // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                                      // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire   [28:0] cpu_data_master_address;                                                                                        // cpu:d_address -> cpu_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                                          // cpu:d_write -> cpu_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                                           // cpu:d_read -> cpu_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                                       // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                                                                    // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire          cpu_data_master_readdatavalid;                                                                                  // cpu_data_master_translator:av_readdatavalid -> cpu:d_readdatavalid
	wire    [3:0] cpu_data_master_byteenable;                                                                                     // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire          cpu_instruction_master_waitrequest;                                                                             // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire   [28:0] cpu_instruction_master_address;                                                                                 // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                                    // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                                // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_readdatavalid;                                                                           // cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	wire          sgdma_rx_descriptor_read_waitrequest;                                                                           // sgdma_rx_descriptor_read_translator:av_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire   [31:0] sgdma_rx_descriptor_read_address;                                                                               // sgdma_rx:descriptor_read_address -> sgdma_rx_descriptor_read_translator:av_address
	wire          sgdma_rx_descriptor_read_read;                                                                                  // sgdma_rx:descriptor_read_read -> sgdma_rx_descriptor_read_translator:av_read
	wire   [31:0] sgdma_rx_descriptor_read_readdata;                                                                              // sgdma_rx_descriptor_read_translator:av_readdata -> sgdma_rx:descriptor_read_readdata
	wire          sgdma_rx_descriptor_read_readdatavalid;                                                                         // sgdma_rx_descriptor_read_translator:av_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire          sgdma_rx_descriptor_write_waitrequest;                                                                          // sgdma_rx_descriptor_write_translator:av_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire   [31:0] sgdma_rx_descriptor_write_writedata;                                                                            // sgdma_rx:descriptor_write_writedata -> sgdma_rx_descriptor_write_translator:av_writedata
	wire   [31:0] sgdma_rx_descriptor_write_address;                                                                              // sgdma_rx:descriptor_write_address -> sgdma_rx_descriptor_write_translator:av_address
	wire          sgdma_rx_descriptor_write_write;                                                                                // sgdma_rx:descriptor_write_write -> sgdma_rx_descriptor_write_translator:av_write
	wire          sgdma_tx_descriptor_read_waitrequest;                                                                           // sgdma_tx_descriptor_read_translator:av_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire   [31:0] sgdma_tx_descriptor_read_address;                                                                               // sgdma_tx:descriptor_read_address -> sgdma_tx_descriptor_read_translator:av_address
	wire          sgdma_tx_descriptor_read_read;                                                                                  // sgdma_tx:descriptor_read_read -> sgdma_tx_descriptor_read_translator:av_read
	wire   [31:0] sgdma_tx_descriptor_read_readdata;                                                                              // sgdma_tx_descriptor_read_translator:av_readdata -> sgdma_tx:descriptor_read_readdata
	wire          sgdma_tx_descriptor_read_readdatavalid;                                                                         // sgdma_tx_descriptor_read_translator:av_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire          sgdma_tx_descriptor_write_waitrequest;                                                                          // sgdma_tx_descriptor_write_translator:av_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire   [31:0] sgdma_tx_descriptor_write_writedata;                                                                            // sgdma_tx:descriptor_write_writedata -> sgdma_tx_descriptor_write_translator:av_writedata
	wire   [31:0] sgdma_tx_descriptor_write_address;                                                                              // sgdma_tx:descriptor_write_address -> sgdma_tx_descriptor_write_translator:av_address
	wire          sgdma_tx_descriptor_write_write;                                                                                // sgdma_tx:descriptor_write_write -> sgdma_tx_descriptor_write_translator:av_write
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                                 // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                                   // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                                // cpu_jtag_debug_module_translator:av_chipselect -> cpu:jtag_debug_module_select
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                     // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                                  // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                             // cpu_jtag_debug_module_translator:av_begintransfer -> cpu:jtag_debug_module_begintransfer
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                               // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                                // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire   [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_writedata;                                                  // descriptor_memory_s1_translator:av_writedata -> descriptor_memory:writedata
	wire    [9:0] descriptor_memory_s1_translator_avalon_anti_slave_0_address;                                                    // descriptor_memory_s1_translator:av_address -> descriptor_memory:address
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect;                                                 // descriptor_memory_s1_translator:av_chipselect -> descriptor_memory:chipselect
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_clken;                                                      // descriptor_memory_s1_translator:av_clken -> descriptor_memory:clken
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_write;                                                      // descriptor_memory_s1_translator:av_write -> descriptor_memory:write
	wire   [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_readdata;                                                   // descriptor_memory:readdata -> descriptor_memory_s1_translator:av_readdata
	wire    [3:0] descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable;                                                 // descriptor_memory_s1_translator:av_byteenable -> descriptor_memory:byteenable
	wire   [31:0] sgdma_rx_csr_translator_avalon_anti_slave_0_writedata;                                                          // sgdma_rx_csr_translator:av_writedata -> sgdma_rx:csr_writedata
	wire    [3:0] sgdma_rx_csr_translator_avalon_anti_slave_0_address;                                                            // sgdma_rx_csr_translator:av_address -> sgdma_rx:csr_address
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect;                                                         // sgdma_rx_csr_translator:av_chipselect -> sgdma_rx:csr_chipselect
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_write;                                                              // sgdma_rx_csr_translator:av_write -> sgdma_rx:csr_write
	wire          sgdma_rx_csr_translator_avalon_anti_slave_0_read;                                                               // sgdma_rx_csr_translator:av_read -> sgdma_rx:csr_read
	wire   [31:0] sgdma_rx_csr_translator_avalon_anti_slave_0_readdata;                                                           // sgdma_rx:csr_readdata -> sgdma_rx_csr_translator:av_readdata
	wire   [31:0] sgdma_tx_csr_translator_avalon_anti_slave_0_writedata;                                                          // sgdma_tx_csr_translator:av_writedata -> sgdma_tx:csr_writedata
	wire    [3:0] sgdma_tx_csr_translator_avalon_anti_slave_0_address;                                                            // sgdma_tx_csr_translator:av_address -> sgdma_tx:csr_address
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect;                                                         // sgdma_tx_csr_translator:av_chipselect -> sgdma_tx:csr_chipselect
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_write;                                                              // sgdma_tx_csr_translator:av_write -> sgdma_tx:csr_write
	wire          sgdma_tx_csr_translator_avalon_anti_slave_0_read;                                                               // sgdma_tx_csr_translator:av_read -> sgdma_tx:csr_read
	wire   [31:0] sgdma_tx_csr_translator_avalon_anti_slave_0_readdata;                                                           // sgdma_tx:csr_readdata -> sgdma_tx_csr_translator:av_readdata
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest;                                                // tse_mac:waitrequest -> tse_mac_control_port_translator:av_waitrequest
	wire   [31:0] tse_mac_control_port_translator_avalon_anti_slave_0_writedata;                                                  // tse_mac_control_port_translator:av_writedata -> tse_mac:writedata
	wire    [7:0] tse_mac_control_port_translator_avalon_anti_slave_0_address;                                                    // tse_mac_control_port_translator:av_address -> tse_mac:address
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_write;                                                      // tse_mac_control_port_translator:av_write -> tse_mac:write
	wire          tse_mac_control_port_translator_avalon_anti_slave_0_read;                                                       // tse_mac_control_port_translator:av_read -> tse_mac:read
	wire   [31:0] tse_mac_control_port_translator_avalon_anti_slave_0_readdata;                                                   // tse_mac:readdata -> tse_mac_control_port_translator:av_readdata
	wire          sls_sdhc_control_translator_avalon_anti_slave_0_waitrequest;                                                    // sls_sdhc:AvS_waitrequest -> sls_sdhc_control_translator:av_waitrequest
	wire   [31:0] sls_sdhc_control_translator_avalon_anti_slave_0_writedata;                                                      // sls_sdhc_control_translator:av_writedata -> sls_sdhc:AvS_writedata
	wire    [4:0] sls_sdhc_control_translator_avalon_anti_slave_0_address;                                                        // sls_sdhc_control_translator:av_address -> sls_sdhc:AvS_address
	wire          sls_sdhc_control_translator_avalon_anti_slave_0_chipselect;                                                     // sls_sdhc_control_translator:av_chipselect -> sls_sdhc:AvS_chipselect
	wire          sls_sdhc_control_translator_avalon_anti_slave_0_write;                                                          // sls_sdhc_control_translator:av_write -> sls_sdhc:AvS_write_n
	wire          sls_sdhc_control_translator_avalon_anti_slave_0_read;                                                           // sls_sdhc_control_translator:av_read -> sls_sdhc:AvS_read_n
	wire   [31:0] sls_sdhc_control_translator_avalon_anti_slave_0_readdata;                                                       // sls_sdhc:AvS_readdata -> sls_sdhc_control_translator:av_readdata
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                           // pipeline_bridge_before_tristate_bridge:s0_waitrequest -> pipeline_bridge_before_tristate_bridge_s0_translator:av_waitrequest
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_burstcount;                            // pipeline_bridge_before_tristate_bridge_s0_translator:av_burstcount -> pipeline_bridge_before_tristate_bridge:s0_burstcount
	wire   [31:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_writedata;                             // pipeline_bridge_before_tristate_bridge_s0_translator:av_writedata -> pipeline_bridge_before_tristate_bridge:s0_writedata
	wire   [26:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_address;                               // pipeline_bridge_before_tristate_bridge_s0_translator:av_address -> pipeline_bridge_before_tristate_bridge:s0_address
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_write;                                 // pipeline_bridge_before_tristate_bridge_s0_translator:av_write -> pipeline_bridge_before_tristate_bridge:s0_write
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_read;                                  // pipeline_bridge_before_tristate_bridge_s0_translator:av_read -> pipeline_bridge_before_tristate_bridge:s0_read
	wire   [31:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_readdata;                              // pipeline_bridge_before_tristate_bridge:s0_readdata -> pipeline_bridge_before_tristate_bridge_s0_translator:av_readdata
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                           // pipeline_bridge_before_tristate_bridge_s0_translator:av_debugaccess -> pipeline_bridge_before_tristate_bridge:s0_debugaccess
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                         // pipeline_bridge_before_tristate_bridge:s0_readdatavalid -> pipeline_bridge_before_tristate_bridge_s0_translator:av_readdatavalid
	wire    [3:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_byteenable;                            // pipeline_bridge_before_tristate_bridge_s0_translator:av_byteenable -> pipeline_bridge_before_tristate_bridge:s0_byteenable
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                             // cpu_ddr_clock_bridge:s0_waitrequest -> cpu_ddr_clock_bridge_s0_translator:av_waitrequest
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                              // cpu_ddr_clock_bridge_s0_translator:av_burstcount -> cpu_ddr_clock_bridge:s0_burstcount
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata;                                               // cpu_ddr_clock_bridge_s0_translator:av_writedata -> cpu_ddr_clock_bridge:s0_writedata
	wire   [26:0] cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address;                                                 // cpu_ddr_clock_bridge_s0_translator:av_address -> cpu_ddr_clock_bridge:s0_address
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write;                                                   // cpu_ddr_clock_bridge_s0_translator:av_write -> cpu_ddr_clock_bridge:s0_write
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read;                                                    // cpu_ddr_clock_bridge_s0_translator:av_read -> cpu_ddr_clock_bridge:s0_read
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata;                                                // cpu_ddr_clock_bridge:s0_readdata -> cpu_ddr_clock_bridge_s0_translator:av_readdata
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                             // cpu_ddr_clock_bridge_s0_translator:av_debugaccess -> cpu_ddr_clock_bridge:s0_debugaccess
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                           // cpu_ddr_clock_bridge:s0_readdatavalid -> cpu_ddr_clock_bridge_s0_translator:av_readdatavalid
	wire    [3:0] cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                              // cpu_ddr_clock_bridge_s0_translator:av_byteenable -> cpu_ddr_clock_bridge:s0_byteenable
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                           // cpu_ddr_1_clock_bridge:s0_waitrequest -> cpu_ddr_1_clock_bridge_s0_translator:av_waitrequest
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                            // cpu_ddr_1_clock_bridge_s0_translator:av_burstcount -> cpu_ddr_1_clock_bridge:s0_burstcount
	wire   [31:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_writedata;                                             // cpu_ddr_1_clock_bridge_s0_translator:av_writedata -> cpu_ddr_1_clock_bridge:s0_writedata
	wire   [25:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_address;                                               // cpu_ddr_1_clock_bridge_s0_translator:av_address -> cpu_ddr_1_clock_bridge:s0_address
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_write;                                                 // cpu_ddr_1_clock_bridge_s0_translator:av_write -> cpu_ddr_1_clock_bridge:s0_write
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_read;                                                  // cpu_ddr_1_clock_bridge_s0_translator:av_read -> cpu_ddr_1_clock_bridge:s0_read
	wire   [31:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_readdata;                                              // cpu_ddr_1_clock_bridge:s0_readdata -> cpu_ddr_1_clock_bridge_s0_translator:av_readdata
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                           // cpu_ddr_1_clock_bridge_s0_translator:av_debugaccess -> cpu_ddr_1_clock_bridge:s0_debugaccess
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                         // cpu_ddr_1_clock_bridge:s0_readdatavalid -> cpu_ddr_1_clock_bridge_s0_translator:av_readdatavalid
	wire    [3:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                            // cpu_ddr_1_clock_bridge_s0_translator:av_byteenable -> cpu_ddr_1_clock_bridge:s0_byteenable
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                           // slow_peripheral_bridge:s0_waitrequest -> slow_peripheral_bridge_s0_translator:av_waitrequest
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                            // slow_peripheral_bridge_s0_translator:av_burstcount -> slow_peripheral_bridge:s0_burstcount
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata;                                             // slow_peripheral_bridge_s0_translator:av_writedata -> slow_peripheral_bridge:s0_writedata
	wire    [9:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address;                                               // slow_peripheral_bridge_s0_translator:av_address -> slow_peripheral_bridge:s0_address
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write;                                                 // slow_peripheral_bridge_s0_translator:av_write -> slow_peripheral_bridge:s0_write
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read;                                                  // slow_peripheral_bridge_s0_translator:av_read -> slow_peripheral_bridge:s0_read
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata;                                              // slow_peripheral_bridge:s0_readdata -> slow_peripheral_bridge_s0_translator:av_readdata
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                           // slow_peripheral_bridge_s0_translator:av_debugaccess -> slow_peripheral_bridge:s0_debugaccess
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                         // slow_peripheral_bridge:s0_readdatavalid -> slow_peripheral_bridge_s0_translator:av_readdatavalid
	wire    [3:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                            // slow_peripheral_bridge_s0_translator:av_byteenable -> slow_peripheral_bridge:s0_byteenable
	wire          lcd_sgdma_descriptor_read_waitrequest;                                                                          // lcd_sgdma_descriptor_read_translator:av_waitrequest -> lcd_sgdma:descriptor_read_waitrequest
	wire   [31:0] lcd_sgdma_descriptor_read_address;                                                                              // lcd_sgdma:descriptor_read_address -> lcd_sgdma_descriptor_read_translator:av_address
	wire          lcd_sgdma_descriptor_read_read;                                                                                 // lcd_sgdma:descriptor_read_read -> lcd_sgdma_descriptor_read_translator:av_read
	wire   [31:0] lcd_sgdma_descriptor_read_readdata;                                                                             // lcd_sgdma_descriptor_read_translator:av_readdata -> lcd_sgdma:descriptor_read_readdata
	wire          lcd_sgdma_descriptor_read_readdatavalid;                                                                        // lcd_sgdma_descriptor_read_translator:av_readdatavalid -> lcd_sgdma:descriptor_read_readdatavalid
	wire          lcd_sgdma_descriptor_write_waitrequest;                                                                         // lcd_sgdma_descriptor_write_translator:av_waitrequest -> lcd_sgdma:descriptor_write_waitrequest
	wire   [31:0] lcd_sgdma_descriptor_write_writedata;                                                                           // lcd_sgdma:descriptor_write_writedata -> lcd_sgdma_descriptor_write_translator:av_writedata
	wire   [31:0] lcd_sgdma_descriptor_write_address;                                                                             // lcd_sgdma:descriptor_write_address -> lcd_sgdma_descriptor_write_translator:av_address
	wire          lcd_sgdma_descriptor_write_write;                                                                               // lcd_sgdma:descriptor_write_write -> lcd_sgdma_descriptor_write_translator:av_write
	wire          lcd_sgdma_m_read_waitrequest;                                                                                   // lcd_sgdma_m_read_translator:av_waitrequest -> lcd_sgdma:m_read_waitrequest
	wire   [31:0] lcd_sgdma_m_read_address;                                                                                       // lcd_sgdma:m_read_address -> lcd_sgdma_m_read_translator:av_address
	wire          lcd_sgdma_m_read_read;                                                                                          // lcd_sgdma:m_read_read -> lcd_sgdma_m_read_translator:av_read
	wire   [63:0] lcd_sgdma_m_read_readdata;                                                                                      // lcd_sgdma_m_read_translator:av_readdata -> lcd_sgdma:m_read_readdata
	wire          lcd_sgdma_m_read_readdatavalid;                                                                                 // lcd_sgdma_m_read_translator:av_readdatavalid -> lcd_sgdma:m_read_readdatavalid
	wire    [0:0] sdhc_ddr_clock_bridge_m0_burstcount;                                                                            // sdhc_ddr_clock_bridge:m0_burstcount -> sdhc_ddr_clock_bridge_m0_translator:av_burstcount
	wire          sdhc_ddr_clock_bridge_m0_waitrequest;                                                                           // sdhc_ddr_clock_bridge_m0_translator:av_waitrequest -> sdhc_ddr_clock_bridge:m0_waitrequest
	wire   [25:0] sdhc_ddr_clock_bridge_m0_address;                                                                               // sdhc_ddr_clock_bridge:m0_address -> sdhc_ddr_clock_bridge_m0_translator:av_address
	wire   [63:0] sdhc_ddr_clock_bridge_m0_writedata;                                                                             // sdhc_ddr_clock_bridge:m0_writedata -> sdhc_ddr_clock_bridge_m0_translator:av_writedata
	wire          sdhc_ddr_clock_bridge_m0_write;                                                                                 // sdhc_ddr_clock_bridge:m0_write -> sdhc_ddr_clock_bridge_m0_translator:av_write
	wire          sdhc_ddr_clock_bridge_m0_read;                                                                                  // sdhc_ddr_clock_bridge:m0_read -> sdhc_ddr_clock_bridge_m0_translator:av_read
	wire   [63:0] sdhc_ddr_clock_bridge_m0_readdata;                                                                              // sdhc_ddr_clock_bridge_m0_translator:av_readdata -> sdhc_ddr_clock_bridge:m0_readdata
	wire          sdhc_ddr_clock_bridge_m0_debugaccess;                                                                           // sdhc_ddr_clock_bridge:m0_debugaccess -> sdhc_ddr_clock_bridge_m0_translator:av_debugaccess
	wire    [7:0] sdhc_ddr_clock_bridge_m0_byteenable;                                                                            // sdhc_ddr_clock_bridge:m0_byteenable -> sdhc_ddr_clock_bridge_m0_translator:av_byteenable
	wire          sdhc_ddr_clock_bridge_m0_readdatavalid;                                                                         // sdhc_ddr_clock_bridge_m0_translator:av_readdatavalid -> sdhc_ddr_clock_bridge:m0_readdatavalid
	wire    [0:0] cpu_ddr_clock_bridge_m0_burstcount;                                                                             // cpu_ddr_clock_bridge:m0_burstcount -> cpu_ddr_clock_bridge_m0_translator:av_burstcount
	wire          cpu_ddr_clock_bridge_m0_waitrequest;                                                                            // cpu_ddr_clock_bridge_m0_translator:av_waitrequest -> cpu_ddr_clock_bridge:m0_waitrequest
	wire   [26:0] cpu_ddr_clock_bridge_m0_address;                                                                                // cpu_ddr_clock_bridge:m0_address -> cpu_ddr_clock_bridge_m0_translator:av_address
	wire   [31:0] cpu_ddr_clock_bridge_m0_writedata;                                                                              // cpu_ddr_clock_bridge:m0_writedata -> cpu_ddr_clock_bridge_m0_translator:av_writedata
	wire          cpu_ddr_clock_bridge_m0_write;                                                                                  // cpu_ddr_clock_bridge:m0_write -> cpu_ddr_clock_bridge_m0_translator:av_write
	wire          cpu_ddr_clock_bridge_m0_read;                                                                                   // cpu_ddr_clock_bridge:m0_read -> cpu_ddr_clock_bridge_m0_translator:av_read
	wire   [31:0] cpu_ddr_clock_bridge_m0_readdata;                                                                               // cpu_ddr_clock_bridge_m0_translator:av_readdata -> cpu_ddr_clock_bridge:m0_readdata
	wire          cpu_ddr_clock_bridge_m0_debugaccess;                                                                            // cpu_ddr_clock_bridge:m0_debugaccess -> cpu_ddr_clock_bridge_m0_translator:av_debugaccess
	wire    [3:0] cpu_ddr_clock_bridge_m0_byteenable;                                                                             // cpu_ddr_clock_bridge:m0_byteenable -> cpu_ddr_clock_bridge_m0_translator:av_byteenable
	wire          cpu_ddr_clock_bridge_m0_readdatavalid;                                                                          // cpu_ddr_clock_bridge_m0_translator:av_readdatavalid -> cpu_ddr_clock_bridge:m0_readdatavalid
	wire    [0:0] tse_ddr_clock_bridge_m0_burstcount;                                                                             // tse_ddr_clock_bridge:m0_burstcount -> tse_ddr_clock_bridge_m0_translator:av_burstcount
	wire          tse_ddr_clock_bridge_m0_waitrequest;                                                                            // tse_ddr_clock_bridge_m0_translator:av_waitrequest -> tse_ddr_clock_bridge:m0_waitrequest
	wire   [25:0] tse_ddr_clock_bridge_m0_address;                                                                                // tse_ddr_clock_bridge:m0_address -> tse_ddr_clock_bridge_m0_translator:av_address
	wire   [31:0] tse_ddr_clock_bridge_m0_writedata;                                                                              // tse_ddr_clock_bridge:m0_writedata -> tse_ddr_clock_bridge_m0_translator:av_writedata
	wire          tse_ddr_clock_bridge_m0_write;                                                                                  // tse_ddr_clock_bridge:m0_write -> tse_ddr_clock_bridge_m0_translator:av_write
	wire          tse_ddr_clock_bridge_m0_read;                                                                                   // tse_ddr_clock_bridge:m0_read -> tse_ddr_clock_bridge_m0_translator:av_read
	wire   [31:0] tse_ddr_clock_bridge_m0_readdata;                                                                               // tse_ddr_clock_bridge_m0_translator:av_readdata -> tse_ddr_clock_bridge:m0_readdata
	wire          tse_ddr_clock_bridge_m0_debugaccess;                                                                            // tse_ddr_clock_bridge:m0_debugaccess -> tse_ddr_clock_bridge_m0_translator:av_debugaccess
	wire    [3:0] tse_ddr_clock_bridge_m0_byteenable;                                                                             // tse_ddr_clock_bridge:m0_byteenable -> tse_ddr_clock_bridge_m0_translator:av_byteenable
	wire          tse_ddr_clock_bridge_m0_readdatavalid;                                                                          // tse_ddr_clock_bridge_m0_translator:av_readdatavalid -> tse_ddr_clock_bridge:m0_readdatavalid
	wire          ddr2_sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                       // ddr2_sdram:local_ready -> ddr2_sdram_s1_translator:av_waitrequest
	wire          ddr2_sdram_s1_translator_avalon_anti_slave_0_burstcount;                                                        // ddr2_sdram_s1_translator:av_burstcount -> ddr2_sdram:local_size
	wire   [63:0] ddr2_sdram_s1_translator_avalon_anti_slave_0_writedata;                                                         // ddr2_sdram_s1_translator:av_writedata -> ddr2_sdram:local_wdata
	wire   [22:0] ddr2_sdram_s1_translator_avalon_anti_slave_0_address;                                                           // ddr2_sdram_s1_translator:av_address -> ddr2_sdram:local_address
	wire          ddr2_sdram_s1_translator_avalon_anti_slave_0_write;                                                             // ddr2_sdram_s1_translator:av_write -> ddr2_sdram:local_write_req
	wire          ddr2_sdram_s1_translator_avalon_anti_slave_0_beginbursttransfer;                                                // ddr2_sdram_s1_translator:av_beginbursttransfer -> ddr2_sdram:local_burstbegin
	wire          ddr2_sdram_s1_translator_avalon_anti_slave_0_read;                                                              // ddr2_sdram_s1_translator:av_read -> ddr2_sdram:local_read_req
	wire   [63:0] ddr2_sdram_s1_translator_avalon_anti_slave_0_readdata;                                                          // ddr2_sdram:local_rdata -> ddr2_sdram_s1_translator:av_readdata
	wire          ddr2_sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                     // ddr2_sdram:local_rdata_valid -> ddr2_sdram_s1_translator:av_readdatavalid
	wire    [7:0] ddr2_sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                        // ddr2_sdram_s1_translator:av_byteenable -> ddr2_sdram:local_be
	wire          ddr2_sdram_reset_request_n_reset;                                                                               // ddr2_sdram:reset_request_n -> [cmd_xbar_mux_010:reset, ddr2_sdram_s1_translator:reset, ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:reset, ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_010:reset, rsp_xbar_demux_010:reset, rst_controller:reset_in3, rst_controller_001:reset_in3, rst_controller_002:reset_in3, rst_controller_003:reset_in3, rst_controller_004:reset_in3, rst_controller_005:reset_in3, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset]
	wire   [31:0] lcd_sgdma_csr_translator_avalon_anti_slave_0_writedata;                                                         // lcd_sgdma_csr_translator:av_writedata -> lcd_sgdma:csr_writedata
	wire    [3:0] lcd_sgdma_csr_translator_avalon_anti_slave_0_address;                                                           // lcd_sgdma_csr_translator:av_address -> lcd_sgdma:csr_address
	wire          lcd_sgdma_csr_translator_avalon_anti_slave_0_chipselect;                                                        // lcd_sgdma_csr_translator:av_chipselect -> lcd_sgdma:csr_chipselect
	wire          lcd_sgdma_csr_translator_avalon_anti_slave_0_write;                                                             // lcd_sgdma_csr_translator:av_write -> lcd_sgdma:csr_write
	wire          lcd_sgdma_csr_translator_avalon_anti_slave_0_read;                                                              // lcd_sgdma_csr_translator:av_read -> lcd_sgdma:csr_read
	wire   [31:0] lcd_sgdma_csr_translator_avalon_anti_slave_0_readdata;                                                          // lcd_sgdma:csr_readdata -> lcd_sgdma_csr_translator:av_readdata
	wire          sls_sdhc_read_master_waitrequest;                                                                               // sls_sdhc_read_master_translator:av_waitrequest -> sls_sdhc:AvM_rd_waitrequest
	wire   [31:0] sls_sdhc_read_master_address;                                                                                   // sls_sdhc:AvM_rd_address -> sls_sdhc_read_master_translator:av_address
	wire          sls_sdhc_read_master_read;                                                                                      // sls_sdhc:AvM_rd_read_n -> sls_sdhc_read_master_translator:av_read
	wire   [31:0] sls_sdhc_read_master_readdata;                                                                                  // sls_sdhc_read_master_translator:av_readdata -> sls_sdhc:AvM_rd_readdata
	wire    [3:0] sls_sdhc_read_master_byteenable;                                                                                // sls_sdhc:AvM_rd_byteenable -> sls_sdhc_read_master_translator:av_byteenable
	wire          sls_sdhc_read_master_readdatavalid;                                                                             // sls_sdhc_read_master_translator:av_readdatavalid -> sls_sdhc:AvM_rd_readdatavalid
	wire          sls_sdhc_write_master_waitrequest;                                                                              // sls_sdhc_write_master_translator:av_waitrequest -> sls_sdhc:AvM_wr_waitrequest
	wire   [31:0] sls_sdhc_write_master_writedata;                                                                                // sls_sdhc:AvM_wr_writedata -> sls_sdhc_write_master_translator:av_writedata
	wire   [31:0] sls_sdhc_write_master_address;                                                                                  // sls_sdhc:AvM_wr_address -> sls_sdhc_write_master_translator:av_address
	wire          sls_sdhc_write_master_chipselect;                                                                               // sls_sdhc:AvM_wr_chipselect -> sls_sdhc_write_master_translator:av_chipselect
	wire          sls_sdhc_write_master_write;                                                                                    // sls_sdhc:AvM_wr_write_n -> sls_sdhc_write_master_translator:av_write
	wire    [3:0] sls_sdhc_write_master_byteenable;                                                                               // sls_sdhc:AvM_wr_byteenable -> sls_sdhc_write_master_translator:av_byteenable
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                            // sdhc_ddr_clock_bridge:s0_waitrequest -> sdhc_ddr_clock_bridge_s0_translator:av_waitrequest
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                             // sdhc_ddr_clock_bridge_s0_translator:av_burstcount -> sdhc_ddr_clock_bridge:s0_burstcount
	wire   [63:0] sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata;                                              // sdhc_ddr_clock_bridge_s0_translator:av_writedata -> sdhc_ddr_clock_bridge:s0_writedata
	wire   [25:0] sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address;                                                // sdhc_ddr_clock_bridge_s0_translator:av_address -> sdhc_ddr_clock_bridge:s0_address
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write;                                                  // sdhc_ddr_clock_bridge_s0_translator:av_write -> sdhc_ddr_clock_bridge:s0_write
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read;                                                   // sdhc_ddr_clock_bridge_s0_translator:av_read -> sdhc_ddr_clock_bridge:s0_read
	wire   [63:0] sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata;                                               // sdhc_ddr_clock_bridge:s0_readdata -> sdhc_ddr_clock_bridge_s0_translator:av_readdata
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                            // sdhc_ddr_clock_bridge_s0_translator:av_debugaccess -> sdhc_ddr_clock_bridge:s0_debugaccess
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                          // sdhc_ddr_clock_bridge:s0_readdatavalid -> sdhc_ddr_clock_bridge_s0_translator:av_readdatavalid
	wire    [7:0] sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                             // sdhc_ddr_clock_bridge_s0_translator:av_byteenable -> sdhc_ddr_clock_bridge:s0_byteenable
	wire    [0:0] cpu_ddr_1_clock_bridge_m0_burstcount;                                                                           // cpu_ddr_1_clock_bridge:m0_burstcount -> cpu_ddr_1_clock_bridge_m0_translator:av_burstcount
	wire          cpu_ddr_1_clock_bridge_m0_waitrequest;                                                                          // cpu_ddr_1_clock_bridge_m0_translator:av_waitrequest -> cpu_ddr_1_clock_bridge:m0_waitrequest
	wire   [25:0] cpu_ddr_1_clock_bridge_m0_address;                                                                              // cpu_ddr_1_clock_bridge:m0_address -> cpu_ddr_1_clock_bridge_m0_translator:av_address
	wire   [31:0] cpu_ddr_1_clock_bridge_m0_writedata;                                                                            // cpu_ddr_1_clock_bridge:m0_writedata -> cpu_ddr_1_clock_bridge_m0_translator:av_writedata
	wire          cpu_ddr_1_clock_bridge_m0_write;                                                                                // cpu_ddr_1_clock_bridge:m0_write -> cpu_ddr_1_clock_bridge_m0_translator:av_write
	wire          cpu_ddr_1_clock_bridge_m0_read;                                                                                 // cpu_ddr_1_clock_bridge:m0_read -> cpu_ddr_1_clock_bridge_m0_translator:av_read
	wire   [31:0] cpu_ddr_1_clock_bridge_m0_readdata;                                                                             // cpu_ddr_1_clock_bridge_m0_translator:av_readdata -> cpu_ddr_1_clock_bridge:m0_readdata
	wire          cpu_ddr_1_clock_bridge_m0_debugaccess;                                                                          // cpu_ddr_1_clock_bridge:m0_debugaccess -> cpu_ddr_1_clock_bridge_m0_translator:av_debugaccess
	wire    [3:0] cpu_ddr_1_clock_bridge_m0_byteenable;                                                                           // cpu_ddr_1_clock_bridge:m0_byteenable -> cpu_ddr_1_clock_bridge_m0_translator:av_byteenable
	wire          cpu_ddr_1_clock_bridge_m0_readdatavalid;                                                                        // cpu_ddr_1_clock_bridge_m0_translator:av_readdatavalid -> cpu_ddr_1_clock_bridge:m0_readdatavalid
	wire          ddr2_sdram_1_s1_translator_avalon_anti_slave_0_waitrequest;                                                     // ddr2_sdram_1:local_ready -> ddr2_sdram_1_s1_translator:av_waitrequest
	wire    [1:0] ddr2_sdram_1_s1_translator_avalon_anti_slave_0_burstcount;                                                      // ddr2_sdram_1_s1_translator:av_burstcount -> ddr2_sdram_1:local_size
	wire   [31:0] ddr2_sdram_1_s1_translator_avalon_anti_slave_0_writedata;                                                       // ddr2_sdram_1_s1_translator:av_writedata -> ddr2_sdram_1:local_wdata
	wire   [23:0] ddr2_sdram_1_s1_translator_avalon_anti_slave_0_address;                                                         // ddr2_sdram_1_s1_translator:av_address -> ddr2_sdram_1:local_address
	wire          ddr2_sdram_1_s1_translator_avalon_anti_slave_0_write;                                                           // ddr2_sdram_1_s1_translator:av_write -> ddr2_sdram_1:local_write_req
	wire          ddr2_sdram_1_s1_translator_avalon_anti_slave_0_beginbursttransfer;                                              // ddr2_sdram_1_s1_translator:av_beginbursttransfer -> ddr2_sdram_1:local_burstbegin
	wire          ddr2_sdram_1_s1_translator_avalon_anti_slave_0_read;                                                            // ddr2_sdram_1_s1_translator:av_read -> ddr2_sdram_1:local_read_req
	wire   [31:0] ddr2_sdram_1_s1_translator_avalon_anti_slave_0_readdata;                                                        // ddr2_sdram_1:local_rdata -> ddr2_sdram_1_s1_translator:av_readdata
	wire          ddr2_sdram_1_s1_translator_avalon_anti_slave_0_readdatavalid;                                                   // ddr2_sdram_1:local_rdata_valid -> ddr2_sdram_1_s1_translator:av_readdatavalid
	wire    [3:0] ddr2_sdram_1_s1_translator_avalon_anti_slave_0_byteenable;                                                      // ddr2_sdram_1_s1_translator:av_byteenable -> ddr2_sdram_1:local_be
	wire          ddr2_sdram_1_reset_request_n_reset;                                                                             // ddr2_sdram_1:reset_request_n -> [ddr2_sdram_1_s1_translator:reset, ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:reset, ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_013:reset, rsp_xbar_demux_013:reset, rst_controller:reset_in4, rst_controller_001:reset_in4, rst_controller_002:reset_in4, rst_controller_003:reset_in4, rst_controller_004:reset_in4, rst_controller_005:reset_in4]
	wire    [0:0] slow_peripheral_bridge_m0_burstcount;                                                                           // slow_peripheral_bridge:m0_burstcount -> slow_peripheral_bridge_m0_translator:av_burstcount
	wire          slow_peripheral_bridge_m0_waitrequest;                                                                          // slow_peripheral_bridge_m0_translator:av_waitrequest -> slow_peripheral_bridge:m0_waitrequest
	wire    [9:0] slow_peripheral_bridge_m0_address;                                                                              // slow_peripheral_bridge:m0_address -> slow_peripheral_bridge_m0_translator:av_address
	wire   [31:0] slow_peripheral_bridge_m0_writedata;                                                                            // slow_peripheral_bridge:m0_writedata -> slow_peripheral_bridge_m0_translator:av_writedata
	wire          slow_peripheral_bridge_m0_write;                                                                                // slow_peripheral_bridge:m0_write -> slow_peripheral_bridge_m0_translator:av_write
	wire          slow_peripheral_bridge_m0_read;                                                                                 // slow_peripheral_bridge:m0_read -> slow_peripheral_bridge_m0_translator:av_read
	wire   [31:0] slow_peripheral_bridge_m0_readdata;                                                                             // slow_peripheral_bridge_m0_translator:av_readdata -> slow_peripheral_bridge:m0_readdata
	wire          slow_peripheral_bridge_m0_debugaccess;                                                                          // slow_peripheral_bridge:m0_debugaccess -> slow_peripheral_bridge_m0_translator:av_debugaccess
	wire    [3:0] slow_peripheral_bridge_m0_byteenable;                                                                           // slow_peripheral_bridge:m0_byteenable -> slow_peripheral_bridge_m0_translator:av_byteenable
	wire          slow_peripheral_bridge_m0_readdatavalid;                                                                        // slow_peripheral_bridge_m0_translator:av_readdatavalid -> slow_peripheral_bridge:m0_readdatavalid
	wire   [31:0] button_pio_s1_translator_avalon_anti_slave_0_writedata;                                                         // button_pio_s1_translator:av_writedata -> button_pio:writedata
	wire    [1:0] button_pio_s1_translator_avalon_anti_slave_0_address;                                                           // button_pio_s1_translator:av_address -> button_pio:address
	wire          button_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                        // button_pio_s1_translator:av_chipselect -> button_pio:chipselect
	wire          button_pio_s1_translator_avalon_anti_slave_0_write;                                                             // button_pio_s1_translator:av_write -> button_pio:write_n
	wire   [31:0] button_pio_s1_translator_avalon_anti_slave_0_readdata;                                                          // button_pio:readdata -> button_pio_s1_translator:av_readdata
	wire   [15:0] high_res_timer_s1_translator_avalon_anti_slave_0_writedata;                                                     // high_res_timer_s1_translator:av_writedata -> high_res_timer:writedata
	wire    [2:0] high_res_timer_s1_translator_avalon_anti_slave_0_address;                                                       // high_res_timer_s1_translator:av_address -> high_res_timer:address
	wire          high_res_timer_s1_translator_avalon_anti_slave_0_chipselect;                                                    // high_res_timer_s1_translator:av_chipselect -> high_res_timer:chipselect
	wire          high_res_timer_s1_translator_avalon_anti_slave_0_write;                                                         // high_res_timer_s1_translator:av_write -> high_res_timer:write_n
	wire   [15:0] high_res_timer_s1_translator_avalon_anti_slave_0_readdata;                                                      // high_res_timer:readdata -> high_res_timer_s1_translator:av_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                         // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                           // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                             // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                          // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                               // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                                // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                            // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] uart1_s1_translator_avalon_anti_slave_0_writedata;                                                              // uart1_s1_translator:av_writedata -> uart1:writedata
	wire    [2:0] uart1_s1_translator_avalon_anti_slave_0_address;                                                                // uart1_s1_translator:av_address -> uart1:address
	wire          uart1_s1_translator_avalon_anti_slave_0_chipselect;                                                             // uart1_s1_translator:av_chipselect -> uart1:chipselect
	wire          uart1_s1_translator_avalon_anti_slave_0_write;                                                                  // uart1_s1_translator:av_write -> uart1:write_n
	wire          uart1_s1_translator_avalon_anti_slave_0_read;                                                                   // uart1_s1_translator:av_read -> uart1:read_n
	wire   [15:0] uart1_s1_translator_avalon_anti_slave_0_readdata;                                                               // uart1:readdata -> uart1_s1_translator:av_readdata
	wire          uart1_s1_translator_avalon_anti_slave_0_begintransfer;                                                          // uart1_s1_translator:av_begintransfer -> uart1:begintransfer
	wire   [31:0] led_pio_s1_translator_avalon_anti_slave_0_writedata;                                                            // led_pio_s1_translator:av_writedata -> led_pio:writedata
	wire    [1:0] led_pio_s1_translator_avalon_anti_slave_0_address;                                                              // led_pio_s1_translator:av_address -> led_pio:address
	wire          led_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                           // led_pio_s1_translator:av_chipselect -> led_pio:chipselect
	wire          led_pio_s1_translator_avalon_anti_slave_0_write;                                                                // led_pio_s1_translator:av_write -> led_pio:write_n
	wire   [31:0] led_pio_s1_translator_avalon_anti_slave_0_readdata;                                                             // led_pio:readdata -> led_pio_s1_translator:av_readdata
	wire   [31:0] performance_counter_control_slave_translator_avalon_anti_slave_0_writedata;                                     // performance_counter_control_slave_translator:av_writedata -> performance_counter:writedata
	wire    [2:0] performance_counter_control_slave_translator_avalon_anti_slave_0_address;                                       // performance_counter_control_slave_translator:av_address -> performance_counter:address
	wire          performance_counter_control_slave_translator_avalon_anti_slave_0_write;                                         // performance_counter_control_slave_translator:av_write -> performance_counter:write
	wire   [31:0] performance_counter_control_slave_translator_avalon_anti_slave_0_readdata;                                      // performance_counter:readdata -> performance_counter_control_slave_translator:av_readdata
	wire          performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer;                                 // performance_counter_control_slave_translator:av_begintransfer -> performance_counter:begintransfer
	wire   [15:0] pll_s1_translator_avalon_anti_slave_0_writedata;                                                                // pll_s1_translator:av_writedata -> pll:writedata
	wire    [2:0] pll_s1_translator_avalon_anti_slave_0_address;                                                                  // pll_s1_translator:av_address -> pll:address
	wire          pll_s1_translator_avalon_anti_slave_0_chipselect;                                                               // pll_s1_translator:av_chipselect -> pll:chipselect
	wire          pll_s1_translator_avalon_anti_slave_0_write;                                                                    // pll_s1_translator:av_write -> pll:write
	wire          pll_s1_translator_avalon_anti_slave_0_read;                                                                     // pll_s1_translator:av_read -> pll:read
	wire   [15:0] pll_s1_translator_avalon_anti_slave_0_readdata;                                                                 // pll:readdata -> pll_s1_translator:av_readdata
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata;                                                      // sys_clk_timer_s1_translator:av_writedata -> sys_clk_timer:writedata
	wire    [2:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_address;                                                        // sys_clk_timer_s1_translator:av_address -> sys_clk_timer:address
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect;                                                     // sys_clk_timer_s1_translator:av_chipselect -> sys_clk_timer:chipselect
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_write;                                                          // sys_clk_timer_s1_translator:av_write -> sys_clk_timer:write_n
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata;                                                       // sys_clk_timer:readdata -> sys_clk_timer_s1_translator:av_readdata
	wire          sysid_control_slave_translator_avalon_anti_slave_0_address;                                                     // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                                    // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [31:0] lcd_i2c_en_s1_translator_avalon_anti_slave_0_writedata;                                                         // lcd_i2c_en_s1_translator:av_writedata -> lcd_i2c_en:writedata
	wire    [1:0] lcd_i2c_en_s1_translator_avalon_anti_slave_0_address;                                                           // lcd_i2c_en_s1_translator:av_address -> lcd_i2c_en:address
	wire          lcd_i2c_en_s1_translator_avalon_anti_slave_0_chipselect;                                                        // lcd_i2c_en_s1_translator:av_chipselect -> lcd_i2c_en:chipselect
	wire          lcd_i2c_en_s1_translator_avalon_anti_slave_0_write;                                                             // lcd_i2c_en_s1_translator:av_write -> lcd_i2c_en:write_n
	wire   [31:0] lcd_i2c_en_s1_translator_avalon_anti_slave_0_readdata;                                                          // lcd_i2c_en:readdata -> lcd_i2c_en_s1_translator:av_readdata
	wire   [31:0] lcd_i2c_scl_s1_translator_avalon_anti_slave_0_writedata;                                                        // lcd_i2c_scl_s1_translator:av_writedata -> lcd_i2c_scl:writedata
	wire    [1:0] lcd_i2c_scl_s1_translator_avalon_anti_slave_0_address;                                                          // lcd_i2c_scl_s1_translator:av_address -> lcd_i2c_scl:address
	wire          lcd_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect;                                                       // lcd_i2c_scl_s1_translator:av_chipselect -> lcd_i2c_scl:chipselect
	wire          lcd_i2c_scl_s1_translator_avalon_anti_slave_0_write;                                                            // lcd_i2c_scl_s1_translator:av_write -> lcd_i2c_scl:write_n
	wire   [31:0] lcd_i2c_scl_s1_translator_avalon_anti_slave_0_readdata;                                                         // lcd_i2c_scl:readdata -> lcd_i2c_scl_s1_translator:av_readdata
	wire   [31:0] lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_writedata;                                                       // lcd_i2c_sdat_s1_translator:av_writedata -> lcd_i2c_sdat:writedata
	wire    [1:0] lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_address;                                                         // lcd_i2c_sdat_s1_translator:av_address -> lcd_i2c_sdat:address
	wire          lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_chipselect;                                                      // lcd_i2c_sdat_s1_translator:av_chipselect -> lcd_i2c_sdat:chipselect
	wire          lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_write;                                                           // lcd_i2c_sdat_s1_translator:av_write -> lcd_i2c_sdat:write_n
	wire   [31:0] lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_readdata;                                                        // lcd_i2c_sdat:readdata -> lcd_i2c_sdat_s1_translator:av_readdata
	wire   [31:0] pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_writedata;                                                  // pio_id_eeprom_dat_s1_translator:av_writedata -> pio_id_eeprom_dat:writedata
	wire    [1:0] pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_address;                                                    // pio_id_eeprom_dat_s1_translator:av_address -> pio_id_eeprom_dat:address
	wire          pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_chipselect;                                                 // pio_id_eeprom_dat_s1_translator:av_chipselect -> pio_id_eeprom_dat:chipselect
	wire          pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_write;                                                      // pio_id_eeprom_dat_s1_translator:av_write -> pio_id_eeprom_dat:write_n
	wire   [31:0] pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_readdata;                                                   // pio_id_eeprom_dat:readdata -> pio_id_eeprom_dat_s1_translator:av_readdata
	wire   [31:0] pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_writedata;                                                  // pio_id_eeprom_scl_s1_translator:av_writedata -> pio_id_eeprom_scl:writedata
	wire    [1:0] pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_address;                                                    // pio_id_eeprom_scl_s1_translator:av_address -> pio_id_eeprom_scl:address
	wire          pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_chipselect;                                                 // pio_id_eeprom_scl_s1_translator:av_chipselect -> pio_id_eeprom_scl:chipselect
	wire          pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_write;                                                      // pio_id_eeprom_scl_s1_translator:av_write -> pio_id_eeprom_scl:write_n
	wire   [31:0] pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_readdata;                                                   // pio_id_eeprom_scl:readdata -> pio_id_eeprom_scl_s1_translator:av_readdata
	wire   [31:0] touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_writedata;                                              // touch_panel_pen_irq_n_s1_translator:av_writedata -> touch_panel_pen_irq_n:writedata
	wire    [1:0] touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_address;                                                // touch_panel_pen_irq_n_s1_translator:av_address -> touch_panel_pen_irq_n:address
	wire          touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_chipselect;                                             // touch_panel_pen_irq_n_s1_translator:av_chipselect -> touch_panel_pen_irq_n:chipselect
	wire          touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_write;                                                  // touch_panel_pen_irq_n_s1_translator:av_write -> touch_panel_pen_irq_n:write_n
	wire   [31:0] touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_readdata;                                               // touch_panel_pen_irq_n:readdata -> touch_panel_pen_irq_n_s1_translator:av_readdata
	wire   [15:0] touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_writedata;                                      // touch_panel_spi_spi_control_port_translator:av_writedata -> touch_panel_spi:data_from_cpu
	wire    [2:0] touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_address;                                        // touch_panel_spi_spi_control_port_translator:av_address -> touch_panel_spi:mem_addr
	wire          touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_chipselect;                                     // touch_panel_spi_spi_control_port_translator:av_chipselect -> touch_panel_spi:spi_select
	wire          touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_write;                                          // touch_panel_spi_spi_control_port_translator:av_write -> touch_panel_spi:write_n
	wire          touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_read;                                           // touch_panel_spi_spi_control_port_translator:av_read -> touch_panel_spi:read_n
	wire   [15:0] touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_readdata;                                       // touch_panel_spi:data_to_cpu -> touch_panel_spi_spi_control_port_translator:av_readdata
	wire          sgdma_rx_m_write_waitrequest;                                                                                   // sgdma_rx_m_write_translator:av_waitrequest -> sgdma_rx:m_write_waitrequest
	wire   [31:0] sgdma_rx_m_write_writedata;                                                                                     // sgdma_rx:m_write_writedata -> sgdma_rx_m_write_translator:av_writedata
	wire   [31:0] sgdma_rx_m_write_address;                                                                                       // sgdma_rx:m_write_address -> sgdma_rx_m_write_translator:av_address
	wire          sgdma_rx_m_write_write;                                                                                         // sgdma_rx:m_write_write -> sgdma_rx_m_write_translator:av_write
	wire    [3:0] sgdma_rx_m_write_byteenable;                                                                                    // sgdma_rx:m_write_byteenable -> sgdma_rx_m_write_translator:av_byteenable
	wire          sgdma_tx_m_read_waitrequest;                                                                                    // sgdma_tx_m_read_translator:av_waitrequest -> sgdma_tx:m_read_waitrequest
	wire   [31:0] sgdma_tx_m_read_address;                                                                                        // sgdma_tx:m_read_address -> sgdma_tx_m_read_translator:av_address
	wire          sgdma_tx_m_read_read;                                                                                           // sgdma_tx:m_read_read -> sgdma_tx_m_read_translator:av_read
	wire   [31:0] sgdma_tx_m_read_readdata;                                                                                       // sgdma_tx_m_read_translator:av_readdata -> sgdma_tx:m_read_readdata
	wire          sgdma_tx_m_read_readdatavalid;                                                                                  // sgdma_tx_m_read_translator:av_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire          tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                             // tse_ddr_clock_bridge:s0_waitrequest -> tse_ddr_clock_bridge_s0_translator:av_waitrequest
	wire          tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                              // tse_ddr_clock_bridge_s0_translator:av_burstcount -> tse_ddr_clock_bridge:s0_burstcount
	wire   [31:0] tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata;                                               // tse_ddr_clock_bridge_s0_translator:av_writedata -> tse_ddr_clock_bridge:s0_writedata
	wire   [25:0] tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address;                                                 // tse_ddr_clock_bridge_s0_translator:av_address -> tse_ddr_clock_bridge:s0_address
	wire          tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write;                                                   // tse_ddr_clock_bridge_s0_translator:av_write -> tse_ddr_clock_bridge:s0_write
	wire          tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read;                                                    // tse_ddr_clock_bridge_s0_translator:av_read -> tse_ddr_clock_bridge:s0_read
	wire   [31:0] tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata;                                                // tse_ddr_clock_bridge:s0_readdata -> tse_ddr_clock_bridge_s0_translator:av_readdata
	wire          tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                             // tse_ddr_clock_bridge_s0_translator:av_debugaccess -> tse_ddr_clock_bridge:s0_debugaccess
	wire          tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                           // tse_ddr_clock_bridge:s0_readdatavalid -> tse_ddr_clock_bridge_s0_translator:av_readdatavalid
	wire    [3:0] tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                              // tse_ddr_clock_bridge_s0_translator:av_byteenable -> tse_ddr_clock_bridge:s0_byteenable
	wire    [0:0] pipeline_bridge_before_tristate_bridge_m0_burstcount;                                                           // pipeline_bridge_before_tristate_bridge:m0_burstcount -> pipeline_bridge_before_tristate_bridge_m0_translator:av_burstcount
	wire          pipeline_bridge_before_tristate_bridge_m0_waitrequest;                                                          // pipeline_bridge_before_tristate_bridge_m0_translator:av_waitrequest -> pipeline_bridge_before_tristate_bridge:m0_waitrequest
	wire   [26:0] pipeline_bridge_before_tristate_bridge_m0_address;                                                              // pipeline_bridge_before_tristate_bridge:m0_address -> pipeline_bridge_before_tristate_bridge_m0_translator:av_address
	wire   [31:0] pipeline_bridge_before_tristate_bridge_m0_writedata;                                                            // pipeline_bridge_before_tristate_bridge:m0_writedata -> pipeline_bridge_before_tristate_bridge_m0_translator:av_writedata
	wire          pipeline_bridge_before_tristate_bridge_m0_write;                                                                // pipeline_bridge_before_tristate_bridge:m0_write -> pipeline_bridge_before_tristate_bridge_m0_translator:av_write
	wire          pipeline_bridge_before_tristate_bridge_m0_read;                                                                 // pipeline_bridge_before_tristate_bridge:m0_read -> pipeline_bridge_before_tristate_bridge_m0_translator:av_read
	wire   [31:0] pipeline_bridge_before_tristate_bridge_m0_readdata;                                                             // pipeline_bridge_before_tristate_bridge_m0_translator:av_readdata -> pipeline_bridge_before_tristate_bridge:m0_readdata
	wire          pipeline_bridge_before_tristate_bridge_m0_debugaccess;                                                          // pipeline_bridge_before_tristate_bridge:m0_debugaccess -> pipeline_bridge_before_tristate_bridge_m0_translator:av_debugaccess
	wire    [3:0] pipeline_bridge_before_tristate_bridge_m0_byteenable;                                                           // pipeline_bridge_before_tristate_bridge:m0_byteenable -> pipeline_bridge_before_tristate_bridge_m0_translator:av_byteenable
	wire          pipeline_bridge_before_tristate_bridge_m0_readdatavalid;                                                        // pipeline_bridge_before_tristate_bridge_m0_translator:av_readdatavalid -> pipeline_bridge_before_tristate_bridge:m0_readdatavalid
	wire          ext_flash_uas_translator_avalon_anti_slave_0_waitrequest;                                                       // ext_flash:uas_waitrequest -> ext_flash_uas_translator:av_waitrequest
	wire    [1:0] ext_flash_uas_translator_avalon_anti_slave_0_burstcount;                                                        // ext_flash_uas_translator:av_burstcount -> ext_flash:uas_burstcount
	wire   [15:0] ext_flash_uas_translator_avalon_anti_slave_0_writedata;                                                         // ext_flash_uas_translator:av_writedata -> ext_flash:uas_writedata
	wire   [25:0] ext_flash_uas_translator_avalon_anti_slave_0_address;                                                           // ext_flash_uas_translator:av_address -> ext_flash:uas_address
	wire          ext_flash_uas_translator_avalon_anti_slave_0_lock;                                                              // ext_flash_uas_translator:av_lock -> ext_flash:uas_lock
	wire          ext_flash_uas_translator_avalon_anti_slave_0_write;                                                             // ext_flash_uas_translator:av_write -> ext_flash:uas_write
	wire          ext_flash_uas_translator_avalon_anti_slave_0_read;                                                              // ext_flash_uas_translator:av_read -> ext_flash:uas_read
	wire   [15:0] ext_flash_uas_translator_avalon_anti_slave_0_readdata;                                                          // ext_flash:uas_readdata -> ext_flash_uas_translator:av_readdata
	wire          ext_flash_uas_translator_avalon_anti_slave_0_debugaccess;                                                       // ext_flash_uas_translator:av_debugaccess -> ext_flash:uas_debugaccess
	wire          ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid;                                                     // ext_flash:uas_readdatavalid -> ext_flash_uas_translator:av_readdatavalid
	wire    [1:0] ext_flash_uas_translator_avalon_anti_slave_0_byteenable;                                                        // ext_flash_uas_translator:av_byteenable -> ext_flash:uas_byteenable
	wire          max2_uas_translator_avalon_anti_slave_0_waitrequest;                                                            // max2:uas_waitrequest -> max2_uas_translator:av_waitrequest
	wire    [2:0] max2_uas_translator_avalon_anti_slave_0_burstcount;                                                             // max2_uas_translator:av_burstcount -> max2:uas_burstcount
	wire   [31:0] max2_uas_translator_avalon_anti_slave_0_writedata;                                                              // max2_uas_translator:av_writedata -> max2:uas_writedata
	wire    [4:0] max2_uas_translator_avalon_anti_slave_0_address;                                                                // max2_uas_translator:av_address -> max2:uas_address
	wire          max2_uas_translator_avalon_anti_slave_0_lock;                                                                   // max2_uas_translator:av_lock -> max2:uas_lock
	wire          max2_uas_translator_avalon_anti_slave_0_write;                                                                  // max2_uas_translator:av_write -> max2:uas_write
	wire          max2_uas_translator_avalon_anti_slave_0_read;                                                                   // max2_uas_translator:av_read -> max2:uas_read
	wire   [31:0] max2_uas_translator_avalon_anti_slave_0_readdata;                                                               // max2:uas_readdata -> max2_uas_translator:av_readdata
	wire          max2_uas_translator_avalon_anti_slave_0_debugaccess;                                                            // max2_uas_translator:av_debugaccess -> max2:uas_debugaccess
	wire          max2_uas_translator_avalon_anti_slave_0_readdatavalid;                                                          // max2:uas_readdatavalid -> max2_uas_translator:av_readdatavalid
	wire    [3:0] max2_uas_translator_avalon_anti_slave_0_byteenable;                                                             // max2_uas_translator:av_byteenable -> max2:uas_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                               // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                                // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                                 // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_address;                                                   // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                                      // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                                     // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                                      // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                                  // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                               // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                                // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                             // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                                        // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                                         // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                                          // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                            // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                               // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                              // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                               // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                                           // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                                        // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                                         // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                      // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest;                                      // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_read_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount;                                       // sgdma_rx_descriptor_read_translator:uav_burstcount -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata;                                        // sgdma_rx_descriptor_read_translator:uav_writedata -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address;                                          // sgdma_rx_descriptor_read_translator:uav_address -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock;                                             // sgdma_rx_descriptor_read_translator:uav_lock -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write;                                            // sgdma_rx_descriptor_read_translator:uav_write -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read;                                             // sgdma_rx_descriptor_read_translator:uav_read -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata;                                         // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_read_translator:uav_readdata
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess;                                      // sgdma_rx_descriptor_read_translator:uav_debugaccess -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable;                                       // sgdma_rx_descriptor_read_translator:uav_byteenable -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                                    // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_read_translator:uav_readdatavalid
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest;                                     // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_write_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount;                                      // sgdma_rx_descriptor_write_translator:uav_burstcount -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata;                                       // sgdma_rx_descriptor_write_translator:uav_writedata -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address;                                         // sgdma_rx_descriptor_write_translator:uav_address -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock;                                            // sgdma_rx_descriptor_write_translator:uav_lock -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write;                                           // sgdma_rx_descriptor_write_translator:uav_write -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read;                                            // sgdma_rx_descriptor_write_translator:uav_read -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata;                                        // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_write_translator:uav_readdata
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess;                                     // sgdma_rx_descriptor_write_translator:uav_debugaccess -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable;                                      // sgdma_rx_descriptor_write_translator:uav_byteenable -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                                   // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_write_translator:uav_readdatavalid
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest;                                      // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_read_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount;                                       // sgdma_tx_descriptor_read_translator:uav_burstcount -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata;                                        // sgdma_tx_descriptor_read_translator:uav_writedata -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address;                                          // sgdma_tx_descriptor_read_translator:uav_address -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock;                                             // sgdma_tx_descriptor_read_translator:uav_lock -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write;                                            // sgdma_tx_descriptor_read_translator:uav_write -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read;                                             // sgdma_tx_descriptor_read_translator:uav_read -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata;                                         // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_read_translator:uav_readdata
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess;                                      // sgdma_tx_descriptor_read_translator:uav_debugaccess -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable;                                       // sgdma_tx_descriptor_read_translator:uav_byteenable -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                                    // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_read_translator:uav_readdatavalid
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest;                                     // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_write_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount;                                      // sgdma_tx_descriptor_write_translator:uav_burstcount -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata;                                       // sgdma_tx_descriptor_write_translator:uav_writedata -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address;                                         // sgdma_tx_descriptor_write_translator:uav_address -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock;                                            // sgdma_tx_descriptor_write_translator:uav_lock -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write;                                           // sgdma_tx_descriptor_write_translator:uav_write -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read;                                            // sgdma_tx_descriptor_write_translator:uav_read -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata;                                        // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_write_translator:uav_readdata
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess;                                     // sgdma_tx_descriptor_write_translator:uav_debugaccess -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable;                                      // sgdma_tx_descriptor_write_translator:uav_byteenable -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                                   // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_write_translator:uav_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // descriptor_memory_s1_translator:uav_waitrequest -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> descriptor_memory_s1_translator:uav_burstcount
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> descriptor_memory_s1_translator:uav_writedata
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> descriptor_memory_s1_translator:uav_address
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> descriptor_memory_s1_translator:uav_write
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> descriptor_memory_s1_translator:uav_lock
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> descriptor_memory_s1_translator:uav_read
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // descriptor_memory_s1_translator:uav_readdata -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // descriptor_memory_s1_translator:uav_readdatavalid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> descriptor_memory_s1_translator:uav_debugaccess
	wire    [3:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> descriptor_memory_s1_translator:uav_byteenable
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // sgdma_rx_csr_translator:uav_waitrequest -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_rx_csr_translator:uav_burstcount
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_rx_csr_translator:uav_writedata
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address;                                              // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_rx_csr_translator:uav_address
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write;                                                // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_rx_csr_translator:uav_write
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_rx_csr_translator:uav_lock
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read;                                                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_rx_csr_translator:uav_read
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // sgdma_rx_csr_translator:uav_readdata -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // sgdma_rx_csr_translator:uav_readdatavalid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_rx_csr_translator:uav_debugaccess
	wire    [3:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_rx_csr_translator:uav_byteenable
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // sgdma_tx_csr_translator:uav_waitrequest -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_tx_csr_translator:uav_burstcount
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_tx_csr_translator:uav_writedata
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address;                                              // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_tx_csr_translator:uav_address
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write;                                                // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_tx_csr_translator:uav_write
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_tx_csr_translator:uav_lock
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read;                                                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_tx_csr_translator:uav_read
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // sgdma_tx_csr_translator:uav_readdata -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // sgdma_tx_csr_translator:uav_readdatavalid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_tx_csr_translator:uav_debugaccess
	wire    [3:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_tx_csr_translator:uav_byteenable
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // tse_mac_control_port_translator:uav_waitrequest -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> tse_mac_control_port_translator:uav_burstcount
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> tse_mac_control_port_translator:uav_writedata
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address;                                      // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_address -> tse_mac_control_port_translator:uav_address
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write;                                        // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_write -> tse_mac_control_port_translator:uav_write
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                                         // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> tse_mac_control_port_translator:uav_lock
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read;                                         // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_read -> tse_mac_control_port_translator:uav_read
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // tse_mac_control_port_translator:uav_readdata -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // tse_mac_control_port_translator:uav_readdatavalid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> tse_mac_control_port_translator:uav_debugaccess
	wire    [3:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> tse_mac_control_port_translator:uav_byteenable
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // sls_sdhc_control_translator:uav_waitrequest -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_burstcount -> sls_sdhc_control_translator:uav_burstcount
	wire   [31:0] sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_writedata -> sls_sdhc_control_translator:uav_writedata
	wire   [31:0] sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_address;                                          // sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_address -> sls_sdhc_control_translator:uav_address
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_write;                                            // sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_write -> sls_sdhc_control_translator:uav_write
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_lock;                                             // sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_lock -> sls_sdhc_control_translator:uav_lock
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_read;                                             // sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_read -> sls_sdhc_control_translator:uav_read
	wire   [31:0] sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // sls_sdhc_control_translator:uav_readdata -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // sls_sdhc_control_translator:uav_readdatavalid -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sls_sdhc_control_translator:uav_debugaccess
	wire    [3:0] sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // sls_sdhc_control_translator_avalon_universal_slave_0_agent:m0_byteenable -> sls_sdhc_control_translator:uav_byteenable
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rf_source_valid -> sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rf_source_data -> sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                // sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                 // sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // pipeline_bridge_before_tristate_bridge_s0_translator:uav_waitrequest -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> pipeline_bridge_before_tristate_bridge_s0_translator:uav_burstcount
	wire   [31:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;               // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> pipeline_bridge_before_tristate_bridge_s0_translator:uav_writedata
	wire   [31:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                 // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> pipeline_bridge_before_tristate_bridge_s0_translator:uav_address
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                   // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> pipeline_bridge_before_tristate_bridge_s0_translator:uav_write
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                    // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> pipeline_bridge_before_tristate_bridge_s0_translator:uav_lock
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                    // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> pipeline_bridge_before_tristate_bridge_s0_translator:uav_read
	wire   [31:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                // pipeline_bridge_before_tristate_bridge_s0_translator:uav_readdata -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // pipeline_bridge_before_tristate_bridge_s0_translator:uav_readdatavalid -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pipeline_bridge_before_tristate_bridge_s0_translator:uav_debugaccess
	wire    [3:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> pipeline_bridge_before_tristate_bridge_s0_translator:uav_byteenable
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;             // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // cpu_ddr_clock_bridge_s0_translator:uav_waitrequest -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_ddr_clock_bridge_s0_translator:uav_burstcount
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_ddr_clock_bridge_s0_translator:uav_writedata
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                                   // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> cpu_ddr_clock_bridge_s0_translator:uav_address
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                                     // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> cpu_ddr_clock_bridge_s0_translator:uav_write
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                      // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_ddr_clock_bridge_s0_translator:uav_lock
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                                      // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> cpu_ddr_clock_bridge_s0_translator:uav_read
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // cpu_ddr_clock_bridge_s0_translator:uav_readdata -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // cpu_ddr_clock_bridge_s0_translator:uav_readdatavalid -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_ddr_clock_bridge_s0_translator:uav_debugaccess
	wire    [3:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_ddr_clock_bridge_s0_translator:uav_byteenable
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                               // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // cpu_ddr_1_clock_bridge_s0_translator:uav_waitrequest -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_ddr_1_clock_bridge_s0_translator:uav_burstcount
	wire   [31:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                               // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_ddr_1_clock_bridge_s0_translator:uav_writedata
	wire   [31:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                                 // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> cpu_ddr_1_clock_bridge_s0_translator:uav_address
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                                   // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> cpu_ddr_1_clock_bridge_s0_translator:uav_write
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                    // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_ddr_1_clock_bridge_s0_translator:uav_lock
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                                    // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> cpu_ddr_1_clock_bridge_s0_translator:uav_read
	wire   [31:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                // cpu_ddr_1_clock_bridge_s0_translator:uav_readdata -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // cpu_ddr_1_clock_bridge_s0_translator:uav_readdatavalid -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_ddr_1_clock_bridge_s0_translator:uav_debugaccess
	wire    [3:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_ddr_1_clock_bridge_s0_translator:uav_byteenable
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                             // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // slow_peripheral_bridge_s0_translator:uav_waitrequest -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> slow_peripheral_bridge_s0_translator:uav_burstcount
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                               // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> slow_peripheral_bridge_s0_translator:uav_writedata
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                                 // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> slow_peripheral_bridge_s0_translator:uav_address
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                                   // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> slow_peripheral_bridge_s0_translator:uav_write
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                    // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> slow_peripheral_bridge_s0_translator:uav_lock
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                                    // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> slow_peripheral_bridge_s0_translator:uav_read
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                // slow_peripheral_bridge_s0_translator:uav_readdata -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // slow_peripheral_bridge_s0_translator:uav_readdatavalid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> slow_peripheral_bridge_s0_translator:uav_debugaccess
	wire    [3:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> slow_peripheral_bridge_s0_translator:uav_byteenable
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                             // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_waitrequest;                                     // lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> lcd_sgdma_descriptor_read_translator:uav_waitrequest
	wire    [2:0] lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_burstcount;                                      // lcd_sgdma_descriptor_read_translator:uav_burstcount -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_writedata;                                       // lcd_sgdma_descriptor_read_translator:uav_writedata -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_address;                                         // lcd_sgdma_descriptor_read_translator:uav_address -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_lock;                                            // lcd_sgdma_descriptor_read_translator:uav_lock -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_write;                                           // lcd_sgdma_descriptor_read_translator:uav_write -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_read;                                            // lcd_sgdma_descriptor_read_translator:uav_read -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_readdata;                                        // lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> lcd_sgdma_descriptor_read_translator:uav_readdata
	wire          lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_debugaccess;                                     // lcd_sgdma_descriptor_read_translator:uav_debugaccess -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_byteenable;                                      // lcd_sgdma_descriptor_read_translator:uav_byteenable -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                                   // lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> lcd_sgdma_descriptor_read_translator:uav_readdatavalid
	wire          lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_waitrequest;                                    // lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> lcd_sgdma_descriptor_write_translator:uav_waitrequest
	wire    [2:0] lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_burstcount;                                     // lcd_sgdma_descriptor_write_translator:uav_burstcount -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_writedata;                                      // lcd_sgdma_descriptor_write_translator:uav_writedata -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_address;                                        // lcd_sgdma_descriptor_write_translator:uav_address -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_lock;                                           // lcd_sgdma_descriptor_write_translator:uav_lock -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_write;                                          // lcd_sgdma_descriptor_write_translator:uav_write -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_read;                                           // lcd_sgdma_descriptor_write_translator:uav_read -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_readdata;                                       // lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> lcd_sgdma_descriptor_write_translator:uav_readdata
	wire          lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_debugaccess;                                    // lcd_sgdma_descriptor_write_translator:uav_debugaccess -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_byteenable;                                     // lcd_sgdma_descriptor_write_translator:uav_byteenable -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                                  // lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> lcd_sgdma_descriptor_write_translator:uav_readdatavalid
	wire          lcd_sgdma_m_read_translator_avalon_universal_master_0_waitrequest;                                              // lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_waitrequest -> lcd_sgdma_m_read_translator:uav_waitrequest
	wire    [3:0] lcd_sgdma_m_read_translator_avalon_universal_master_0_burstcount;                                               // lcd_sgdma_m_read_translator:uav_burstcount -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [63:0] lcd_sgdma_m_read_translator_avalon_universal_master_0_writedata;                                                // lcd_sgdma_m_read_translator:uav_writedata -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] lcd_sgdma_m_read_translator_avalon_universal_master_0_address;                                                  // lcd_sgdma_m_read_translator:uav_address -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_address
	wire          lcd_sgdma_m_read_translator_avalon_universal_master_0_lock;                                                     // lcd_sgdma_m_read_translator:uav_lock -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_lock
	wire          lcd_sgdma_m_read_translator_avalon_universal_master_0_write;                                                    // lcd_sgdma_m_read_translator:uav_write -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_write
	wire          lcd_sgdma_m_read_translator_avalon_universal_master_0_read;                                                     // lcd_sgdma_m_read_translator:uav_read -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_read
	wire   [63:0] lcd_sgdma_m_read_translator_avalon_universal_master_0_readdata;                                                 // lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_readdata -> lcd_sgdma_m_read_translator:uav_readdata
	wire          lcd_sgdma_m_read_translator_avalon_universal_master_0_debugaccess;                                              // lcd_sgdma_m_read_translator:uav_debugaccess -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [7:0] lcd_sgdma_m_read_translator_avalon_universal_master_0_byteenable;                                               // lcd_sgdma_m_read_translator:uav_byteenable -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          lcd_sgdma_m_read_translator_avalon_universal_master_0_readdatavalid;                                            // lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> lcd_sgdma_m_read_translator:uav_readdatavalid
	wire          sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest;                                      // sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> sdhc_ddr_clock_bridge_m0_translator:uav_waitrequest
	wire    [3:0] sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount;                                       // sdhc_ddr_clock_bridge_m0_translator:uav_burstcount -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [63:0] sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata;                                        // sdhc_ddr_clock_bridge_m0_translator:uav_writedata -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address;                                          // sdhc_ddr_clock_bridge_m0_translator:uav_address -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock;                                             // sdhc_ddr_clock_bridge_m0_translator:uav_lock -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write;                                            // sdhc_ddr_clock_bridge_m0_translator:uav_write -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read;                                             // sdhc_ddr_clock_bridge_m0_translator:uav_read -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [63:0] sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata;                                         // sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> sdhc_ddr_clock_bridge_m0_translator:uav_readdata
	wire          sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess;                                      // sdhc_ddr_clock_bridge_m0_translator:uav_debugaccess -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [7:0] sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable;                                       // sdhc_ddr_clock_bridge_m0_translator:uav_byteenable -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                                    // sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> sdhc_ddr_clock_bridge_m0_translator:uav_readdatavalid
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest;                                       // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_ddr_clock_bridge_m0_translator:uav_waitrequest
	wire    [2:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount;                                        // cpu_ddr_clock_bridge_m0_translator:uav_burstcount -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata;                                         // cpu_ddr_clock_bridge_m0_translator:uav_writedata -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address;                                           // cpu_ddr_clock_bridge_m0_translator:uav_address -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock;                                              // cpu_ddr_clock_bridge_m0_translator:uav_lock -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write;                                             // cpu_ddr_clock_bridge_m0_translator:uav_write -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read;                                              // cpu_ddr_clock_bridge_m0_translator:uav_read -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata;                                          // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> cpu_ddr_clock_bridge_m0_translator:uav_readdata
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess;                                       // cpu_ddr_clock_bridge_m0_translator:uav_debugaccess -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable;                                        // cpu_ddr_clock_bridge_m0_translator:uav_byteenable -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                                     // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_ddr_clock_bridge_m0_translator:uav_readdatavalid
	wire          tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest;                                       // tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> tse_ddr_clock_bridge_m0_translator:uav_waitrequest
	wire    [2:0] tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount;                                        // tse_ddr_clock_bridge_m0_translator:uav_burstcount -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata;                                         // tse_ddr_clock_bridge_m0_translator:uav_writedata -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address;                                           // tse_ddr_clock_bridge_m0_translator:uav_address -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock;                                              // tse_ddr_clock_bridge_m0_translator:uav_lock -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write;                                             // tse_ddr_clock_bridge_m0_translator:uav_write -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read;                                              // tse_ddr_clock_bridge_m0_translator:uav_read -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata;                                          // tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> tse_ddr_clock_bridge_m0_translator:uav_readdata
	wire          tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess;                                       // tse_ddr_clock_bridge_m0_translator:uav_debugaccess -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable;                                        // tse_ddr_clock_bridge_m0_translator:uav_byteenable -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                                     // tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> tse_ddr_clock_bridge_m0_translator:uav_readdatavalid
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                         // ddr2_sdram_s1_translator:uav_waitrequest -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [3:0] ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                          // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_sdram_s1_translator:uav_burstcount
	wire   [63:0] ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                           // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_sdram_s1_translator:uav_writedata
	wire   [31:0] ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                             // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_sdram_s1_translator:uav_address
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                               // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_sdram_s1_translator:uav_write
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_sdram_s1_translator:uav_lock
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_sdram_s1_translator:uav_read
	wire   [63:0] ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                            // ddr2_sdram_s1_translator:uav_readdata -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                       // ddr2_sdram_s1_translator:uav_readdatavalid -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                         // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_sdram_s1_translator:uav_debugaccess
	wire    [7:0] ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                          // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_sdram_s1_translator:uav_byteenable
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                  // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                        // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [125:0] ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                         // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                        // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                               // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                     // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                             // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [125:0] ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                      // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                     // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                   // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [63:0] ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                    // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                   // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                         // lcd_sgdma_csr_translator:uav_waitrequest -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                                          // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_sgdma_csr_translator:uav_burstcount
	wire   [31:0] lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                           // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_sgdma_csr_translator:uav_writedata
	wire   [31:0] lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_address;                                             // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_address -> lcd_sgdma_csr_translator:uav_address
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_write;                                               // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_write -> lcd_sgdma_csr_translator:uav_write
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                                // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_sgdma_csr_translator:uav_lock
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_read;                                                // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_read -> lcd_sgdma_csr_translator:uav_read
	wire   [31:0] lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                            // lcd_sgdma_csr_translator:uav_readdata -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                       // lcd_sgdma_csr_translator:uav_readdatavalid -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                         // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_sgdma_csr_translator:uav_debugaccess
	wire    [3:0] lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                                          // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_sgdma_csr_translator:uav_byteenable
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                  // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                                        // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                                         // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                                        // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                               // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                     // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                             // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                      // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                     // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                   // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                    // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                   // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sls_sdhc_read_master_translator_avalon_universal_master_0_waitrequest;                                          // sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_waitrequest -> sls_sdhc_read_master_translator:uav_waitrequest
	wire    [2:0] sls_sdhc_read_master_translator_avalon_universal_master_0_burstcount;                                           // sls_sdhc_read_master_translator:uav_burstcount -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sls_sdhc_read_master_translator_avalon_universal_master_0_writedata;                                            // sls_sdhc_read_master_translator:uav_writedata -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sls_sdhc_read_master_translator_avalon_universal_master_0_address;                                              // sls_sdhc_read_master_translator:uav_address -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_address
	wire          sls_sdhc_read_master_translator_avalon_universal_master_0_lock;                                                 // sls_sdhc_read_master_translator:uav_lock -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_lock
	wire          sls_sdhc_read_master_translator_avalon_universal_master_0_write;                                                // sls_sdhc_read_master_translator:uav_write -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_write
	wire          sls_sdhc_read_master_translator_avalon_universal_master_0_read;                                                 // sls_sdhc_read_master_translator:uav_read -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sls_sdhc_read_master_translator_avalon_universal_master_0_readdata;                                             // sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_readdata -> sls_sdhc_read_master_translator:uav_readdata
	wire          sls_sdhc_read_master_translator_avalon_universal_master_0_debugaccess;                                          // sls_sdhc_read_master_translator:uav_debugaccess -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sls_sdhc_read_master_translator_avalon_universal_master_0_byteenable;                                           // sls_sdhc_read_master_translator:uav_byteenable -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sls_sdhc_read_master_translator_avalon_universal_master_0_readdatavalid;                                        // sls_sdhc_read_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> sls_sdhc_read_master_translator:uav_readdatavalid
	wire          sls_sdhc_write_master_translator_avalon_universal_master_0_waitrequest;                                         // sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_waitrequest -> sls_sdhc_write_master_translator:uav_waitrequest
	wire    [2:0] sls_sdhc_write_master_translator_avalon_universal_master_0_burstcount;                                          // sls_sdhc_write_master_translator:uav_burstcount -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sls_sdhc_write_master_translator_avalon_universal_master_0_writedata;                                           // sls_sdhc_write_master_translator:uav_writedata -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sls_sdhc_write_master_translator_avalon_universal_master_0_address;                                             // sls_sdhc_write_master_translator:uav_address -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_address
	wire          sls_sdhc_write_master_translator_avalon_universal_master_0_lock;                                                // sls_sdhc_write_master_translator:uav_lock -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_lock
	wire          sls_sdhc_write_master_translator_avalon_universal_master_0_write;                                               // sls_sdhc_write_master_translator:uav_write -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_write
	wire          sls_sdhc_write_master_translator_avalon_universal_master_0_read;                                                // sls_sdhc_write_master_translator:uav_read -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sls_sdhc_write_master_translator_avalon_universal_master_0_readdata;                                            // sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_readdata -> sls_sdhc_write_master_translator:uav_readdata
	wire          sls_sdhc_write_master_translator_avalon_universal_master_0_debugaccess;                                         // sls_sdhc_write_master_translator:uav_debugaccess -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sls_sdhc_write_master_translator_avalon_universal_master_0_byteenable;                                          // sls_sdhc_write_master_translator:uav_byteenable -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sls_sdhc_write_master_translator_avalon_universal_master_0_readdatavalid;                                       // sls_sdhc_write_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> sls_sdhc_write_master_translator:uav_readdatavalid
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // sdhc_ddr_clock_bridge_s0_translator:uav_waitrequest -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [3:0] sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdhc_ddr_clock_bridge_s0_translator:uav_burstcount
	wire   [63:0] sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> sdhc_ddr_clock_bridge_s0_translator:uav_writedata
	wire   [31:0] sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                                  // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> sdhc_ddr_clock_bridge_s0_translator:uav_address
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                                    // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> sdhc_ddr_clock_bridge_s0_translator:uav_write
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                     // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> sdhc_ddr_clock_bridge_s0_translator:uav_lock
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                                     // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> sdhc_ddr_clock_bridge_s0_translator:uav_read
	wire   [63:0] sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // sdhc_ddr_clock_bridge_s0_translator:uav_readdata -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // sdhc_ddr_clock_bridge_s0_translator:uav_readdatavalid -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdhc_ddr_clock_bridge_s0_translator:uav_debugaccess
	wire    [7:0] sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdhc_ddr_clock_bridge_s0_translator:uav_byteenable
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [123:0] sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                              // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [123:0] sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [63:0] sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                        // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [63:0] sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                         // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                        // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest;                                     // cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_ddr_1_clock_bridge_m0_translator:uav_waitrequest
	wire    [2:0] cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_burstcount;                                      // cpu_ddr_1_clock_bridge_m0_translator:uav_burstcount -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_writedata;                                       // cpu_ddr_1_clock_bridge_m0_translator:uav_writedata -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_address;                                         // cpu_ddr_1_clock_bridge_m0_translator:uav_address -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_lock;                                            // cpu_ddr_1_clock_bridge_m0_translator:uav_lock -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_write;                                           // cpu_ddr_1_clock_bridge_m0_translator:uav_write -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_read;                                            // cpu_ddr_1_clock_bridge_m0_translator:uav_read -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_readdata;                                        // cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> cpu_ddr_1_clock_bridge_m0_translator:uav_readdata
	wire          cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess;                                     // cpu_ddr_1_clock_bridge_m0_translator:uav_debugaccess -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_byteenable;                                      // cpu_ddr_1_clock_bridge_m0_translator:uav_byteenable -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                                   // cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_ddr_1_clock_bridge_m0_translator:uav_readdatavalid
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // ddr2_sdram_1_s1_translator:uav_waitrequest -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [3:0] ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_sdram_1_s1_translator:uav_burstcount
	wire   [31:0] ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_sdram_1_s1_translator:uav_writedata
	wire   [25:0] ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_sdram_1_s1_translator:uav_address
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_sdram_1_s1_translator:uav_write
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_sdram_1_s1_translator:uav_lock
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_sdram_1_s1_translator:uav_read
	wire   [31:0] ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // ddr2_sdram_1_s1_translator:uav_readdata -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // ddr2_sdram_1_s1_translator:uav_readdatavalid -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_sdram_1_s1_translator:uav_debugaccess
	wire    [3:0] ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_sdram_1_s1_translator:uav_byteenable
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [79:0] ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [79:0] ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest;                                     // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> slow_peripheral_bridge_m0_translator:uav_waitrequest
	wire    [2:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount;                                      // slow_peripheral_bridge_m0_translator:uav_burstcount -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata;                                       // slow_peripheral_bridge_m0_translator:uav_writedata -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire    [9:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address;                                         // slow_peripheral_bridge_m0_translator:uav_address -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock;                                            // slow_peripheral_bridge_m0_translator:uav_lock -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write;                                           // slow_peripheral_bridge_m0_translator:uav_write -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read;                                            // slow_peripheral_bridge_m0_translator:uav_read -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata;                                        // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> slow_peripheral_bridge_m0_translator:uav_readdata
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess;                                     // slow_peripheral_bridge_m0_translator:uav_debugaccess -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable;                                      // slow_peripheral_bridge_m0_translator:uav_byteenable -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                                   // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> slow_peripheral_bridge_m0_translator:uav_readdatavalid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                         // button_pio_s1_translator:uav_waitrequest -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                          // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_pio_s1_translator:uav_burstcount
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                           // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_pio_s1_translator:uav_writedata
	wire    [9:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                             // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_pio_s1_translator:uav_address
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                               // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_pio_s1_translator:uav_write
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_pio_s1_translator:uav_lock
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_pio_s1_translator:uav_read
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                            // button_pio_s1_translator:uav_readdata -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                       // button_pio_s1_translator:uav_readdatavalid -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                         // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_pio_s1_translator:uav_debugaccess
	wire    [3:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                          // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_pio_s1_translator:uav_byteenable
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                         // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                               // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                             // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                      // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                   // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                    // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                   // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // high_res_timer_s1_translator:uav_waitrequest -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_res_timer_s1_translator:uav_burstcount
	wire   [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_res_timer_s1_translator:uav_writedata
	wire    [9:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_res_timer_s1_translator:uav_address
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_res_timer_s1_translator:uav_write
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_res_timer_s1_translator:uav_lock
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_res_timer_s1_translator:uav_read
	wire   [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // high_res_timer_s1_translator:uav_readdata -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // high_res_timer_s1_translator:uav_readdatavalid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_res_timer_s1_translator:uav_debugaccess
	wire    [3:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_res_timer_s1_translator:uav_byteenable
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire    [9:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                              // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                              // uart1_s1_translator:uav_waitrequest -> uart1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] uart1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                               // uart1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart1_s1_translator:uav_burstcount
	wire   [31:0] uart1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                // uart1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart1_s1_translator:uav_writedata
	wire    [9:0] uart1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                  // uart1_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart1_s1_translator:uav_address
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                    // uart1_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart1_s1_translator:uav_write
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                     // uart1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart1_s1_translator:uav_lock
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                     // uart1_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart1_s1_translator:uav_read
	wire   [31:0] uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                 // uart1_s1_translator:uav_readdata -> uart1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                            // uart1_s1_translator:uav_readdatavalid -> uart1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                              // uart1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart1_s1_translator:uav_debugaccess
	wire    [3:0] uart1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                               // uart1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart1_s1_translator:uav_byteenable
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                       // uart1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                             // uart1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                     // uart1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                              // uart1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                             // uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                    // uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                          // uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                  // uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                           // uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                          // uart1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                        // uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                         // uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                        // uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                            // led_pio_s1_translator:uav_waitrequest -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                             // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_pio_s1_translator:uav_burstcount
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                              // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_pio_s1_translator:uav_writedata
	wire    [9:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_pio_s1_translator:uav_address
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                  // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_pio_s1_translator:uav_write
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                   // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_pio_s1_translator:uav_lock
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                   // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_pio_s1_translator:uav_read
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                               // led_pio_s1_translator:uav_readdata -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                          // led_pio_s1_translator:uav_readdatavalid -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                            // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_pio_s1_translator:uav_debugaccess
	wire    [3:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                             // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_pio_s1_translator:uav_byteenable
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                           // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                   // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                            // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                           // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                  // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                        // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                         // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                        // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                      // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                       // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                      // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // performance_counter_control_slave_translator:uav_waitrequest -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> performance_counter_control_slave_translator:uav_burstcount
	wire   [31:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> performance_counter_control_slave_translator:uav_writedata
	wire    [9:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> performance_counter_control_slave_translator:uav_address
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> performance_counter_control_slave_translator:uav_write
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> performance_counter_control_slave_translator:uav_lock
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> performance_counter_control_slave_translator:uav_read
	wire   [31:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // performance_counter_control_slave_translator:uav_readdata -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // performance_counter_control_slave_translator:uav_readdatavalid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> performance_counter_control_slave_translator:uav_debugaccess
	wire    [3:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> performance_counter_control_slave_translator:uav_byteenable
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pll_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // pll_s1_translator:uav_waitrequest -> pll_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pll_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // pll_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pll_s1_translator:uav_burstcount
	wire   [31:0] pll_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // pll_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pll_s1_translator:uav_writedata
	wire    [9:0] pll_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // pll_s1_translator_avalon_universal_slave_0_agent:m0_address -> pll_s1_translator:uav_address
	wire          pll_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // pll_s1_translator_avalon_universal_slave_0_agent:m0_write -> pll_s1_translator:uav_write
	wire          pll_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // pll_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pll_s1_translator:uav_lock
	wire          pll_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // pll_s1_translator_avalon_universal_slave_0_agent:m0_read -> pll_s1_translator:uav_read
	wire   [31:0] pll_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // pll_s1_translator:uav_readdata -> pll_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pll_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // pll_s1_translator:uav_readdatavalid -> pll_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pll_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // pll_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pll_s1_translator:uav_debugaccess
	wire    [3:0] pll_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // pll_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pll_s1_translator:uav_byteenable
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // pll_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // pll_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // pll_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] pll_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // pll_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pll_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pll_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pll_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pll_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pll_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // pll_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // pll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // pll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                          // pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                           // pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                          // pll_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // sys_clk_timer_s1_translator:uav_waitrequest -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sys_clk_timer_s1_translator:uav_burstcount
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sys_clk_timer_s1_translator:uav_writedata
	wire    [9:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sys_clk_timer_s1_translator:uav_address
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sys_clk_timer_s1_translator:uav_write
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sys_clk_timer_s1_translator:uav_lock
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sys_clk_timer_s1_translator:uav_read
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // sys_clk_timer_s1_translator:uav_readdata -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // sys_clk_timer_s1_translator:uav_readdatavalid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sys_clk_timer_s1_translator:uav_debugaccess
	wire    [3:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sys_clk_timer_s1_translator:uav_byteenable
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire    [9:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                         // lcd_i2c_en_s1_translator:uav_waitrequest -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                          // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_i2c_en_s1_translator:uav_burstcount
	wire   [31:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                           // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_i2c_en_s1_translator:uav_writedata
	wire    [9:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_address;                                             // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_i2c_en_s1_translator:uav_address
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_write;                                               // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_i2c_en_s1_translator:uav_write
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_i2c_en_s1_translator:uav_lock
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_i2c_en_s1_translator:uav_read
	wire   [31:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                            // lcd_i2c_en_s1_translator:uav_readdata -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                       // lcd_i2c_en_s1_translator:uav_readdatavalid -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                         // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_i2c_en_s1_translator:uav_debugaccess
	wire    [3:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                          // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_i2c_en_s1_translator:uav_byteenable
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                  // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                        // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                         // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                        // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                               // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                     // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                             // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                      // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                     // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                   // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                    // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                   // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // lcd_i2c_scl_s1_translator:uav_waitrequest -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_i2c_scl_s1_translator:uav_burstcount
	wire   [31:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_i2c_scl_s1_translator:uav_writedata
	wire    [9:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address;                                            // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_i2c_scl_s1_translator:uav_address
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                              // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_i2c_scl_s1_translator:uav_write
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                               // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_i2c_scl_s1_translator:uav_lock
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                               // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_i2c_scl_s1_translator:uav_read
	wire   [31:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // lcd_i2c_scl_s1_translator:uav_readdata -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // lcd_i2c_scl_s1_translator:uav_readdatavalid -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_i2c_scl_s1_translator:uav_debugaccess
	wire    [3:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_i2c_scl_s1_translator:uav_byteenable
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // lcd_i2c_sdat_s1_translator:uav_waitrequest -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_i2c_sdat_s1_translator:uav_burstcount
	wire   [31:0] lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_i2c_sdat_s1_translator:uav_writedata
	wire    [9:0] lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_i2c_sdat_s1_translator:uav_address
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_i2c_sdat_s1_translator:uav_write
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_i2c_sdat_s1_translator:uav_lock
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_i2c_sdat_s1_translator:uav_read
	wire   [31:0] lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // lcd_i2c_sdat_s1_translator:uav_readdata -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // lcd_i2c_sdat_s1_translator:uav_readdatavalid -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_i2c_sdat_s1_translator:uav_debugaccess
	wire    [3:0] lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_i2c_sdat_s1_translator:uav_byteenable
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // pio_id_eeprom_dat_s1_translator:uav_waitrequest -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_id_eeprom_dat_s1_translator:uav_burstcount
	wire   [31:0] pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_id_eeprom_dat_s1_translator:uav_writedata
	wire    [9:0] pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_id_eeprom_dat_s1_translator:uav_address
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_id_eeprom_dat_s1_translator:uav_write
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_id_eeprom_dat_s1_translator:uav_lock
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_id_eeprom_dat_s1_translator:uav_read
	wire   [31:0] pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // pio_id_eeprom_dat_s1_translator:uav_readdata -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // pio_id_eeprom_dat_s1_translator:uav_readdatavalid -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_id_eeprom_dat_s1_translator:uav_debugaccess
	wire    [3:0] pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_id_eeprom_dat_s1_translator:uav_byteenable
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // pio_id_eeprom_scl_s1_translator:uav_waitrequest -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_id_eeprom_scl_s1_translator:uav_burstcount
	wire   [31:0] pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_id_eeprom_scl_s1_translator:uav_writedata
	wire    [9:0] pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_id_eeprom_scl_s1_translator:uav_address
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_id_eeprom_scl_s1_translator:uav_write
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_id_eeprom_scl_s1_translator:uav_lock
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_id_eeprom_scl_s1_translator:uav_read
	wire   [31:0] pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // pio_id_eeprom_scl_s1_translator:uav_readdata -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // pio_id_eeprom_scl_s1_translator:uav_readdatavalid -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_id_eeprom_scl_s1_translator:uav_debugaccess
	wire    [3:0] pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_id_eeprom_scl_s1_translator:uav_byteenable
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // touch_panel_pen_irq_n_s1_translator:uav_waitrequest -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> touch_panel_pen_irq_n_s1_translator:uav_burstcount
	wire   [31:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> touch_panel_pen_irq_n_s1_translator:uav_writedata
	wire    [9:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_address -> touch_panel_pen_irq_n_s1_translator:uav_address
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_write -> touch_panel_pen_irq_n_s1_translator:uav_write
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_lock -> touch_panel_pen_irq_n_s1_translator:uav_lock
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_read -> touch_panel_pen_irq_n_s1_translator:uav_read
	wire   [31:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // touch_panel_pen_irq_n_s1_translator:uav_readdata -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // touch_panel_pen_irq_n_s1_translator:uav_readdatavalid -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> touch_panel_pen_irq_n_s1_translator:uav_debugaccess
	wire    [3:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> touch_panel_pen_irq_n_s1_translator:uav_byteenable
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // touch_panel_spi_spi_control_port_translator:uav_waitrequest -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> touch_panel_spi_spi_control_port_translator:uav_burstcount
	wire   [31:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                        // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> touch_panel_spi_spi_control_port_translator:uav_writedata
	wire    [9:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address;                          // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> touch_panel_spi_spi_control_port_translator:uav_address
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write;                            // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> touch_panel_spi_spi_control_port_translator:uav_write
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                             // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> touch_panel_spi_spi_control_port_translator:uav_lock
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read;                             // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> touch_panel_spi_spi_control_port_translator:uav_read
	wire   [31:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                         // touch_panel_spi_spi_control_port_translator:uav_readdata -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // touch_panel_spi_spi_control_port_translator:uav_readdatavalid -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> touch_panel_spi_spi_control_port_translator:uav_debugaccess
	wire    [3:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> touch_panel_spi_spi_control_port_translator:uav_byteenable
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [69:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                      // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [69:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest;                                              // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_m_write_translator:uav_waitrequest
	wire    [2:0] sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount;                                               // sgdma_rx_m_write_translator:uav_burstcount -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_writedata;                                                // sgdma_rx_m_write_translator:uav_writedata -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_address;                                                  // sgdma_rx_m_write_translator:uav_address -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_lock;                                                     // sgdma_rx_m_write_translator:uav_lock -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_write;                                                    // sgdma_rx_m_write_translator:uav_write -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_read;                                                     // sgdma_rx_m_write_translator:uav_read -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_readdata;                                                 // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_m_write_translator:uav_readdata
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess;                                              // sgdma_rx_m_write_translator:uav_debugaccess -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable;                                               // sgdma_rx_m_write_translator:uav_byteenable -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid;                                            // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_m_write_translator:uav_readdatavalid
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest;                                               // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_m_read_translator:uav_waitrequest
	wire    [2:0] sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount;                                                // sgdma_tx_m_read_translator:uav_burstcount -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_writedata;                                                 // sgdma_tx_m_read_translator:uav_writedata -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_address;                                                   // sgdma_tx_m_read_translator:uav_address -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_lock;                                                      // sgdma_tx_m_read_translator:uav_lock -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_write;                                                     // sgdma_tx_m_read_translator:uav_write -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_read;                                                      // sgdma_tx_m_read_translator:uav_read -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_readdata;                                                  // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_m_read_translator:uav_readdata
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess;                                               // sgdma_tx_m_read_translator:uav_debugaccess -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable;                                                // sgdma_tx_m_read_translator:uav_byteenable -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid;                                             // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_m_read_translator:uav_readdatavalid
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // tse_ddr_clock_bridge_s0_translator:uav_waitrequest -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> tse_ddr_clock_bridge_s0_translator:uav_burstcount
	wire   [31:0] tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> tse_ddr_clock_bridge_s0_translator:uav_writedata
	wire   [31:0] tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                                   // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> tse_ddr_clock_bridge_s0_translator:uav_address
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                                     // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> tse_ddr_clock_bridge_s0_translator:uav_write
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                      // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> tse_ddr_clock_bridge_s0_translator:uav_lock
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                                      // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> tse_ddr_clock_bridge_s0_translator:uav_read
	wire   [31:0] tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // tse_ddr_clock_bridge_s0_translator:uav_readdata -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // tse_ddr_clock_bridge_s0_translator:uav_readdatavalid -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> tse_ddr_clock_bridge_s0_translator:uav_debugaccess
	wire    [3:0] tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> tse_ddr_clock_bridge_s0_translator:uav_byteenable
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                               // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_waitrequest;                     // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> pipeline_bridge_before_tristate_bridge_m0_translator:uav_waitrequest
	wire    [2:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_burstcount;                      // pipeline_bridge_before_tristate_bridge_m0_translator:uav_burstcount -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_writedata;                       // pipeline_bridge_before_tristate_bridge_m0_translator:uav_writedata -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [26:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_address;                         // pipeline_bridge_before_tristate_bridge_m0_translator:uav_address -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_lock;                            // pipeline_bridge_before_tristate_bridge_m0_translator:uav_lock -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_write;                           // pipeline_bridge_before_tristate_bridge_m0_translator:uav_write -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_read;                            // pipeline_bridge_before_tristate_bridge_m0_translator:uav_read -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdata;                        // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> pipeline_bridge_before_tristate_bridge_m0_translator:uav_readdata
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_debugaccess;                     // pipeline_bridge_before_tristate_bridge_m0_translator:uav_debugaccess -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_byteenable;                      // pipeline_bridge_before_tristate_bridge_m0_translator:uav_byteenable -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                   // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> pipeline_bridge_before_tristate_bridge_m0_translator:uav_readdatavalid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                         // ext_flash_uas_translator:uav_waitrequest -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                          // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> ext_flash_uas_translator:uav_burstcount
	wire   [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                           // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> ext_flash_uas_translator:uav_writedata
	wire   [26:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address;                                             // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_address -> ext_flash_uas_translator:uav_address
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write;                                               // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_write -> ext_flash_uas_translator:uav_write
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                                // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_lock -> ext_flash_uas_translator:uav_lock
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read;                                                // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_read -> ext_flash_uas_translator:uav_read
	wire   [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                            // ext_flash_uas_translator:uav_readdata -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                       // ext_flash_uas_translator:uav_readdatavalid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                         // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ext_flash_uas_translator:uav_debugaccess
	wire    [1:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                          // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> ext_flash_uas_translator:uav_byteenable
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                  // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                                        // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [62:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                                         // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                                        // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                               // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                     // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                             // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [62:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                      // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                     // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                   // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                    // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                   // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          max2_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                              // max2_uas_translator:uav_waitrequest -> max2_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] max2_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                               // max2_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> max2_uas_translator:uav_burstcount
	wire   [31:0] max2_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                                // max2_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> max2_uas_translator:uav_writedata
	wire   [26:0] max2_uas_translator_avalon_universal_slave_0_agent_m0_address;                                                  // max2_uas_translator_avalon_universal_slave_0_agent:m0_address -> max2_uas_translator:uav_address
	wire          max2_uas_translator_avalon_universal_slave_0_agent_m0_write;                                                    // max2_uas_translator_avalon_universal_slave_0_agent:m0_write -> max2_uas_translator:uav_write
	wire          max2_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                                     // max2_uas_translator_avalon_universal_slave_0_agent:m0_lock -> max2_uas_translator:uav_lock
	wire          max2_uas_translator_avalon_universal_slave_0_agent_m0_read;                                                     // max2_uas_translator_avalon_universal_slave_0_agent:m0_read -> max2_uas_translator:uav_read
	wire   [31:0] max2_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                                 // max2_uas_translator:uav_readdata -> max2_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          max2_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                            // max2_uas_translator:uav_readdatavalid -> max2_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          max2_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                              // max2_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> max2_uas_translator:uav_debugaccess
	wire    [3:0] max2_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                               // max2_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> max2_uas_translator:uav_byteenable
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                       // max2_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                                             // max2_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                     // max2_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [80:0] max2_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                                              // max2_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                                             // max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> max2_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                    // max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> max2_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                          // max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> max2_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                  // max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> max2_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [80:0] max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                           // max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> max2_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                          // max2_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                        // max2_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> max2_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] max2_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                         // max2_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> max2_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                        // max2_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> max2_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                      // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                            // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                    // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire   [88:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                             // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                            // addr_router:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                               // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                     // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                             // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire   [88:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                      // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                     // addr_router_001:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                             // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                                   // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                           // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [88:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                                    // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                                   // addr_router_002:sink_ready -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                                  // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire   [88:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                                   // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router_003:sink_ready -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                             // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                                   // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                           // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire   [88:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                                    // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                                   // addr_router_004:sink_ready -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                                  // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire   [88:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                                   // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router_005:sink_ready -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire   [88:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [88:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_001:sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                                // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [88:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data;                                                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_002:sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                                // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire   [88:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data;                                                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_003:sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                                        // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire   [88:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data;                                         // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_004:sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_valid;                                            // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire   [88:0] sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_data;                                             // sls_sdhc_control_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_005:sink_ready -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                   // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [88:0] pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                    // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_006:sink_ready -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                     // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [88:0] cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                                      // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_007:sink_ready -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                   // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [88:0] cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                                    // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_008:sink_ready -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                   // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire   [88:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                                    // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_009:sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	wire          lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                                  // lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	wire          lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	wire   [88:0] lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                                   // lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	wire          lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router_006:sink_ready -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                           // lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_007:sink_endofpacket
	wire          lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                                 // lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_007:sink_valid
	wire          lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                         // lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_007:sink_startofpacket
	wire   [88:0] lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                                  // lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_007:sink_data
	wire          lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                                 // addr_router_007:sink_ready -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                                     // lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_008:sink_endofpacket
	wire          lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_valid;                                           // lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_008:sink_valid
	wire          lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                                   // lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_008:sink_startofpacket
	wire  [124:0] lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_data;                                            // lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_008:sink_data
	wire          lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_ready;                                           // addr_router_008:sink_ready -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                             // sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_009:sink_endofpacket
	wire          sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                                   // sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_009:sink_valid
	wire          sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                           // sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_009:sink_startofpacket
	wire  [124:0] sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                                    // sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_009:sink_data
	wire          sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                                   // addr_router_009:sink_ready -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                              // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_010:sink_endofpacket
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                                    // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_010:sink_valid
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                            // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_010:sink_startofpacket
	wire   [88:0] cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                                     // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_010:sink_data
	wire          cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                                    // addr_router_010:sink_ready -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                              // tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_011:sink_endofpacket
	wire          tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                                    // tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_011:sink_valid
	wire          tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                            // tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_011:sink_startofpacket
	wire   [88:0] tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                                     // tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_011:sink_data
	wire          tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                                    // addr_router_011:sink_ready -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                         // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                               // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                       // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [124:0] ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                               // id_router_010:sink_ready -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                         // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                               // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                       // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire   [88:0] lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_data;                                                // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                               // id_router_011:sink_ready -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                 // sls_sdhc_read_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_012:sink_endofpacket
	wire          sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_valid;                                       // sls_sdhc_read_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_012:sink_valid
	wire          sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                               // sls_sdhc_read_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_012:sink_startofpacket
	wire   [86:0] sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_data;                                        // sls_sdhc_read_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_012:sink_data
	wire          sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_ready;                                       // addr_router_012:sink_ready -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                // sls_sdhc_write_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_013:sink_endofpacket
	wire          sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_valid;                                      // sls_sdhc_write_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_013:sink_valid
	wire          sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                              // sls_sdhc_write_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_013:sink_startofpacket
	wire   [86:0] sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_data;                                       // sls_sdhc_write_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_013:sink_data
	wire          sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_ready;                                      // addr_router_013:sink_ready -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                    // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [122:0] sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                                     // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_012:sink_ready -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_014:sink_endofpacket
	wire          cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                                  // cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_014:sink_valid
	wire          cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_014:sink_startofpacket
	wire   [78:0] cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                                   // cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_014:sink_data
	wire          cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router_014:sink_ready -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire   [78:0] ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_013:sink_ready -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_015:sink_endofpacket
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                                  // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_015:sink_valid
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_015:sink_startofpacket
	wire   [68:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                                   // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_015:sink_data
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router_015:sink_ready -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                         // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                               // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                       // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire   [68:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                               // id_router_014:sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire   [68:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_015:sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire   [68:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_016:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                              // uart1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                    // uart1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                            // uart1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire   [68:0] uart1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                     // uart1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                    // id_router_017:sink_ready -> uart1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                            // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                  // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                          // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire   [68:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                   // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                  // id_router_018:sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire   [68:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_019:sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // pll_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // pll_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // pll_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire   [68:0] pll_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // pll_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          pll_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_020:sink_ready -> pll_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire   [68:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_021:sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire   [68:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_022:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                         // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                               // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                       // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire   [68:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                               // id_router_023:sink_ready -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                              // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire   [68:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                               // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_024:sink_ready -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire   [68:0] lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire          lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_025:sink_ready -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire   [68:0] pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire          pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_026:sink_ready -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire   [68:0] pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire          pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_027:sink_ready -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire   [68:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_028:sink_ready -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                            // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	wire   [68:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data;                             // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_029:sink_ready -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                                     // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_016:sink_endofpacket
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid;                                           // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_016:sink_valid
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                                   // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_016:sink_startofpacket
	wire   [84:0] sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data;                                            // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_016:sink_data
	wire          sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready;                                           // addr_router_016:sink_ready -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                                      // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_017:sink_endofpacket
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid;                                            // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_017:sink_valid
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                                    // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_017:sink_startofpacket
	wire   [84:0] sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data;                                             // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_017:sink_data
	wire          sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready;                                            // addr_router_017:sink_ready -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                     // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	wire   [84:0] tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                                      // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	wire          tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_030:sink_ready -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;            // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_018:sink_endofpacket
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                  // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_018:sink_valid
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;          // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_018:sink_startofpacket
	wire   [79:0] pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                   // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_018:sink_data
	wire          pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                  // addr_router_018:sink_ready -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                         // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_031:sink_endofpacket
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                               // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_031:sink_valid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                       // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_031:sink_startofpacket
	wire   [61:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data;                                                // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_031:sink_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                               // id_router_031:sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                              // max2_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_032:sink_endofpacket
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                                    // max2_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_032:sink_valid
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                            // max2_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_032:sink_startofpacket
	wire   [79:0] max2_uas_translator_avalon_universal_slave_0_agent_rp_data;                                                     // max2_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_032:sink_data
	wire          max2_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                                    // id_router_032:sink_ready -> max2_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                                    // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                          // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                                  // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire   [88:0] addr_router_src_data;                                                                                           // addr_router:src_data -> limiter:cmd_sink_data
	wire    [9:0] addr_router_src_channel;                                                                                        // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                          // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                                    // limiter:rsp_src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                          // limiter:rsp_src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                                  // limiter:rsp_src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] limiter_rsp_src_data;                                                                                           // limiter:rsp_src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [9:0] limiter_rsp_src_channel;                                                                                        // limiter:rsp_src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                          // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                                // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                      // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                              // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire   [88:0] addr_router_001_src_data;                                                                                       // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire    [9:0] addr_router_001_src_channel;                                                                                    // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                                      // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                                // limiter_001:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                                      // limiter_001:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                              // limiter_001:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] limiter_001_rsp_src_data;                                                                                       // limiter_001:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [9:0] limiter_001_rsp_src_channel;                                                                                    // limiter_001:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                                      // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          addr_router_002_src_endofpacket;                                                                                // addr_router_002:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                      // addr_router_002:src_valid -> limiter_002:cmd_sink_valid
	wire          addr_router_002_src_startofpacket;                                                                              // addr_router_002:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire   [88:0] addr_router_002_src_data;                                                                                       // addr_router_002:src_data -> limiter_002:cmd_sink_data
	wire    [9:0] addr_router_002_src_channel;                                                                                    // addr_router_002:src_channel -> limiter_002:cmd_sink_channel
	wire          addr_router_002_src_ready;                                                                                      // limiter_002:cmd_sink_ready -> addr_router_002:src_ready
	wire          limiter_002_rsp_src_endofpacket;                                                                                // limiter_002:rsp_src_endofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_002_rsp_src_valid;                                                                                      // limiter_002:rsp_src_valid -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_002_rsp_src_startofpacket;                                                                              // limiter_002:rsp_src_startofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] limiter_002_rsp_src_data;                                                                                       // limiter_002:rsp_src_data -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire    [9:0] limiter_002_rsp_src_channel;                                                                                    // limiter_002:rsp_src_channel -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_002_rsp_src_ready;                                                                                      // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire          addr_router_003_src_endofpacket;                                                                                // addr_router_003:src_endofpacket -> limiter_003:cmd_sink_endofpacket
	wire          addr_router_003_src_valid;                                                                                      // addr_router_003:src_valid -> limiter_003:cmd_sink_valid
	wire          addr_router_003_src_startofpacket;                                                                              // addr_router_003:src_startofpacket -> limiter_003:cmd_sink_startofpacket
	wire   [88:0] addr_router_003_src_data;                                                                                       // addr_router_003:src_data -> limiter_003:cmd_sink_data
	wire    [9:0] addr_router_003_src_channel;                                                                                    // addr_router_003:src_channel -> limiter_003:cmd_sink_channel
	wire          addr_router_003_src_ready;                                                                                      // limiter_003:cmd_sink_ready -> addr_router_003:src_ready
	wire          limiter_003_rsp_src_endofpacket;                                                                                // limiter_003:rsp_src_endofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_003_rsp_src_valid;                                                                                      // limiter_003:rsp_src_valid -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_003_rsp_src_startofpacket;                                                                              // limiter_003:rsp_src_startofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] limiter_003_rsp_src_data;                                                                                       // limiter_003:rsp_src_data -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire    [9:0] limiter_003_rsp_src_channel;                                                                                    // limiter_003:rsp_src_channel -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_003_rsp_src_ready;                                                                                      // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> limiter_003:rsp_src_ready
	wire          addr_router_004_src_endofpacket;                                                                                // addr_router_004:src_endofpacket -> limiter_004:cmd_sink_endofpacket
	wire          addr_router_004_src_valid;                                                                                      // addr_router_004:src_valid -> limiter_004:cmd_sink_valid
	wire          addr_router_004_src_startofpacket;                                                                              // addr_router_004:src_startofpacket -> limiter_004:cmd_sink_startofpacket
	wire   [88:0] addr_router_004_src_data;                                                                                       // addr_router_004:src_data -> limiter_004:cmd_sink_data
	wire    [9:0] addr_router_004_src_channel;                                                                                    // addr_router_004:src_channel -> limiter_004:cmd_sink_channel
	wire          addr_router_004_src_ready;                                                                                      // limiter_004:cmd_sink_ready -> addr_router_004:src_ready
	wire          limiter_004_rsp_src_endofpacket;                                                                                // limiter_004:rsp_src_endofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_004_rsp_src_valid;                                                                                      // limiter_004:rsp_src_valid -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_004_rsp_src_startofpacket;                                                                              // limiter_004:rsp_src_startofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] limiter_004_rsp_src_data;                                                                                       // limiter_004:rsp_src_data -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire    [9:0] limiter_004_rsp_src_channel;                                                                                    // limiter_004:rsp_src_channel -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_004_rsp_src_ready;                                                                                      // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> limiter_004:rsp_src_ready
	wire          addr_router_005_src_endofpacket;                                                                                // addr_router_005:src_endofpacket -> limiter_005:cmd_sink_endofpacket
	wire          addr_router_005_src_valid;                                                                                      // addr_router_005:src_valid -> limiter_005:cmd_sink_valid
	wire          addr_router_005_src_startofpacket;                                                                              // addr_router_005:src_startofpacket -> limiter_005:cmd_sink_startofpacket
	wire   [88:0] addr_router_005_src_data;                                                                                       // addr_router_005:src_data -> limiter_005:cmd_sink_data
	wire    [9:0] addr_router_005_src_channel;                                                                                    // addr_router_005:src_channel -> limiter_005:cmd_sink_channel
	wire          addr_router_005_src_ready;                                                                                      // limiter_005:cmd_sink_ready -> addr_router_005:src_ready
	wire          limiter_005_rsp_src_endofpacket;                                                                                // limiter_005:rsp_src_endofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_005_rsp_src_valid;                                                                                      // limiter_005:rsp_src_valid -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_005_rsp_src_startofpacket;                                                                              // limiter_005:rsp_src_startofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] limiter_005_rsp_src_data;                                                                                       // limiter_005:rsp_src_data -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire    [9:0] limiter_005_rsp_src_channel;                                                                                    // limiter_005:rsp_src_channel -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_005_rsp_src_ready;                                                                                      // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> limiter_005:rsp_src_ready
	wire          addr_router_006_src_endofpacket;                                                                                // addr_router_006:src_endofpacket -> limiter_006:cmd_sink_endofpacket
	wire          addr_router_006_src_valid;                                                                                      // addr_router_006:src_valid -> limiter_006:cmd_sink_valid
	wire          addr_router_006_src_startofpacket;                                                                              // addr_router_006:src_startofpacket -> limiter_006:cmd_sink_startofpacket
	wire   [88:0] addr_router_006_src_data;                                                                                       // addr_router_006:src_data -> limiter_006:cmd_sink_data
	wire    [5:0] addr_router_006_src_channel;                                                                                    // addr_router_006:src_channel -> limiter_006:cmd_sink_channel
	wire          addr_router_006_src_ready;                                                                                      // limiter_006:cmd_sink_ready -> addr_router_006:src_ready
	wire          limiter_006_rsp_src_endofpacket;                                                                                // limiter_006:rsp_src_endofpacket -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_006_rsp_src_valid;                                                                                      // limiter_006:rsp_src_valid -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_006_rsp_src_startofpacket;                                                                              // limiter_006:rsp_src_startofpacket -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] limiter_006_rsp_src_data;                                                                                       // limiter_006:rsp_src_data -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_006_rsp_src_channel;                                                                                    // limiter_006:rsp_src_channel -> lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_006_rsp_src_ready;                                                                                      // lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> limiter_006:rsp_src_ready
	wire          addr_router_007_src_endofpacket;                                                                                // addr_router_007:src_endofpacket -> limiter_007:cmd_sink_endofpacket
	wire          addr_router_007_src_valid;                                                                                      // addr_router_007:src_valid -> limiter_007:cmd_sink_valid
	wire          addr_router_007_src_startofpacket;                                                                              // addr_router_007:src_startofpacket -> limiter_007:cmd_sink_startofpacket
	wire   [88:0] addr_router_007_src_data;                                                                                       // addr_router_007:src_data -> limiter_007:cmd_sink_data
	wire    [5:0] addr_router_007_src_channel;                                                                                    // addr_router_007:src_channel -> limiter_007:cmd_sink_channel
	wire          addr_router_007_src_ready;                                                                                      // limiter_007:cmd_sink_ready -> addr_router_007:src_ready
	wire          limiter_007_rsp_src_endofpacket;                                                                                // limiter_007:rsp_src_endofpacket -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_007_rsp_src_valid;                                                                                      // limiter_007:rsp_src_valid -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_007_rsp_src_startofpacket;                                                                              // limiter_007:rsp_src_startofpacket -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] limiter_007_rsp_src_data;                                                                                       // limiter_007:rsp_src_data -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_007_rsp_src_channel;                                                                                    // limiter_007:rsp_src_channel -> lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_007_rsp_src_ready;                                                                                      // lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> limiter_007:rsp_src_ready
	wire          addr_router_008_src_endofpacket;                                                                                // addr_router_008:src_endofpacket -> limiter_008:cmd_sink_endofpacket
	wire          addr_router_008_src_valid;                                                                                      // addr_router_008:src_valid -> limiter_008:cmd_sink_valid
	wire          addr_router_008_src_startofpacket;                                                                              // addr_router_008:src_startofpacket -> limiter_008:cmd_sink_startofpacket
	wire  [124:0] addr_router_008_src_data;                                                                                       // addr_router_008:src_data -> limiter_008:cmd_sink_data
	wire    [5:0] addr_router_008_src_channel;                                                                                    // addr_router_008:src_channel -> limiter_008:cmd_sink_channel
	wire          addr_router_008_src_ready;                                                                                      // limiter_008:cmd_sink_ready -> addr_router_008:src_ready
	wire          limiter_008_rsp_src_endofpacket;                                                                                // limiter_008:rsp_src_endofpacket -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_008_rsp_src_valid;                                                                                      // limiter_008:rsp_src_valid -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_008_rsp_src_startofpacket;                                                                              // limiter_008:rsp_src_startofpacket -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [124:0] limiter_008_rsp_src_data;                                                                                       // limiter_008:rsp_src_data -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_008_rsp_src_channel;                                                                                    // limiter_008:rsp_src_channel -> lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_008_rsp_src_ready;                                                                                      // lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:rp_ready -> limiter_008:rsp_src_ready
	wire          addr_router_009_src_endofpacket;                                                                                // addr_router_009:src_endofpacket -> limiter_009:cmd_sink_endofpacket
	wire          addr_router_009_src_valid;                                                                                      // addr_router_009:src_valid -> limiter_009:cmd_sink_valid
	wire          addr_router_009_src_startofpacket;                                                                              // addr_router_009:src_startofpacket -> limiter_009:cmd_sink_startofpacket
	wire  [124:0] addr_router_009_src_data;                                                                                       // addr_router_009:src_data -> limiter_009:cmd_sink_data
	wire    [5:0] addr_router_009_src_channel;                                                                                    // addr_router_009:src_channel -> limiter_009:cmd_sink_channel
	wire          addr_router_009_src_ready;                                                                                      // limiter_009:cmd_sink_ready -> addr_router_009:src_ready
	wire          limiter_009_rsp_src_endofpacket;                                                                                // limiter_009:rsp_src_endofpacket -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_009_rsp_src_valid;                                                                                      // limiter_009:rsp_src_valid -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_009_rsp_src_startofpacket;                                                                              // limiter_009:rsp_src_startofpacket -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [124:0] limiter_009_rsp_src_data;                                                                                       // limiter_009:rsp_src_data -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_009_rsp_src_channel;                                                                                    // limiter_009:rsp_src_channel -> sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_009_rsp_src_ready;                                                                                      // sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_009:rsp_src_ready
	wire          addr_router_010_src_endofpacket;                                                                                // addr_router_010:src_endofpacket -> limiter_010:cmd_sink_endofpacket
	wire          addr_router_010_src_valid;                                                                                      // addr_router_010:src_valid -> limiter_010:cmd_sink_valid
	wire          addr_router_010_src_startofpacket;                                                                              // addr_router_010:src_startofpacket -> limiter_010:cmd_sink_startofpacket
	wire   [88:0] addr_router_010_src_data;                                                                                       // addr_router_010:src_data -> limiter_010:cmd_sink_data
	wire    [5:0] addr_router_010_src_channel;                                                                                    // addr_router_010:src_channel -> limiter_010:cmd_sink_channel
	wire          addr_router_010_src_ready;                                                                                      // limiter_010:cmd_sink_ready -> addr_router_010:src_ready
	wire          limiter_010_rsp_src_endofpacket;                                                                                // limiter_010:rsp_src_endofpacket -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_010_rsp_src_valid;                                                                                      // limiter_010:rsp_src_valid -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_010_rsp_src_startofpacket;                                                                              // limiter_010:rsp_src_startofpacket -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] limiter_010_rsp_src_data;                                                                                       // limiter_010:rsp_src_data -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_010_rsp_src_channel;                                                                                    // limiter_010:rsp_src_channel -> cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_010_rsp_src_ready;                                                                                      // cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_010:rsp_src_ready
	wire          addr_router_011_src_endofpacket;                                                                                // addr_router_011:src_endofpacket -> limiter_011:cmd_sink_endofpacket
	wire          addr_router_011_src_valid;                                                                                      // addr_router_011:src_valid -> limiter_011:cmd_sink_valid
	wire          addr_router_011_src_startofpacket;                                                                              // addr_router_011:src_startofpacket -> limiter_011:cmd_sink_startofpacket
	wire   [88:0] addr_router_011_src_data;                                                                                       // addr_router_011:src_data -> limiter_011:cmd_sink_data
	wire    [5:0] addr_router_011_src_channel;                                                                                    // addr_router_011:src_channel -> limiter_011:cmd_sink_channel
	wire          addr_router_011_src_ready;                                                                                      // limiter_011:cmd_sink_ready -> addr_router_011:src_ready
	wire          limiter_011_rsp_src_endofpacket;                                                                                // limiter_011:rsp_src_endofpacket -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_011_rsp_src_valid;                                                                                      // limiter_011:rsp_src_valid -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_011_rsp_src_startofpacket;                                                                              // limiter_011:rsp_src_startofpacket -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] limiter_011_rsp_src_data;                                                                                       // limiter_011:rsp_src_data -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_011_rsp_src_channel;                                                                                    // limiter_011:rsp_src_channel -> tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_011_rsp_src_ready;                                                                                      // tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_011:rsp_src_ready
	wire          addr_router_015_src_endofpacket;                                                                                // addr_router_015:src_endofpacket -> limiter_012:cmd_sink_endofpacket
	wire          addr_router_015_src_valid;                                                                                      // addr_router_015:src_valid -> limiter_012:cmd_sink_valid
	wire          addr_router_015_src_startofpacket;                                                                              // addr_router_015:src_startofpacket -> limiter_012:cmd_sink_startofpacket
	wire   [68:0] addr_router_015_src_data;                                                                                       // addr_router_015:src_data -> limiter_012:cmd_sink_data
	wire   [15:0] addr_router_015_src_channel;                                                                                    // addr_router_015:src_channel -> limiter_012:cmd_sink_channel
	wire          addr_router_015_src_ready;                                                                                      // limiter_012:cmd_sink_ready -> addr_router_015:src_ready
	wire          limiter_012_rsp_src_endofpacket;                                                                                // limiter_012:rsp_src_endofpacket -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_012_rsp_src_valid;                                                                                      // limiter_012:rsp_src_valid -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_012_rsp_src_startofpacket;                                                                              // limiter_012:rsp_src_startofpacket -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [68:0] limiter_012_rsp_src_data;                                                                                       // limiter_012:rsp_src_data -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] limiter_012_rsp_src_channel;                                                                                    // limiter_012:rsp_src_channel -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_012_rsp_src_ready;                                                                                      // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_012:rsp_src_ready
	wire          addr_router_018_src_endofpacket;                                                                                // addr_router_018:src_endofpacket -> limiter_013:cmd_sink_endofpacket
	wire          addr_router_018_src_valid;                                                                                      // addr_router_018:src_valid -> limiter_013:cmd_sink_valid
	wire          addr_router_018_src_startofpacket;                                                                              // addr_router_018:src_startofpacket -> limiter_013:cmd_sink_startofpacket
	wire   [79:0] addr_router_018_src_data;                                                                                       // addr_router_018:src_data -> limiter_013:cmd_sink_data
	wire    [1:0] addr_router_018_src_channel;                                                                                    // addr_router_018:src_channel -> limiter_013:cmd_sink_channel
	wire          addr_router_018_src_ready;                                                                                      // limiter_013:cmd_sink_ready -> addr_router_018:src_ready
	wire          limiter_013_rsp_src_endofpacket;                                                                                // limiter_013:rsp_src_endofpacket -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_013_rsp_src_valid;                                                                                      // limiter_013:rsp_src_valid -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_013_rsp_src_startofpacket;                                                                              // limiter_013:rsp_src_startofpacket -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [79:0] limiter_013_rsp_src_data;                                                                                       // limiter_013:rsp_src_data -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] limiter_013_rsp_src_channel;                                                                                    // limiter_013:rsp_src_channel -> pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_013_rsp_src_ready;                                                                                      // pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_013:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                              // burst_adapter:source0_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                    // burst_adapter:source0_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                            // burst_adapter:source0_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [61:0] burst_adapter_source0_data;                                                                                     // burst_adapter:source0_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                    // ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [1:0] burst_adapter_source0_channel;                                                                                  // burst_adapter:source0_channel -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                 // rst_controller:reset_out -> [addr_router_012:reset, addr_router_013:reset, cmd_xbar_demux_012:reset, cmd_xbar_demux_013:reset, crosser:out_reset, crosser_001:in_reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:out_reset, crosser_005:out_reset, crosser_006:out_reset, crosser_007:in_reset, ddr2_sdram:soft_reset_n, id_router_005:reset, id_router_020:reset, irq_synchronizer_008:receiver_reset, pll:reset_n, pll_s1_translator:reset, pll_s1_translator_avalon_universal_slave_0_agent:reset, pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_020:reset, sls_sdhc:reset_n, sls_sdhc_control_translator:reset, sls_sdhc_control_translator_avalon_universal_slave_0_agent:reset, sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sls_sdhc_read_master_translator:reset, sls_sdhc_read_master_translator_avalon_universal_master_0_agent:reset, sls_sdhc_write_master_translator:reset, sls_sdhc_write_master_translator_avalon_universal_master_0_agent:reset]
	wire          pll_resetrequest_reset;                                                                                         // pll:resetrequest -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in2, rst_controller_003:reset_in2, rst_controller_004:reset_in2, rst_controller_005:reset_in2]
	wire          cpu_jtag_debug_module_reset_reset;                                                                              // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in5, rst_controller_001:reset_in5, rst_controller_002:reset_in5, rst_controller_003:reset_in5, rst_controller_004:reset_in5, rst_controller_005:reset_in5]
	wire          rst_controller_001_reset_out_reset;                                                                             // rst_controller_001:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, addr_router_005:reset, addr_router_016:reset, addr_router_017:reset, addr_router_018:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, cmd_xbar_demux_016:reset, cmd_xbar_demux_017:reset, cmd_xbar_demux_018:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_012:reset, cmd_xbar_mux_030:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_ddr_1_clock_bridge:s0_reset, cpu_ddr_1_clock_bridge_s0_translator:reset, cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:reset, cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu_ddr_clock_bridge:s0_reset, cpu_ddr_clock_bridge_s0_translator:reset, cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:reset, cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:in_reset, crosser_001:out_reset, crosser_002:out_reset, crosser_003:out_reset, crosser_004:in_reset, crosser_005:in_reset, descriptor_memory:reset, descriptor_memory_s1_translator:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ext_flash:reset_reset, ext_flash_uas_translator:reset, ext_flash_uas_translator_avalon_universal_slave_0_agent:reset, ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, flash_tristate_bridge_bridge_0:reset, flash_tristate_bridge_pinSharer_0:reset_reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_012:reset, id_router_030:reset, id_router_031:reset, id_router_032:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, irq_synchronizer_007:sender_reset, irq_synchronizer_008:sender_reset, lcd_32_to_8_bits_dfa:reset_n, lcd_64_to_32_bits_dfa:reset_n, lcd_pixel_converter:reset_n, lcd_pixel_fifo:rdreset_n, lcd_sync_generator:reset_n, lcd_ta_fifo_to_dfa:reset_n, limiter:reset, limiter_001:reset, limiter_002:reset, limiter_003:reset, limiter_004:reset, limiter_005:reset, limiter_013:reset, max2:reset_reset, max2_uas_translator:reset, max2_uas_translator_avalon_universal_slave_0_agent:reset, max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pipeline_bridge_before_tristate_bridge:reset, pipeline_bridge_before_tristate_bridge_m0_translator:reset, pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent:reset, pipeline_bridge_before_tristate_bridge_s0_translator:reset, pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:reset, pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_030:reset, rsp_xbar_demux_031:reset, rsp_xbar_demux_032:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_018:reset, sdhc_ddr_clock_bridge:s0_reset, sdhc_ddr_clock_bridge_s0_translator:reset, sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:reset, sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_rx:system_reset_n, sgdma_rx_csr_translator:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_rx_descriptor_read_translator:reset, sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_rx_descriptor_write_translator:reset, sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_rx_m_write_translator:reset, sgdma_rx_m_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx:system_reset_n, sgdma_tx_csr_translator:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_tx_descriptor_read_translator:reset, sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_tx_descriptor_write_translator:reset, sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx_m_read_translator:reset, sgdma_tx_m_read_translator_avalon_universal_master_0_agent:reset, slow_peripheral_bridge:s0_reset, slow_peripheral_bridge_s0_translator:reset, slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:reset, slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tse_ddr_clock_bridge:s0_reset, tse_ddr_clock_bridge_s0_translator:reset, tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:reset, tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tse_mac:reset, tse_mac_control_port_translator:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter_008:reset, width_adapter_009:reset, width_adapter_010:reset, width_adapter_011:reset]
	wire          rst_controller_002_reset_out_reset;                                                                             // rst_controller_002:reset_out -> ddr2_sdram_1:soft_reset_n
	wire          rst_controller_003_reset_out_reset;                                                                             // rst_controller_003:reset_out -> [addr_router_006:reset, addr_router_007:reset, addr_router_008:reset, addr_router_009:reset, addr_router_010:reset, addr_router_011:reset, cmd_xbar_demux_006:reset, cmd_xbar_demux_007:reset, cmd_xbar_demux_008:reset, cmd_xbar_demux_009:reset, cmd_xbar_demux_010:reset, cmd_xbar_demux_011:reset, cpu_ddr_clock_bridge:m0_reset, cpu_ddr_clock_bridge_m0_translator:reset, cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:reset, id_router_011:reset, irq_synchronizer_003:receiver_reset, lcd_pixel_fifo:wrreset_n, lcd_sgdma:system_reset_n, lcd_sgdma_csr_translator:reset, lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:reset, lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_sgdma_descriptor_read_translator:reset, lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent:reset, lcd_sgdma_descriptor_write_translator:reset, lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent:reset, lcd_sgdma_m_read_translator:reset, lcd_sgdma_m_read_translator_avalon_universal_master_0_agent:reset, lcd_ta_sgdma_to_fifo:reset_n, limiter_006:reset, limiter_007:reset, limiter_008:reset, limiter_009:reset, limiter_010:reset, limiter_011:reset, rsp_xbar_demux_011:reset, rsp_xbar_mux_010:reset, sdhc_ddr_clock_bridge:m0_reset, sdhc_ddr_clock_bridge_m0_translator:reset, sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:reset, tse_ddr_clock_bridge:m0_reset, tse_ddr_clock_bridge_m0_translator:reset, tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          rst_controller_004_reset_out_reset;                                                                             // rst_controller_004:reset_out -> [addr_router_015:reset, button_pio:reset_n, button_pio_s1_translator:reset, button_pio_s1_translator_avalon_universal_slave_0_agent:reset, button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux_015:reset, crosser_006:in_reset, crosser_007:out_reset, high_res_timer:reset_n, high_res_timer_s1_translator:reset, high_res_timer_s1_translator_avalon_universal_slave_0_agent:reset, high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_021:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, id_router_025:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, id_router_029:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, irq_synchronizer_006:receiver_reset, irq_synchronizer_007:receiver_reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_i2c_en:reset_n, lcd_i2c_en_s1_translator:reset, lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:reset, lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_i2c_scl:reset_n, lcd_i2c_scl_s1_translator:reset, lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:reset, lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_i2c_sdat:reset_n, lcd_i2c_sdat_s1_translator:reset, lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:reset, lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_pio:reset_n, led_pio_s1_translator:reset, led_pio_s1_translator_avalon_universal_slave_0_agent:reset, led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_012:reset, performance_counter:reset_n, performance_counter_control_slave_translator:reset, performance_counter_control_slave_translator_avalon_universal_slave_0_agent:reset, performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_id_eeprom_dat:reset_n, pio_id_eeprom_dat_s1_translator:reset, pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:reset, pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_id_eeprom_scl:reset_n, pio_id_eeprom_scl_s1_translator:reset, pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:reset, pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_demux_029:reset, rsp_xbar_mux_015:reset, slow_peripheral_bridge:m0_reset, slow_peripheral_bridge_m0_translator:reset, slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:reset, sys_clk_timer:reset_n, sys_clk_timer_s1_translator:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, touch_panel_pen_irq_n:reset_n, touch_panel_pen_irq_n_s1_translator:reset, touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:reset, touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, touch_panel_spi:reset_n, touch_panel_spi_spi_control_port_translator:reset, touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:reset, touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart1:reset_n, uart1_s1_translator:reset, uart1_s1_translator_avalon_universal_slave_0_agent:reset, uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_005_reset_out_reset;                                                                             // rst_controller_005:reset_out -> [addr_router_014:reset, cmd_xbar_demux_014:reset, cpu_ddr_1_clock_bridge:m0_reset, cpu_ddr_1_clock_bridge_m0_translator:reset, cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                      // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                              // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire   [88:0] cmd_xbar_demux_src0_data;                                                                                       // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire    [9:0] cmd_xbar_demux_src0_channel;                                                                                    // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                      // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                      // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                              // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire   [88:0] cmd_xbar_demux_src1_data;                                                                                       // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire    [9:0] cmd_xbar_demux_src1_channel;                                                                                    // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                      // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                                // cmd_xbar_demux:src2_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                      // cmd_xbar_demux:src2_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                              // cmd_xbar_demux:src2_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_demux_src2_data;                                                                                       // cmd_xbar_demux:src2_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [9:0] cmd_xbar_demux_src2_channel;                                                                                    // cmd_xbar_demux:src2_channel -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src3_endofpacket;                                                                                // cmd_xbar_demux:src3_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                                      // cmd_xbar_demux:src3_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                              // cmd_xbar_demux:src3_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_demux_src3_data;                                                                                       // cmd_xbar_demux:src3_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [9:0] cmd_xbar_demux_src3_channel;                                                                                    // cmd_xbar_demux:src3_channel -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src4_endofpacket;                                                                                // cmd_xbar_demux:src4_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                                      // cmd_xbar_demux:src4_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                                              // cmd_xbar_demux:src4_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_demux_src4_data;                                                                                       // cmd_xbar_demux:src4_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire    [9:0] cmd_xbar_demux_src4_channel;                                                                                    // cmd_xbar_demux:src4_channel -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src6_endofpacket;                                                                                // cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire          cmd_xbar_demux_src6_valid;                                                                                      // cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire          cmd_xbar_demux_src6_startofpacket;                                                                              // cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire   [88:0] cmd_xbar_demux_src6_data;                                                                                       // cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	wire    [9:0] cmd_xbar_demux_src6_channel;                                                                                    // cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire          cmd_xbar_demux_src6_ready;                                                                                      // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	wire          cmd_xbar_demux_src7_endofpacket;                                                                                // cmd_xbar_demux:src7_endofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src7_valid;                                                                                      // cmd_xbar_demux:src7_valid -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src7_startofpacket;                                                                              // cmd_xbar_demux:src7_startofpacket -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_demux_src7_data;                                                                                       // cmd_xbar_demux:src7_data -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [9:0] cmd_xbar_demux_src7_channel;                                                                                    // cmd_xbar_demux:src7_channel -> cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src8_endofpacket;                                                                                // cmd_xbar_demux:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire          cmd_xbar_demux_src8_valid;                                                                                      // cmd_xbar_demux:src8_valid -> cmd_xbar_mux_008:sink0_valid
	wire          cmd_xbar_demux_src8_startofpacket;                                                                              // cmd_xbar_demux:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire   [88:0] cmd_xbar_demux_src8_data;                                                                                       // cmd_xbar_demux:src8_data -> cmd_xbar_mux_008:sink0_data
	wire    [9:0] cmd_xbar_demux_src8_channel;                                                                                    // cmd_xbar_demux:src8_channel -> cmd_xbar_mux_008:sink0_channel
	wire          cmd_xbar_demux_src8_ready;                                                                                      // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux:src8_ready
	wire          cmd_xbar_demux_src9_endofpacket;                                                                                // cmd_xbar_demux:src9_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src9_valid;                                                                                      // cmd_xbar_demux:src9_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src9_startofpacket;                                                                              // cmd_xbar_demux:src9_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_demux_src9_data;                                                                                       // cmd_xbar_demux:src9_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [9:0] cmd_xbar_demux_src9_channel;                                                                                    // cmd_xbar_demux:src9_channel -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                            // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                  // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                          // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire   [88:0] cmd_xbar_demux_001_src0_data;                                                                                   // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire    [9:0] cmd_xbar_demux_001_src0_channel;                                                                                // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                  // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                            // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                  // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_006:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                          // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire   [88:0] cmd_xbar_demux_001_src1_data;                                                                                   // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_006:sink1_data
	wire    [9:0] cmd_xbar_demux_001_src1_channel;                                                                                // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_006:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                  // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                            // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                  // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_008:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                          // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire   [88:0] cmd_xbar_demux_001_src2_data;                                                                                   // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_008:sink1_data
	wire    [9:0] cmd_xbar_demux_001_src2_channel;                                                                                // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_008:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                                  // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                            // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                                  // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                          // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire   [88:0] cmd_xbar_demux_002_src0_data;                                                                                   // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_001:sink1_data
	wire    [9:0] cmd_xbar_demux_002_src0_channel;                                                                                // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                                  // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                            // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                                  // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_001:sink2_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                          // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire   [88:0] cmd_xbar_demux_003_src0_data;                                                                                   // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_001:sink2_data
	wire    [9:0] cmd_xbar_demux_003_src0_channel;                                                                                // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_001:sink2_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                                  // cmd_xbar_mux_001:sink2_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                            // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_001:sink3_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                                  // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_001:sink3_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                                          // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_001:sink3_startofpacket
	wire   [88:0] cmd_xbar_demux_004_src0_data;                                                                                   // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_001:sink3_data
	wire    [9:0] cmd_xbar_demux_004_src0_channel;                                                                                // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_001:sink3_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                                  // cmd_xbar_mux_001:sink3_ready -> cmd_xbar_demux_004:src0_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                            // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_001:sink4_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                                  // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_001:sink4_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                                          // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_001:sink4_startofpacket
	wire   [88:0] cmd_xbar_demux_005_src0_data;                                                                                   // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_001:sink4_data
	wire    [9:0] cmd_xbar_demux_005_src0_channel;                                                                                // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_001:sink4_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                                  // cmd_xbar_mux_001:sink4_ready -> cmd_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                      // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                              // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire   [88:0] rsp_xbar_demux_src0_data;                                                                                       // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [9:0] rsp_xbar_demux_src0_channel;                                                                                    // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                      // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                      // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                              // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire   [88:0] rsp_xbar_demux_src1_data;                                                                                       // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [9:0] rsp_xbar_demux_src1_channel;                                                                                    // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                      // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                            // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                  // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                          // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src0_data;                                                                                   // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [9:0] rsp_xbar_demux_001_src0_channel;                                                                                // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                  // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                            // rsp_xbar_demux_001:src1_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                  // rsp_xbar_demux_001:src1_valid -> limiter_002:rsp_sink_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                          // rsp_xbar_demux_001:src1_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src1_data;                                                                                   // rsp_xbar_demux_001:src1_data -> limiter_002:rsp_sink_data
	wire    [9:0] rsp_xbar_demux_001_src1_channel;                                                                                // rsp_xbar_demux_001:src1_channel -> limiter_002:rsp_sink_channel
	wire          rsp_xbar_demux_001_src2_endofpacket;                                                                            // rsp_xbar_demux_001:src2_endofpacket -> limiter_003:rsp_sink_endofpacket
	wire          rsp_xbar_demux_001_src2_valid;                                                                                  // rsp_xbar_demux_001:src2_valid -> limiter_003:rsp_sink_valid
	wire          rsp_xbar_demux_001_src2_startofpacket;                                                                          // rsp_xbar_demux_001:src2_startofpacket -> limiter_003:rsp_sink_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src2_data;                                                                                   // rsp_xbar_demux_001:src2_data -> limiter_003:rsp_sink_data
	wire    [9:0] rsp_xbar_demux_001_src2_channel;                                                                                // rsp_xbar_demux_001:src2_channel -> limiter_003:rsp_sink_channel
	wire          rsp_xbar_demux_001_src3_endofpacket;                                                                            // rsp_xbar_demux_001:src3_endofpacket -> limiter_004:rsp_sink_endofpacket
	wire          rsp_xbar_demux_001_src3_valid;                                                                                  // rsp_xbar_demux_001:src3_valid -> limiter_004:rsp_sink_valid
	wire          rsp_xbar_demux_001_src3_startofpacket;                                                                          // rsp_xbar_demux_001:src3_startofpacket -> limiter_004:rsp_sink_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src3_data;                                                                                   // rsp_xbar_demux_001:src3_data -> limiter_004:rsp_sink_data
	wire    [9:0] rsp_xbar_demux_001_src3_channel;                                                                                // rsp_xbar_demux_001:src3_channel -> limiter_004:rsp_sink_channel
	wire          rsp_xbar_demux_001_src4_endofpacket;                                                                            // rsp_xbar_demux_001:src4_endofpacket -> limiter_005:rsp_sink_endofpacket
	wire          rsp_xbar_demux_001_src4_valid;                                                                                  // rsp_xbar_demux_001:src4_valid -> limiter_005:rsp_sink_valid
	wire          rsp_xbar_demux_001_src4_startofpacket;                                                                          // rsp_xbar_demux_001:src4_startofpacket -> limiter_005:rsp_sink_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src4_data;                                                                                   // rsp_xbar_demux_001:src4_data -> limiter_005:rsp_sink_data
	wire    [9:0] rsp_xbar_demux_001_src4_channel;                                                                                // rsp_xbar_demux_001:src4_channel -> limiter_005:rsp_sink_channel
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                            // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                  // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                          // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire   [88:0] rsp_xbar_demux_002_src0_data;                                                                                   // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [9:0] rsp_xbar_demux_002_src0_channel;                                                                                // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                  // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                            // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                  // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                          // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire   [88:0] rsp_xbar_demux_003_src0_data;                                                                                   // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire    [9:0] rsp_xbar_demux_003_src0_channel;                                                                                // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                  // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                            // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                  // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                          // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire   [88:0] rsp_xbar_demux_004_src0_data;                                                                                   // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire    [9:0] rsp_xbar_demux_004_src0_channel;                                                                                // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                  // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                            // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                  // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                          // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire   [88:0] rsp_xbar_demux_006_src0_data;                                                                                   // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire    [9:0] rsp_xbar_demux_006_src0_channel;                                                                                // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                  // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_006_src1_endofpacket;                                                                            // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_006_src1_valid;                                                                                  // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_006_src1_startofpacket;                                                                          // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire   [88:0] rsp_xbar_demux_006_src1_data;                                                                                   // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink1_data
	wire    [9:0] rsp_xbar_demux_006_src1_channel;                                                                                // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_006_src1_ready;                                                                                  // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_006:src1_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                            // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                  // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                          // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire   [88:0] rsp_xbar_demux_007_src0_data;                                                                                   // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire    [9:0] rsp_xbar_demux_007_src0_channel;                                                                                // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                  // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                            // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                  // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                          // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire   [88:0] rsp_xbar_demux_008_src0_data;                                                                                   // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	wire    [9:0] rsp_xbar_demux_008_src0_channel;                                                                                // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                  // rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_008_src1_endofpacket;                                                                            // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_008_src1_valid;                                                                                  // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_008_src1_startofpacket;                                                                          // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire   [88:0] rsp_xbar_demux_008_src1_data;                                                                                   // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_001:sink2_data
	wire    [9:0] rsp_xbar_demux_008_src1_channel;                                                                                // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_008_src1_ready;                                                                                  // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_008:src1_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                            // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                  // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                          // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	wire   [88:0] rsp_xbar_demux_009_src0_data;                                                                                   // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	wire    [9:0] rsp_xbar_demux_009_src0_channel;                                                                                // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                  // rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                                    // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                                  // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire   [88:0] limiter_cmd_src_data;                                                                                           // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [9:0] limiter_cmd_src_channel;                                                                                        // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                          // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                   // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                         // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                 // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire   [88:0] rsp_xbar_mux_src_data;                                                                                          // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [9:0] rsp_xbar_mux_src_channel;                                                                                       // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                         // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                                // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                              // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire   [88:0] limiter_001_cmd_src_data;                                                                                       // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire    [9:0] limiter_001_cmd_src_channel;                                                                                    // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                                      // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                               // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                     // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                             // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire   [88:0] rsp_xbar_mux_001_src_data;                                                                                      // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire    [9:0] rsp_xbar_mux_001_src_channel;                                                                                   // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                     // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          limiter_002_cmd_src_endofpacket;                                                                                // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          limiter_002_cmd_src_startofpacket;                                                                              // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [88:0] limiter_002_cmd_src_data;                                                                                       // limiter_002:cmd_src_data -> cmd_xbar_demux_002:sink_data
	wire    [9:0] limiter_002_cmd_src_channel;                                                                                    // limiter_002:cmd_src_channel -> cmd_xbar_demux_002:sink_channel
	wire          limiter_002_cmd_src_ready;                                                                                      // cmd_xbar_demux_002:sink_ready -> limiter_002:cmd_src_ready
	wire          rsp_xbar_demux_001_src1_ready;                                                                                  // limiter_002:rsp_sink_ready -> rsp_xbar_demux_001:src1_ready
	wire          limiter_003_cmd_src_endofpacket;                                                                                // limiter_003:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          limiter_003_cmd_src_startofpacket;                                                                              // limiter_003:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire   [88:0] limiter_003_cmd_src_data;                                                                                       // limiter_003:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire    [9:0] limiter_003_cmd_src_channel;                                                                                    // limiter_003:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire          limiter_003_cmd_src_ready;                                                                                      // cmd_xbar_demux_003:sink_ready -> limiter_003:cmd_src_ready
	wire          rsp_xbar_demux_001_src2_ready;                                                                                  // limiter_003:rsp_sink_ready -> rsp_xbar_demux_001:src2_ready
	wire          limiter_004_cmd_src_endofpacket;                                                                                // limiter_004:cmd_src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          limiter_004_cmd_src_startofpacket;                                                                              // limiter_004:cmd_src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire   [88:0] limiter_004_cmd_src_data;                                                                                       // limiter_004:cmd_src_data -> cmd_xbar_demux_004:sink_data
	wire    [9:0] limiter_004_cmd_src_channel;                                                                                    // limiter_004:cmd_src_channel -> cmd_xbar_demux_004:sink_channel
	wire          limiter_004_cmd_src_ready;                                                                                      // cmd_xbar_demux_004:sink_ready -> limiter_004:cmd_src_ready
	wire          rsp_xbar_demux_001_src3_ready;                                                                                  // limiter_004:rsp_sink_ready -> rsp_xbar_demux_001:src3_ready
	wire          limiter_005_cmd_src_endofpacket;                                                                                // limiter_005:cmd_src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          limiter_005_cmd_src_startofpacket;                                                                              // limiter_005:cmd_src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire   [88:0] limiter_005_cmd_src_data;                                                                                       // limiter_005:cmd_src_data -> cmd_xbar_demux_005:sink_data
	wire    [9:0] limiter_005_cmd_src_channel;                                                                                    // limiter_005:cmd_src_channel -> cmd_xbar_demux_005:sink_channel
	wire          limiter_005_cmd_src_ready;                                                                                      // cmd_xbar_demux_005:sink_ready -> limiter_005:cmd_src_ready
	wire          rsp_xbar_demux_001_src4_ready;                                                                                  // limiter_005:rsp_sink_ready -> rsp_xbar_demux_001:src4_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                   // cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                         // cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                 // cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_mux_src_data;                                                                                          // cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire    [9:0] cmd_xbar_mux_src_channel;                                                                                       // cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                      // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                            // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                    // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire   [88:0] id_router_src_data;                                                                                             // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [9:0] id_router_src_channel;                                                                                          // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                            // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                               // cmd_xbar_mux_001:src_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                     // cmd_xbar_mux_001:src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                             // cmd_xbar_mux_001:src_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_mux_001_src_data;                                                                                      // cmd_xbar_mux_001:src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [9:0] cmd_xbar_mux_001_src_channel;                                                                                   // cmd_xbar_mux_001:src_channel -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                     // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                                  // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                        // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [88:0] id_router_001_src_data;                                                                                         // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [9:0] id_router_001_src_channel;                                                                                      // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                        // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_src2_ready;                                                                                      // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire          id_router_002_src_endofpacket;                                                                                  // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                        // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                                // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [88:0] id_router_002_src_data;                                                                                         // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [9:0] id_router_002_src_channel;                                                                                      // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                        // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_src3_ready;                                                                                      // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src3_ready
	wire          id_router_003_src_endofpacket;                                                                                  // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                        // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire   [88:0] id_router_003_src_data;                                                                                         // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [9:0] id_router_003_src_channel;                                                                                      // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                        // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_src4_ready;                                                                                      // tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src4_ready
	wire          id_router_004_src_endofpacket;                                                                                  // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                        // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire   [88:0] id_router_004_src_data;                                                                                         // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [9:0] id_router_004_src_channel;                                                                                      // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                        // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          crosser_out_ready;                                                                                              // sls_sdhc_control_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_005_src_endofpacket;                                                                                  // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                        // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                                // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire   [88:0] id_router_005_src_data;                                                                                         // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire    [9:0] id_router_005_src_channel;                                                                                      // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                        // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_mux_006_src_endofpacket;                                                                               // cmd_xbar_mux_006:src_endofpacket -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_006_src_valid;                                                                                     // cmd_xbar_mux_006:src_valid -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_006_src_startofpacket;                                                                             // cmd_xbar_mux_006:src_startofpacket -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_mux_006_src_data;                                                                                      // cmd_xbar_mux_006:src_data -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [9:0] cmd_xbar_mux_006_src_channel;                                                                                   // cmd_xbar_mux_006:src_channel -> pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_006_src_ready;                                                                                     // pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	wire          id_router_006_src_endofpacket;                                                                                  // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                        // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [88:0] id_router_006_src_data;                                                                                         // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire    [9:0] id_router_006_src_channel;                                                                                      // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                        // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_src7_ready;                                                                                      // cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src7_ready
	wire          id_router_007_src_endofpacket;                                                                                  // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                        // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [88:0] id_router_007_src_data;                                                                                         // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire    [9:0] id_router_007_src_channel;                                                                                      // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                        // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_mux_008_src_endofpacket;                                                                               // cmd_xbar_mux_008:src_endofpacket -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_008_src_valid;                                                                                     // cmd_xbar_mux_008:src_valid -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_008_src_startofpacket;                                                                             // cmd_xbar_mux_008:src_startofpacket -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_mux_008_src_data;                                                                                      // cmd_xbar_mux_008:src_data -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [9:0] cmd_xbar_mux_008_src_channel;                                                                                   // cmd_xbar_mux_008:src_channel -> cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_008_src_ready;                                                                                     // cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire          id_router_008_src_endofpacket;                                                                                  // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                        // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [88:0] id_router_008_src_data;                                                                                         // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire    [9:0] id_router_008_src_channel;                                                                                      // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                        // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_src9_ready;                                                                                      // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src9_ready
	wire          id_router_009_src_endofpacket;                                                                                  // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                        // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire   [88:0] id_router_009_src_data;                                                                                         // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire    [9:0] id_router_009_src_channel;                                                                                      // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                        // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_008_src0_endofpacket;                                                                            // cmd_xbar_demux_008:src0_endofpacket -> cmd_xbar_mux_010:sink2_endofpacket
	wire          cmd_xbar_demux_008_src0_valid;                                                                                  // cmd_xbar_demux_008:src0_valid -> cmd_xbar_mux_010:sink2_valid
	wire          cmd_xbar_demux_008_src0_startofpacket;                                                                          // cmd_xbar_demux_008:src0_startofpacket -> cmd_xbar_mux_010:sink2_startofpacket
	wire  [124:0] cmd_xbar_demux_008_src0_data;                                                                                   // cmd_xbar_demux_008:src0_data -> cmd_xbar_mux_010:sink2_data
	wire    [5:0] cmd_xbar_demux_008_src0_channel;                                                                                // cmd_xbar_demux_008:src0_channel -> cmd_xbar_mux_010:sink2_channel
	wire          cmd_xbar_demux_008_src0_ready;                                                                                  // cmd_xbar_mux_010:sink2_ready -> cmd_xbar_demux_008:src0_ready
	wire          cmd_xbar_demux_009_src0_endofpacket;                                                                            // cmd_xbar_demux_009:src0_endofpacket -> cmd_xbar_mux_010:sink3_endofpacket
	wire          cmd_xbar_demux_009_src0_valid;                                                                                  // cmd_xbar_demux_009:src0_valid -> cmd_xbar_mux_010:sink3_valid
	wire          cmd_xbar_demux_009_src0_startofpacket;                                                                          // cmd_xbar_demux_009:src0_startofpacket -> cmd_xbar_mux_010:sink3_startofpacket
	wire  [124:0] cmd_xbar_demux_009_src0_data;                                                                                   // cmd_xbar_demux_009:src0_data -> cmd_xbar_mux_010:sink3_data
	wire    [5:0] cmd_xbar_demux_009_src0_channel;                                                                                // cmd_xbar_demux_009:src0_channel -> cmd_xbar_mux_010:sink3_channel
	wire          cmd_xbar_demux_009_src0_ready;                                                                                  // cmd_xbar_mux_010:sink3_ready -> cmd_xbar_demux_009:src0_ready
	wire          cmd_xbar_demux_010_src1_endofpacket;                                                                            // cmd_xbar_demux_010:src1_endofpacket -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_010_src1_valid;                                                                                  // cmd_xbar_demux_010:src1_valid -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_010_src1_startofpacket;                                                                          // cmd_xbar_demux_010:src1_startofpacket -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_demux_010_src1_data;                                                                                   // cmd_xbar_demux_010:src1_data -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_demux_010_src1_channel;                                                                                // cmd_xbar_demux_010:src1_channel -> lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_010_src2_endofpacket;                                                                            // rsp_xbar_demux_010:src2_endofpacket -> limiter_008:rsp_sink_endofpacket
	wire          rsp_xbar_demux_010_src2_valid;                                                                                  // rsp_xbar_demux_010:src2_valid -> limiter_008:rsp_sink_valid
	wire          rsp_xbar_demux_010_src2_startofpacket;                                                                          // rsp_xbar_demux_010:src2_startofpacket -> limiter_008:rsp_sink_startofpacket
	wire  [124:0] rsp_xbar_demux_010_src2_data;                                                                                   // rsp_xbar_demux_010:src2_data -> limiter_008:rsp_sink_data
	wire    [5:0] rsp_xbar_demux_010_src2_channel;                                                                                // rsp_xbar_demux_010:src2_channel -> limiter_008:rsp_sink_channel
	wire          rsp_xbar_demux_010_src3_endofpacket;                                                                            // rsp_xbar_demux_010:src3_endofpacket -> limiter_009:rsp_sink_endofpacket
	wire          rsp_xbar_demux_010_src3_valid;                                                                                  // rsp_xbar_demux_010:src3_valid -> limiter_009:rsp_sink_valid
	wire          rsp_xbar_demux_010_src3_startofpacket;                                                                          // rsp_xbar_demux_010:src3_startofpacket -> limiter_009:rsp_sink_startofpacket
	wire  [124:0] rsp_xbar_demux_010_src3_data;                                                                                   // rsp_xbar_demux_010:src3_data -> limiter_009:rsp_sink_data
	wire    [5:0] rsp_xbar_demux_010_src3_channel;                                                                                // rsp_xbar_demux_010:src3_channel -> limiter_009:rsp_sink_channel
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                            // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_010:sink1_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                  // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_010:sink1_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                          // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_010:sink1_startofpacket
	wire   [88:0] rsp_xbar_demux_011_src0_data;                                                                                   // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_010:sink1_data
	wire    [5:0] rsp_xbar_demux_011_src0_channel;                                                                                // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_010:sink1_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                  // rsp_xbar_mux_010:sink1_ready -> rsp_xbar_demux_011:src0_ready
	wire          limiter_006_cmd_src_endofpacket;                                                                                // limiter_006:cmd_src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	wire          limiter_006_cmd_src_startofpacket;                                                                              // limiter_006:cmd_src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	wire   [88:0] limiter_006_cmd_src_data;                                                                                       // limiter_006:cmd_src_data -> cmd_xbar_demux_006:sink_data
	wire    [5:0] limiter_006_cmd_src_channel;                                                                                    // limiter_006:cmd_src_channel -> cmd_xbar_demux_006:sink_channel
	wire          limiter_006_cmd_src_ready;                                                                                      // cmd_xbar_demux_006:sink_ready -> limiter_006:cmd_src_ready
	wire          width_adapter_004_src_ready;                                                                                    // limiter_006:rsp_sink_ready -> width_adapter_004:out_ready
	wire          limiter_007_cmd_src_endofpacket;                                                                                // limiter_007:cmd_src_endofpacket -> cmd_xbar_demux_007:sink_endofpacket
	wire          limiter_007_cmd_src_startofpacket;                                                                              // limiter_007:cmd_src_startofpacket -> cmd_xbar_demux_007:sink_startofpacket
	wire   [88:0] limiter_007_cmd_src_data;                                                                                       // limiter_007:cmd_src_data -> cmd_xbar_demux_007:sink_data
	wire    [5:0] limiter_007_cmd_src_channel;                                                                                    // limiter_007:cmd_src_channel -> cmd_xbar_demux_007:sink_channel
	wire          limiter_007_cmd_src_ready;                                                                                      // cmd_xbar_demux_007:sink_ready -> limiter_007:cmd_src_ready
	wire          width_adapter_005_src_ready;                                                                                    // limiter_007:rsp_sink_ready -> width_adapter_005:out_ready
	wire          limiter_008_cmd_src_endofpacket;                                                                                // limiter_008:cmd_src_endofpacket -> cmd_xbar_demux_008:sink_endofpacket
	wire          limiter_008_cmd_src_startofpacket;                                                                              // limiter_008:cmd_src_startofpacket -> cmd_xbar_demux_008:sink_startofpacket
	wire  [124:0] limiter_008_cmd_src_data;                                                                                       // limiter_008:cmd_src_data -> cmd_xbar_demux_008:sink_data
	wire    [5:0] limiter_008_cmd_src_channel;                                                                                    // limiter_008:cmd_src_channel -> cmd_xbar_demux_008:sink_channel
	wire          limiter_008_cmd_src_ready;                                                                                      // cmd_xbar_demux_008:sink_ready -> limiter_008:cmd_src_ready
	wire          rsp_xbar_demux_010_src2_ready;                                                                                  // limiter_008:rsp_sink_ready -> rsp_xbar_demux_010:src2_ready
	wire          limiter_009_cmd_src_endofpacket;                                                                                // limiter_009:cmd_src_endofpacket -> cmd_xbar_demux_009:sink_endofpacket
	wire          limiter_009_cmd_src_startofpacket;                                                                              // limiter_009:cmd_src_startofpacket -> cmd_xbar_demux_009:sink_startofpacket
	wire  [124:0] limiter_009_cmd_src_data;                                                                                       // limiter_009:cmd_src_data -> cmd_xbar_demux_009:sink_data
	wire    [5:0] limiter_009_cmd_src_channel;                                                                                    // limiter_009:cmd_src_channel -> cmd_xbar_demux_009:sink_channel
	wire          limiter_009_cmd_src_ready;                                                                                      // cmd_xbar_demux_009:sink_ready -> limiter_009:cmd_src_ready
	wire          rsp_xbar_demux_010_src3_ready;                                                                                  // limiter_009:rsp_sink_ready -> rsp_xbar_demux_010:src3_ready
	wire          limiter_010_cmd_src_endofpacket;                                                                                // limiter_010:cmd_src_endofpacket -> cmd_xbar_demux_010:sink_endofpacket
	wire          limiter_010_cmd_src_startofpacket;                                                                              // limiter_010:cmd_src_startofpacket -> cmd_xbar_demux_010:sink_startofpacket
	wire   [88:0] limiter_010_cmd_src_data;                                                                                       // limiter_010:cmd_src_data -> cmd_xbar_demux_010:sink_data
	wire    [5:0] limiter_010_cmd_src_channel;                                                                                    // limiter_010:cmd_src_channel -> cmd_xbar_demux_010:sink_channel
	wire          limiter_010_cmd_src_ready;                                                                                      // cmd_xbar_demux_010:sink_ready -> limiter_010:cmd_src_ready
	wire          rsp_xbar_mux_010_src_endofpacket;                                                                               // rsp_xbar_mux_010:src_endofpacket -> limiter_010:rsp_sink_endofpacket
	wire          rsp_xbar_mux_010_src_valid;                                                                                     // rsp_xbar_mux_010:src_valid -> limiter_010:rsp_sink_valid
	wire          rsp_xbar_mux_010_src_startofpacket;                                                                             // rsp_xbar_mux_010:src_startofpacket -> limiter_010:rsp_sink_startofpacket
	wire   [88:0] rsp_xbar_mux_010_src_data;                                                                                      // rsp_xbar_mux_010:src_data -> limiter_010:rsp_sink_data
	wire    [5:0] rsp_xbar_mux_010_src_channel;                                                                                   // rsp_xbar_mux_010:src_channel -> limiter_010:rsp_sink_channel
	wire          rsp_xbar_mux_010_src_ready;                                                                                     // limiter_010:rsp_sink_ready -> rsp_xbar_mux_010:src_ready
	wire          limiter_011_cmd_src_endofpacket;                                                                                // limiter_011:cmd_src_endofpacket -> cmd_xbar_demux_011:sink_endofpacket
	wire          limiter_011_cmd_src_startofpacket;                                                                              // limiter_011:cmd_src_startofpacket -> cmd_xbar_demux_011:sink_startofpacket
	wire   [88:0] limiter_011_cmd_src_data;                                                                                       // limiter_011:cmd_src_data -> cmd_xbar_demux_011:sink_data
	wire    [5:0] limiter_011_cmd_src_channel;                                                                                    // limiter_011:cmd_src_channel -> cmd_xbar_demux_011:sink_channel
	wire          limiter_011_cmd_src_ready;                                                                                      // cmd_xbar_demux_011:sink_ready -> limiter_011:cmd_src_ready
	wire          width_adapter_007_src_ready;                                                                                    // limiter_011:rsp_sink_ready -> width_adapter_007:out_ready
	wire          cmd_xbar_mux_010_src_endofpacket;                                                                               // cmd_xbar_mux_010:src_endofpacket -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_010_src_valid;                                                                                     // cmd_xbar_mux_010:src_valid -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_010_src_startofpacket;                                                                             // cmd_xbar_mux_010:src_startofpacket -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [124:0] cmd_xbar_mux_010_src_data;                                                                                      // cmd_xbar_mux_010:src_data -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_010_src_channel;                                                                                   // cmd_xbar_mux_010:src_channel -> ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_010_src_ready;                                                                                     // ddr2_sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	wire          id_router_010_src_endofpacket;                                                                                  // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                        // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                                // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [124:0] id_router_010_src_data;                                                                                         // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire    [5:0] id_router_010_src_channel;                                                                                      // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                        // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_010_src1_ready;                                                                                  // lcd_sgdma_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_010:src1_ready
	wire          id_router_011_src_endofpacket;                                                                                  // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                        // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                                // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire   [88:0] id_router_011_src_data;                                                                                         // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire    [5:0] id_router_011_src_channel;                                                                                      // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                        // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          addr_router_012_src_endofpacket;                                                                                // addr_router_012:src_endofpacket -> cmd_xbar_demux_012:sink_endofpacket
	wire          addr_router_012_src_valid;                                                                                      // addr_router_012:src_valid -> cmd_xbar_demux_012:sink_valid
	wire          addr_router_012_src_startofpacket;                                                                              // addr_router_012:src_startofpacket -> cmd_xbar_demux_012:sink_startofpacket
	wire   [86:0] addr_router_012_src_data;                                                                                       // addr_router_012:src_data -> cmd_xbar_demux_012:sink_data
	wire    [1:0] addr_router_012_src_channel;                                                                                    // addr_router_012:src_channel -> cmd_xbar_demux_012:sink_channel
	wire          addr_router_012_src_ready;                                                                                      // cmd_xbar_demux_012:sink_ready -> addr_router_012:src_ready
	wire          crosser_004_out_ready;                                                                                          // sls_sdhc_read_master_translator_avalon_universal_master_0_agent:rp_ready -> crosser_004:out_ready
	wire          addr_router_013_src_endofpacket;                                                                                // addr_router_013:src_endofpacket -> cmd_xbar_demux_013:sink_endofpacket
	wire          addr_router_013_src_valid;                                                                                      // addr_router_013:src_valid -> cmd_xbar_demux_013:sink_valid
	wire          addr_router_013_src_startofpacket;                                                                              // addr_router_013:src_startofpacket -> cmd_xbar_demux_013:sink_startofpacket
	wire   [86:0] addr_router_013_src_data;                                                                                       // addr_router_013:src_data -> cmd_xbar_demux_013:sink_data
	wire    [1:0] addr_router_013_src_channel;                                                                                    // addr_router_013:src_channel -> cmd_xbar_demux_013:sink_channel
	wire          addr_router_013_src_ready;                                                                                      // cmd_xbar_demux_013:sink_ready -> addr_router_013:src_ready
	wire          crosser_005_out_ready;                                                                                          // sls_sdhc_write_master_translator_avalon_universal_master_0_agent:rp_ready -> crosser_005:out_ready
	wire          cmd_xbar_demux_014_src0_endofpacket;                                                                            // cmd_xbar_demux_014:src0_endofpacket -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_014_src0_valid;                                                                                  // cmd_xbar_demux_014:src0_valid -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_014_src0_startofpacket;                                                                          // cmd_xbar_demux_014:src0_startofpacket -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [78:0] cmd_xbar_demux_014_src0_data;                                                                                   // cmd_xbar_demux_014:src0_data -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [0:0] cmd_xbar_demux_014_src0_channel;                                                                                // cmd_xbar_demux_014:src0_channel -> ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                            // rsp_xbar_demux_013:src0_endofpacket -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                  // rsp_xbar_demux_013:src0_valid -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                          // rsp_xbar_demux_013:src0_startofpacket -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [78:0] rsp_xbar_demux_013_src0_data;                                                                                   // rsp_xbar_demux_013:src0_data -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [0:0] rsp_xbar_demux_013_src0_channel;                                                                                // rsp_xbar_demux_013:src0_channel -> cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_014_src_endofpacket;                                                                                // addr_router_014:src_endofpacket -> cmd_xbar_demux_014:sink_endofpacket
	wire          addr_router_014_src_valid;                                                                                      // addr_router_014:src_valid -> cmd_xbar_demux_014:sink_valid
	wire          addr_router_014_src_startofpacket;                                                                              // addr_router_014:src_startofpacket -> cmd_xbar_demux_014:sink_startofpacket
	wire   [78:0] addr_router_014_src_data;                                                                                       // addr_router_014:src_data -> cmd_xbar_demux_014:sink_data
	wire    [0:0] addr_router_014_src_channel;                                                                                    // addr_router_014:src_channel -> cmd_xbar_demux_014:sink_channel
	wire          addr_router_014_src_ready;                                                                                      // cmd_xbar_demux_014:sink_ready -> addr_router_014:src_ready
	wire          rsp_xbar_demux_013_src0_ready;                                                                                  // cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_013:src0_ready
	wire          cmd_xbar_demux_014_src0_ready;                                                                                  // ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_014:src0_ready
	wire          id_router_013_src_endofpacket;                                                                                  // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                        // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                                // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire   [78:0] id_router_013_src_data;                                                                                         // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire    [0:0] id_router_013_src_channel;                                                                                      // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                        // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_015_src0_endofpacket;                                                                            // cmd_xbar_demux_015:src0_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src0_valid;                                                                                  // cmd_xbar_demux_015:src0_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src0_startofpacket;                                                                          // cmd_xbar_demux_015:src0_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src0_data;                                                                                   // cmd_xbar_demux_015:src0_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src0_channel;                                                                                // cmd_xbar_demux_015:src0_channel -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src1_endofpacket;                                                                            // cmd_xbar_demux_015:src1_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src1_valid;                                                                                  // cmd_xbar_demux_015:src1_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src1_startofpacket;                                                                          // cmd_xbar_demux_015:src1_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src1_data;                                                                                   // cmd_xbar_demux_015:src1_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src1_channel;                                                                                // cmd_xbar_demux_015:src1_channel -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src2_endofpacket;                                                                            // cmd_xbar_demux_015:src2_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src2_valid;                                                                                  // cmd_xbar_demux_015:src2_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src2_startofpacket;                                                                          // cmd_xbar_demux_015:src2_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src2_data;                                                                                   // cmd_xbar_demux_015:src2_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src2_channel;                                                                                // cmd_xbar_demux_015:src2_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src3_endofpacket;                                                                            // cmd_xbar_demux_015:src3_endofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src3_valid;                                                                                  // cmd_xbar_demux_015:src3_valid -> uart1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src3_startofpacket;                                                                          // cmd_xbar_demux_015:src3_startofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src3_data;                                                                                   // cmd_xbar_demux_015:src3_data -> uart1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src3_channel;                                                                                // cmd_xbar_demux_015:src3_channel -> uart1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src4_endofpacket;                                                                            // cmd_xbar_demux_015:src4_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src4_valid;                                                                                  // cmd_xbar_demux_015:src4_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src4_startofpacket;                                                                          // cmd_xbar_demux_015:src4_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src4_data;                                                                                   // cmd_xbar_demux_015:src4_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src4_channel;                                                                                // cmd_xbar_demux_015:src4_channel -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src5_endofpacket;                                                                            // cmd_xbar_demux_015:src5_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src5_valid;                                                                                  // cmd_xbar_demux_015:src5_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src5_startofpacket;                                                                          // cmd_xbar_demux_015:src5_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src5_data;                                                                                   // cmd_xbar_demux_015:src5_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src5_channel;                                                                                // cmd_xbar_demux_015:src5_channel -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src7_endofpacket;                                                                            // cmd_xbar_demux_015:src7_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src7_valid;                                                                                  // cmd_xbar_demux_015:src7_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src7_startofpacket;                                                                          // cmd_xbar_demux_015:src7_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src7_data;                                                                                   // cmd_xbar_demux_015:src7_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src7_channel;                                                                                // cmd_xbar_demux_015:src7_channel -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src8_endofpacket;                                                                            // cmd_xbar_demux_015:src8_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src8_valid;                                                                                  // cmd_xbar_demux_015:src8_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src8_startofpacket;                                                                          // cmd_xbar_demux_015:src8_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src8_data;                                                                                   // cmd_xbar_demux_015:src8_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src8_channel;                                                                                // cmd_xbar_demux_015:src8_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src9_endofpacket;                                                                            // cmd_xbar_demux_015:src9_endofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src9_valid;                                                                                  // cmd_xbar_demux_015:src9_valid -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src9_startofpacket;                                                                          // cmd_xbar_demux_015:src9_startofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src9_data;                                                                                   // cmd_xbar_demux_015:src9_data -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src9_channel;                                                                                // cmd_xbar_demux_015:src9_channel -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src10_endofpacket;                                                                           // cmd_xbar_demux_015:src10_endofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src10_valid;                                                                                 // cmd_xbar_demux_015:src10_valid -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src10_startofpacket;                                                                         // cmd_xbar_demux_015:src10_startofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src10_data;                                                                                  // cmd_xbar_demux_015:src10_data -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src10_channel;                                                                               // cmd_xbar_demux_015:src10_channel -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src11_endofpacket;                                                                           // cmd_xbar_demux_015:src11_endofpacket -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src11_valid;                                                                                 // cmd_xbar_demux_015:src11_valid -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src11_startofpacket;                                                                         // cmd_xbar_demux_015:src11_startofpacket -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src11_data;                                                                                  // cmd_xbar_demux_015:src11_data -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src11_channel;                                                                               // cmd_xbar_demux_015:src11_channel -> lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src12_endofpacket;                                                                           // cmd_xbar_demux_015:src12_endofpacket -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src12_valid;                                                                                 // cmd_xbar_demux_015:src12_valid -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src12_startofpacket;                                                                         // cmd_xbar_demux_015:src12_startofpacket -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src12_data;                                                                                  // cmd_xbar_demux_015:src12_data -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src12_channel;                                                                               // cmd_xbar_demux_015:src12_channel -> pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src13_endofpacket;                                                                           // cmd_xbar_demux_015:src13_endofpacket -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src13_valid;                                                                                 // cmd_xbar_demux_015:src13_valid -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src13_startofpacket;                                                                         // cmd_xbar_demux_015:src13_startofpacket -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src13_data;                                                                                  // cmd_xbar_demux_015:src13_data -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src13_channel;                                                                               // cmd_xbar_demux_015:src13_channel -> pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src14_endofpacket;                                                                           // cmd_xbar_demux_015:src14_endofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src14_valid;                                                                                 // cmd_xbar_demux_015:src14_valid -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src14_startofpacket;                                                                         // cmd_xbar_demux_015:src14_startofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src14_data;                                                                                  // cmd_xbar_demux_015:src14_data -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src14_channel;                                                                               // cmd_xbar_demux_015:src14_channel -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src15_endofpacket;                                                                           // cmd_xbar_demux_015:src15_endofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_015_src15_valid;                                                                                 // cmd_xbar_demux_015:src15_valid -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_015_src15_startofpacket;                                                                         // cmd_xbar_demux_015:src15_startofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src15_data;                                                                                  // cmd_xbar_demux_015:src15_data -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_015_src15_channel;                                                                               // cmd_xbar_demux_015:src15_channel -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                            // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_015:sink0_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                                  // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_015:sink0_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                          // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_015:sink0_startofpacket
	wire   [68:0] rsp_xbar_demux_014_src0_data;                                                                                   // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_015:sink0_data
	wire   [15:0] rsp_xbar_demux_014_src0_channel;                                                                                // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_015:sink0_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                                  // rsp_xbar_mux_015:sink0_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                            // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_015:sink1_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                                  // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_015:sink1_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                          // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_015:sink1_startofpacket
	wire   [68:0] rsp_xbar_demux_015_src0_data;                                                                                   // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_015:sink1_data
	wire   [15:0] rsp_xbar_demux_015_src0_channel;                                                                                // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_015:sink1_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                                  // rsp_xbar_mux_015:sink1_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                            // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_015:sink2_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                                  // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_015:sink2_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                          // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_015:sink2_startofpacket
	wire   [68:0] rsp_xbar_demux_016_src0_data;                                                                                   // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_015:sink2_data
	wire   [15:0] rsp_xbar_demux_016_src0_channel;                                                                                // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_015:sink2_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                                  // rsp_xbar_mux_015:sink2_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                            // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_015:sink3_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                                  // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_015:sink3_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                          // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_015:sink3_startofpacket
	wire   [68:0] rsp_xbar_demux_017_src0_data;                                                                                   // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_015:sink3_data
	wire   [15:0] rsp_xbar_demux_017_src0_channel;                                                                                // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_015:sink3_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                                  // rsp_xbar_mux_015:sink3_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                            // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_015:sink4_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                                  // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_015:sink4_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                          // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_015:sink4_startofpacket
	wire   [68:0] rsp_xbar_demux_018_src0_data;                                                                                   // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_015:sink4_data
	wire   [15:0] rsp_xbar_demux_018_src0_channel;                                                                                // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_015:sink4_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                                  // rsp_xbar_mux_015:sink4_ready -> rsp_xbar_demux_018:src0_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                                            // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_015:sink5_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                                  // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_015:sink5_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                                          // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_015:sink5_startofpacket
	wire   [68:0] rsp_xbar_demux_019_src0_data;                                                                                   // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_015:sink5_data
	wire   [15:0] rsp_xbar_demux_019_src0_channel;                                                                                // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_015:sink5_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                                  // rsp_xbar_mux_015:sink5_ready -> rsp_xbar_demux_019:src0_ready
	wire          rsp_xbar_demux_021_src0_endofpacket;                                                                            // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_015:sink7_endofpacket
	wire          rsp_xbar_demux_021_src0_valid;                                                                                  // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_015:sink7_valid
	wire          rsp_xbar_demux_021_src0_startofpacket;                                                                          // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_015:sink7_startofpacket
	wire   [68:0] rsp_xbar_demux_021_src0_data;                                                                                   // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_015:sink7_data
	wire   [15:0] rsp_xbar_demux_021_src0_channel;                                                                                // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_015:sink7_channel
	wire          rsp_xbar_demux_021_src0_ready;                                                                                  // rsp_xbar_mux_015:sink7_ready -> rsp_xbar_demux_021:src0_ready
	wire          rsp_xbar_demux_022_src0_endofpacket;                                                                            // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_015:sink8_endofpacket
	wire          rsp_xbar_demux_022_src0_valid;                                                                                  // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_015:sink8_valid
	wire          rsp_xbar_demux_022_src0_startofpacket;                                                                          // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_015:sink8_startofpacket
	wire   [68:0] rsp_xbar_demux_022_src0_data;                                                                                   // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_015:sink8_data
	wire   [15:0] rsp_xbar_demux_022_src0_channel;                                                                                // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_015:sink8_channel
	wire          rsp_xbar_demux_022_src0_ready;                                                                                  // rsp_xbar_mux_015:sink8_ready -> rsp_xbar_demux_022:src0_ready
	wire          rsp_xbar_demux_023_src0_endofpacket;                                                                            // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_015:sink9_endofpacket
	wire          rsp_xbar_demux_023_src0_valid;                                                                                  // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_015:sink9_valid
	wire          rsp_xbar_demux_023_src0_startofpacket;                                                                          // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_015:sink9_startofpacket
	wire   [68:0] rsp_xbar_demux_023_src0_data;                                                                                   // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_015:sink9_data
	wire   [15:0] rsp_xbar_demux_023_src0_channel;                                                                                // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_015:sink9_channel
	wire          rsp_xbar_demux_023_src0_ready;                                                                                  // rsp_xbar_mux_015:sink9_ready -> rsp_xbar_demux_023:src0_ready
	wire          rsp_xbar_demux_024_src0_endofpacket;                                                                            // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_015:sink10_endofpacket
	wire          rsp_xbar_demux_024_src0_valid;                                                                                  // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_015:sink10_valid
	wire          rsp_xbar_demux_024_src0_startofpacket;                                                                          // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_015:sink10_startofpacket
	wire   [68:0] rsp_xbar_demux_024_src0_data;                                                                                   // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_015:sink10_data
	wire   [15:0] rsp_xbar_demux_024_src0_channel;                                                                                // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_015:sink10_channel
	wire          rsp_xbar_demux_024_src0_ready;                                                                                  // rsp_xbar_mux_015:sink10_ready -> rsp_xbar_demux_024:src0_ready
	wire          rsp_xbar_demux_025_src0_endofpacket;                                                                            // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_015:sink11_endofpacket
	wire          rsp_xbar_demux_025_src0_valid;                                                                                  // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_015:sink11_valid
	wire          rsp_xbar_demux_025_src0_startofpacket;                                                                          // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_015:sink11_startofpacket
	wire   [68:0] rsp_xbar_demux_025_src0_data;                                                                                   // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_015:sink11_data
	wire   [15:0] rsp_xbar_demux_025_src0_channel;                                                                                // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_015:sink11_channel
	wire          rsp_xbar_demux_025_src0_ready;                                                                                  // rsp_xbar_mux_015:sink11_ready -> rsp_xbar_demux_025:src0_ready
	wire          rsp_xbar_demux_026_src0_endofpacket;                                                                            // rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_015:sink12_endofpacket
	wire          rsp_xbar_demux_026_src0_valid;                                                                                  // rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_015:sink12_valid
	wire          rsp_xbar_demux_026_src0_startofpacket;                                                                          // rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_015:sink12_startofpacket
	wire   [68:0] rsp_xbar_demux_026_src0_data;                                                                                   // rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_015:sink12_data
	wire   [15:0] rsp_xbar_demux_026_src0_channel;                                                                                // rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_015:sink12_channel
	wire          rsp_xbar_demux_026_src0_ready;                                                                                  // rsp_xbar_mux_015:sink12_ready -> rsp_xbar_demux_026:src0_ready
	wire          rsp_xbar_demux_027_src0_endofpacket;                                                                            // rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux_015:sink13_endofpacket
	wire          rsp_xbar_demux_027_src0_valid;                                                                                  // rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux_015:sink13_valid
	wire          rsp_xbar_demux_027_src0_startofpacket;                                                                          // rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux_015:sink13_startofpacket
	wire   [68:0] rsp_xbar_demux_027_src0_data;                                                                                   // rsp_xbar_demux_027:src0_data -> rsp_xbar_mux_015:sink13_data
	wire   [15:0] rsp_xbar_demux_027_src0_channel;                                                                                // rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux_015:sink13_channel
	wire          rsp_xbar_demux_027_src0_ready;                                                                                  // rsp_xbar_mux_015:sink13_ready -> rsp_xbar_demux_027:src0_ready
	wire          rsp_xbar_demux_028_src0_endofpacket;                                                                            // rsp_xbar_demux_028:src0_endofpacket -> rsp_xbar_mux_015:sink14_endofpacket
	wire          rsp_xbar_demux_028_src0_valid;                                                                                  // rsp_xbar_demux_028:src0_valid -> rsp_xbar_mux_015:sink14_valid
	wire          rsp_xbar_demux_028_src0_startofpacket;                                                                          // rsp_xbar_demux_028:src0_startofpacket -> rsp_xbar_mux_015:sink14_startofpacket
	wire   [68:0] rsp_xbar_demux_028_src0_data;                                                                                   // rsp_xbar_demux_028:src0_data -> rsp_xbar_mux_015:sink14_data
	wire   [15:0] rsp_xbar_demux_028_src0_channel;                                                                                // rsp_xbar_demux_028:src0_channel -> rsp_xbar_mux_015:sink14_channel
	wire          rsp_xbar_demux_028_src0_ready;                                                                                  // rsp_xbar_mux_015:sink14_ready -> rsp_xbar_demux_028:src0_ready
	wire          rsp_xbar_demux_029_src0_endofpacket;                                                                            // rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux_015:sink15_endofpacket
	wire          rsp_xbar_demux_029_src0_valid;                                                                                  // rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux_015:sink15_valid
	wire          rsp_xbar_demux_029_src0_startofpacket;                                                                          // rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux_015:sink15_startofpacket
	wire   [68:0] rsp_xbar_demux_029_src0_data;                                                                                   // rsp_xbar_demux_029:src0_data -> rsp_xbar_mux_015:sink15_data
	wire   [15:0] rsp_xbar_demux_029_src0_channel;                                                                                // rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux_015:sink15_channel
	wire          rsp_xbar_demux_029_src0_ready;                                                                                  // rsp_xbar_mux_015:sink15_ready -> rsp_xbar_demux_029:src0_ready
	wire          limiter_012_cmd_src_endofpacket;                                                                                // limiter_012:cmd_src_endofpacket -> cmd_xbar_demux_015:sink_endofpacket
	wire          limiter_012_cmd_src_startofpacket;                                                                              // limiter_012:cmd_src_startofpacket -> cmd_xbar_demux_015:sink_startofpacket
	wire   [68:0] limiter_012_cmd_src_data;                                                                                       // limiter_012:cmd_src_data -> cmd_xbar_demux_015:sink_data
	wire   [15:0] limiter_012_cmd_src_channel;                                                                                    // limiter_012:cmd_src_channel -> cmd_xbar_demux_015:sink_channel
	wire          limiter_012_cmd_src_ready;                                                                                      // cmd_xbar_demux_015:sink_ready -> limiter_012:cmd_src_ready
	wire          rsp_xbar_mux_015_src_endofpacket;                                                                               // rsp_xbar_mux_015:src_endofpacket -> limiter_012:rsp_sink_endofpacket
	wire          rsp_xbar_mux_015_src_valid;                                                                                     // rsp_xbar_mux_015:src_valid -> limiter_012:rsp_sink_valid
	wire          rsp_xbar_mux_015_src_startofpacket;                                                                             // rsp_xbar_mux_015:src_startofpacket -> limiter_012:rsp_sink_startofpacket
	wire   [68:0] rsp_xbar_mux_015_src_data;                                                                                      // rsp_xbar_mux_015:src_data -> limiter_012:rsp_sink_data
	wire   [15:0] rsp_xbar_mux_015_src_channel;                                                                                   // rsp_xbar_mux_015:src_channel -> limiter_012:rsp_sink_channel
	wire          rsp_xbar_mux_015_src_ready;                                                                                     // limiter_012:rsp_sink_ready -> rsp_xbar_mux_015:src_ready
	wire          cmd_xbar_demux_015_src0_ready;                                                                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src0_ready
	wire          id_router_014_src_endofpacket;                                                                                  // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                        // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                                // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire   [68:0] id_router_014_src_data;                                                                                         // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [15:0] id_router_014_src_channel;                                                                                      // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                        // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_015_src1_ready;                                                                                  // high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src1_ready
	wire          id_router_015_src_endofpacket;                                                                                  // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                        // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                                // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire   [68:0] id_router_015_src_data;                                                                                         // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [15:0] id_router_015_src_channel;                                                                                      // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                        // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_015_src2_ready;                                                                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src2_ready
	wire          id_router_016_src_endofpacket;                                                                                  // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                        // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                                // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire   [68:0] id_router_016_src_data;                                                                                         // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [15:0] id_router_016_src_channel;                                                                                      // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                        // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_015_src3_ready;                                                                                  // uart1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src3_ready
	wire          id_router_017_src_endofpacket;                                                                                  // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                        // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                                // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire   [68:0] id_router_017_src_data;                                                                                         // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [15:0] id_router_017_src_channel;                                                                                      // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                        // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_015_src4_ready;                                                                                  // led_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src4_ready
	wire          id_router_018_src_endofpacket;                                                                                  // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                                        // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                                // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire   [68:0] id_router_018_src_data;                                                                                         // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [15:0] id_router_018_src_channel;                                                                                      // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                                        // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_015_src5_ready;                                                                                  // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src5_ready
	wire          id_router_019_src_endofpacket;                                                                                  // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                                        // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                                // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire   [68:0] id_router_019_src_data;                                                                                         // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [15:0] id_router_019_src_channel;                                                                                      // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                                        // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          crosser_006_out_ready;                                                                                          // pll_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_006:out_ready
	wire          id_router_020_src_endofpacket;                                                                                  // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                                        // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                                // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire   [68:0] id_router_020_src_data;                                                                                         // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [15:0] id_router_020_src_channel;                                                                                      // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                                        // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          cmd_xbar_demux_015_src7_ready;                                                                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src7_ready
	wire          id_router_021_src_endofpacket;                                                                                  // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire          id_router_021_src_valid;                                                                                        // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire          id_router_021_src_startofpacket;                                                                                // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire   [68:0] id_router_021_src_data;                                                                                         // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire   [15:0] id_router_021_src_channel;                                                                                      // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire          id_router_021_src_ready;                                                                                        // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire          cmd_xbar_demux_015_src8_ready;                                                                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src8_ready
	wire          id_router_022_src_endofpacket;                                                                                  // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire          id_router_022_src_valid;                                                                                        // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire          id_router_022_src_startofpacket;                                                                                // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire   [68:0] id_router_022_src_data;                                                                                         // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire   [15:0] id_router_022_src_channel;                                                                                      // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire          id_router_022_src_ready;                                                                                        // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire          cmd_xbar_demux_015_src9_ready;                                                                                  // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src9_ready
	wire          id_router_023_src_endofpacket;                                                                                  // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire          id_router_023_src_valid;                                                                                        // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire          id_router_023_src_startofpacket;                                                                                // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire   [68:0] id_router_023_src_data;                                                                                         // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire   [15:0] id_router_023_src_channel;                                                                                      // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire          id_router_023_src_ready;                                                                                        // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire          cmd_xbar_demux_015_src10_ready;                                                                                 // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src10_ready
	wire          id_router_024_src_endofpacket;                                                                                  // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire          id_router_024_src_valid;                                                                                        // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire          id_router_024_src_startofpacket;                                                                                // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire   [68:0] id_router_024_src_data;                                                                                         // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire   [15:0] id_router_024_src_channel;                                                                                      // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire          id_router_024_src_ready;                                                                                        // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire          cmd_xbar_demux_015_src11_ready;                                                                                 // lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src11_ready
	wire          id_router_025_src_endofpacket;                                                                                  // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire          id_router_025_src_valid;                                                                                        // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire          id_router_025_src_startofpacket;                                                                                // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire   [68:0] id_router_025_src_data;                                                                                         // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire   [15:0] id_router_025_src_channel;                                                                                      // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire          id_router_025_src_ready;                                                                                        // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire          cmd_xbar_demux_015_src12_ready;                                                                                 // pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src12_ready
	wire          id_router_026_src_endofpacket;                                                                                  // id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire          id_router_026_src_valid;                                                                                        // id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	wire          id_router_026_src_startofpacket;                                                                                // id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire   [68:0] id_router_026_src_data;                                                                                         // id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	wire   [15:0] id_router_026_src_channel;                                                                                      // id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	wire          id_router_026_src_ready;                                                                                        // rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	wire          cmd_xbar_demux_015_src13_ready;                                                                                 // pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src13_ready
	wire          id_router_027_src_endofpacket;                                                                                  // id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire          id_router_027_src_valid;                                                                                        // id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	wire          id_router_027_src_startofpacket;                                                                                // id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire   [68:0] id_router_027_src_data;                                                                                         // id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	wire   [15:0] id_router_027_src_channel;                                                                                      // id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	wire          id_router_027_src_ready;                                                                                        // rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	wire          cmd_xbar_demux_015_src14_ready;                                                                                 // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src14_ready
	wire          id_router_028_src_endofpacket;                                                                                  // id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire          id_router_028_src_valid;                                                                                        // id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	wire          id_router_028_src_startofpacket;                                                                                // id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire   [68:0] id_router_028_src_data;                                                                                         // id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	wire   [15:0] id_router_028_src_channel;                                                                                      // id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	wire          id_router_028_src_ready;                                                                                        // rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	wire          cmd_xbar_demux_015_src15_ready;                                                                                 // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_015:src15_ready
	wire          id_router_029_src_endofpacket;                                                                                  // id_router_029:src_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	wire          id_router_029_src_valid;                                                                                        // id_router_029:src_valid -> rsp_xbar_demux_029:sink_valid
	wire          id_router_029_src_startofpacket;                                                                                // id_router_029:src_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	wire   [68:0] id_router_029_src_data;                                                                                         // id_router_029:src_data -> rsp_xbar_demux_029:sink_data
	wire   [15:0] id_router_029_src_channel;                                                                                      // id_router_029:src_channel -> rsp_xbar_demux_029:sink_channel
	wire          id_router_029_src_ready;                                                                                        // rsp_xbar_demux_029:sink_ready -> id_router_029:src_ready
	wire          cmd_xbar_demux_016_src0_endofpacket;                                                                            // cmd_xbar_demux_016:src0_endofpacket -> cmd_xbar_mux_030:sink0_endofpacket
	wire          cmd_xbar_demux_016_src0_valid;                                                                                  // cmd_xbar_demux_016:src0_valid -> cmd_xbar_mux_030:sink0_valid
	wire          cmd_xbar_demux_016_src0_startofpacket;                                                                          // cmd_xbar_demux_016:src0_startofpacket -> cmd_xbar_mux_030:sink0_startofpacket
	wire   [84:0] cmd_xbar_demux_016_src0_data;                                                                                   // cmd_xbar_demux_016:src0_data -> cmd_xbar_mux_030:sink0_data
	wire    [1:0] cmd_xbar_demux_016_src0_channel;                                                                                // cmd_xbar_demux_016:src0_channel -> cmd_xbar_mux_030:sink0_channel
	wire          cmd_xbar_demux_016_src0_ready;                                                                                  // cmd_xbar_mux_030:sink0_ready -> cmd_xbar_demux_016:src0_ready
	wire          cmd_xbar_demux_017_src0_endofpacket;                                                                            // cmd_xbar_demux_017:src0_endofpacket -> cmd_xbar_mux_030:sink1_endofpacket
	wire          cmd_xbar_demux_017_src0_valid;                                                                                  // cmd_xbar_demux_017:src0_valid -> cmd_xbar_mux_030:sink1_valid
	wire          cmd_xbar_demux_017_src0_startofpacket;                                                                          // cmd_xbar_demux_017:src0_startofpacket -> cmd_xbar_mux_030:sink1_startofpacket
	wire   [84:0] cmd_xbar_demux_017_src0_data;                                                                                   // cmd_xbar_demux_017:src0_data -> cmd_xbar_mux_030:sink1_data
	wire    [1:0] cmd_xbar_demux_017_src0_channel;                                                                                // cmd_xbar_demux_017:src0_channel -> cmd_xbar_mux_030:sink1_channel
	wire          cmd_xbar_demux_017_src0_ready;                                                                                  // cmd_xbar_mux_030:sink1_ready -> cmd_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_030_src0_endofpacket;                                                                            // rsp_xbar_demux_030:src0_endofpacket -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_030_src0_valid;                                                                                  // rsp_xbar_demux_030:src0_valid -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_030_src0_startofpacket;                                                                          // rsp_xbar_demux_030:src0_startofpacket -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [84:0] rsp_xbar_demux_030_src0_data;                                                                                   // rsp_xbar_demux_030:src0_data -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] rsp_xbar_demux_030_src0_channel;                                                                                // rsp_xbar_demux_030:src0_channel -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_030_src1_endofpacket;                                                                            // rsp_xbar_demux_030:src1_endofpacket -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_030_src1_valid;                                                                                  // rsp_xbar_demux_030:src1_valid -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_030_src1_startofpacket;                                                                          // rsp_xbar_demux_030:src1_startofpacket -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [84:0] rsp_xbar_demux_030_src1_data;                                                                                   // rsp_xbar_demux_030:src1_data -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] rsp_xbar_demux_030_src1_channel;                                                                                // rsp_xbar_demux_030:src1_channel -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_016_src_endofpacket;                                                                                // addr_router_016:src_endofpacket -> cmd_xbar_demux_016:sink_endofpacket
	wire          addr_router_016_src_valid;                                                                                      // addr_router_016:src_valid -> cmd_xbar_demux_016:sink_valid
	wire          addr_router_016_src_startofpacket;                                                                              // addr_router_016:src_startofpacket -> cmd_xbar_demux_016:sink_startofpacket
	wire   [84:0] addr_router_016_src_data;                                                                                       // addr_router_016:src_data -> cmd_xbar_demux_016:sink_data
	wire    [1:0] addr_router_016_src_channel;                                                                                    // addr_router_016:src_channel -> cmd_xbar_demux_016:sink_channel
	wire          addr_router_016_src_ready;                                                                                      // cmd_xbar_demux_016:sink_ready -> addr_router_016:src_ready
	wire          rsp_xbar_demux_030_src0_ready;                                                                                  // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_030:src0_ready
	wire          addr_router_017_src_endofpacket;                                                                                // addr_router_017:src_endofpacket -> cmd_xbar_demux_017:sink_endofpacket
	wire          addr_router_017_src_valid;                                                                                      // addr_router_017:src_valid -> cmd_xbar_demux_017:sink_valid
	wire          addr_router_017_src_startofpacket;                                                                              // addr_router_017:src_startofpacket -> cmd_xbar_demux_017:sink_startofpacket
	wire   [84:0] addr_router_017_src_data;                                                                                       // addr_router_017:src_data -> cmd_xbar_demux_017:sink_data
	wire    [1:0] addr_router_017_src_channel;                                                                                    // addr_router_017:src_channel -> cmd_xbar_demux_017:sink_channel
	wire          addr_router_017_src_ready;                                                                                      // cmd_xbar_demux_017:sink_ready -> addr_router_017:src_ready
	wire          rsp_xbar_demux_030_src1_ready;                                                                                  // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_030:src1_ready
	wire          cmd_xbar_mux_030_src_endofpacket;                                                                               // cmd_xbar_mux_030:src_endofpacket -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_030_src_valid;                                                                                     // cmd_xbar_mux_030:src_valid -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_030_src_startofpacket;                                                                             // cmd_xbar_mux_030:src_startofpacket -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_mux_030_src_data;                                                                                      // cmd_xbar_mux_030:src_data -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [1:0] cmd_xbar_mux_030_src_channel;                                                                                   // cmd_xbar_mux_030:src_channel -> tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_030_src_ready;                                                                                     // tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_030:src_ready
	wire          id_router_030_src_endofpacket;                                                                                  // id_router_030:src_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	wire          id_router_030_src_valid;                                                                                        // id_router_030:src_valid -> rsp_xbar_demux_030:sink_valid
	wire          id_router_030_src_startofpacket;                                                                                // id_router_030:src_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	wire   [84:0] id_router_030_src_data;                                                                                         // id_router_030:src_data -> rsp_xbar_demux_030:sink_data
	wire    [1:0] id_router_030_src_channel;                                                                                      // id_router_030:src_channel -> rsp_xbar_demux_030:sink_channel
	wire          id_router_030_src_ready;                                                                                        // rsp_xbar_demux_030:sink_ready -> id_router_030:src_ready
	wire          cmd_xbar_demux_018_src0_endofpacket;                                                                            // cmd_xbar_demux_018:src0_endofpacket -> width_adapter_010:in_endofpacket
	wire          cmd_xbar_demux_018_src0_valid;                                                                                  // cmd_xbar_demux_018:src0_valid -> width_adapter_010:in_valid
	wire          cmd_xbar_demux_018_src0_startofpacket;                                                                          // cmd_xbar_demux_018:src0_startofpacket -> width_adapter_010:in_startofpacket
	wire   [79:0] cmd_xbar_demux_018_src0_data;                                                                                   // cmd_xbar_demux_018:src0_data -> width_adapter_010:in_data
	wire    [1:0] cmd_xbar_demux_018_src0_channel;                                                                                // cmd_xbar_demux_018:src0_channel -> width_adapter_010:in_channel
	wire          cmd_xbar_demux_018_src1_endofpacket;                                                                            // cmd_xbar_demux_018:src1_endofpacket -> max2_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_018_src1_valid;                                                                                  // cmd_xbar_demux_018:src1_valid -> max2_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_018_src1_startofpacket;                                                                          // cmd_xbar_demux_018:src1_startofpacket -> max2_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [79:0] cmd_xbar_demux_018_src1_data;                                                                                   // cmd_xbar_demux_018:src1_data -> max2_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire    [1:0] cmd_xbar_demux_018_src1_channel;                                                                                // cmd_xbar_demux_018:src1_channel -> max2_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_031_src0_endofpacket;                                                                            // rsp_xbar_demux_031:src0_endofpacket -> rsp_xbar_mux_018:sink0_endofpacket
	wire          rsp_xbar_demux_031_src0_valid;                                                                                  // rsp_xbar_demux_031:src0_valid -> rsp_xbar_mux_018:sink0_valid
	wire          rsp_xbar_demux_031_src0_startofpacket;                                                                          // rsp_xbar_demux_031:src0_startofpacket -> rsp_xbar_mux_018:sink0_startofpacket
	wire   [79:0] rsp_xbar_demux_031_src0_data;                                                                                   // rsp_xbar_demux_031:src0_data -> rsp_xbar_mux_018:sink0_data
	wire    [1:0] rsp_xbar_demux_031_src0_channel;                                                                                // rsp_xbar_demux_031:src0_channel -> rsp_xbar_mux_018:sink0_channel
	wire          rsp_xbar_demux_031_src0_ready;                                                                                  // rsp_xbar_mux_018:sink0_ready -> rsp_xbar_demux_031:src0_ready
	wire          rsp_xbar_demux_032_src0_endofpacket;                                                                            // rsp_xbar_demux_032:src0_endofpacket -> rsp_xbar_mux_018:sink1_endofpacket
	wire          rsp_xbar_demux_032_src0_valid;                                                                                  // rsp_xbar_demux_032:src0_valid -> rsp_xbar_mux_018:sink1_valid
	wire          rsp_xbar_demux_032_src0_startofpacket;                                                                          // rsp_xbar_demux_032:src0_startofpacket -> rsp_xbar_mux_018:sink1_startofpacket
	wire   [79:0] rsp_xbar_demux_032_src0_data;                                                                                   // rsp_xbar_demux_032:src0_data -> rsp_xbar_mux_018:sink1_data
	wire    [1:0] rsp_xbar_demux_032_src0_channel;                                                                                // rsp_xbar_demux_032:src0_channel -> rsp_xbar_mux_018:sink1_channel
	wire          rsp_xbar_demux_032_src0_ready;                                                                                  // rsp_xbar_mux_018:sink1_ready -> rsp_xbar_demux_032:src0_ready
	wire          limiter_013_cmd_src_endofpacket;                                                                                // limiter_013:cmd_src_endofpacket -> cmd_xbar_demux_018:sink_endofpacket
	wire          limiter_013_cmd_src_startofpacket;                                                                              // limiter_013:cmd_src_startofpacket -> cmd_xbar_demux_018:sink_startofpacket
	wire   [79:0] limiter_013_cmd_src_data;                                                                                       // limiter_013:cmd_src_data -> cmd_xbar_demux_018:sink_data
	wire    [1:0] limiter_013_cmd_src_channel;                                                                                    // limiter_013:cmd_src_channel -> cmd_xbar_demux_018:sink_channel
	wire          limiter_013_cmd_src_ready;                                                                                      // cmd_xbar_demux_018:sink_ready -> limiter_013:cmd_src_ready
	wire          rsp_xbar_mux_018_src_endofpacket;                                                                               // rsp_xbar_mux_018:src_endofpacket -> limiter_013:rsp_sink_endofpacket
	wire          rsp_xbar_mux_018_src_valid;                                                                                     // rsp_xbar_mux_018:src_valid -> limiter_013:rsp_sink_valid
	wire          rsp_xbar_mux_018_src_startofpacket;                                                                             // rsp_xbar_mux_018:src_startofpacket -> limiter_013:rsp_sink_startofpacket
	wire   [79:0] rsp_xbar_mux_018_src_data;                                                                                      // rsp_xbar_mux_018:src_data -> limiter_013:rsp_sink_data
	wire    [1:0] rsp_xbar_mux_018_src_channel;                                                                                   // rsp_xbar_mux_018:src_channel -> limiter_013:rsp_sink_channel
	wire          rsp_xbar_mux_018_src_ready;                                                                                     // limiter_013:rsp_sink_ready -> rsp_xbar_mux_018:src_ready
	wire          cmd_xbar_demux_018_src1_ready;                                                                                  // max2_uas_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_018:src1_ready
	wire          id_router_032_src_endofpacket;                                                                                  // id_router_032:src_endofpacket -> rsp_xbar_demux_032:sink_endofpacket
	wire          id_router_032_src_valid;                                                                                        // id_router_032:src_valid -> rsp_xbar_demux_032:sink_valid
	wire          id_router_032_src_startofpacket;                                                                                // id_router_032:src_startofpacket -> rsp_xbar_demux_032:sink_startofpacket
	wire   [79:0] id_router_032_src_data;                                                                                         // id_router_032:src_data -> rsp_xbar_demux_032:sink_data
	wire    [1:0] id_router_032_src_channel;                                                                                      // id_router_032:src_channel -> rsp_xbar_demux_032:sink_channel
	wire          id_router_032_src_ready;                                                                                        // rsp_xbar_demux_032:sink_ready -> id_router_032:src_ready
	wire          cmd_xbar_demux_006_src0_endofpacket;                                                                            // cmd_xbar_demux_006:src0_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_006_src0_valid;                                                                                  // cmd_xbar_demux_006:src0_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_006_src0_startofpacket;                                                                          // cmd_xbar_demux_006:src0_startofpacket -> width_adapter:in_startofpacket
	wire   [88:0] cmd_xbar_demux_006_src0_data;                                                                                   // cmd_xbar_demux_006:src0_data -> width_adapter:in_data
	wire    [5:0] cmd_xbar_demux_006_src0_channel;                                                                                // cmd_xbar_demux_006:src0_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_006_src0_ready;                                                                                  // width_adapter:in_ready -> cmd_xbar_demux_006:src0_ready
	wire          width_adapter_src_endofpacket;                                                                                  // width_adapter:out_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                        // width_adapter:out_valid -> cmd_xbar_mux_010:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                                // width_adapter:out_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [124:0] width_adapter_src_data;                                                                                         // width_adapter:out_data -> cmd_xbar_mux_010:sink0_data
	wire          width_adapter_src_ready;                                                                                        // cmd_xbar_mux_010:sink0_ready -> width_adapter:out_ready
	wire    [5:0] width_adapter_src_channel;                                                                                      // width_adapter:out_channel -> cmd_xbar_mux_010:sink0_channel
	wire          cmd_xbar_demux_007_src0_endofpacket;                                                                            // cmd_xbar_demux_007:src0_endofpacket -> width_adapter_001:in_endofpacket
	wire          cmd_xbar_demux_007_src0_valid;                                                                                  // cmd_xbar_demux_007:src0_valid -> width_adapter_001:in_valid
	wire          cmd_xbar_demux_007_src0_startofpacket;                                                                          // cmd_xbar_demux_007:src0_startofpacket -> width_adapter_001:in_startofpacket
	wire   [88:0] cmd_xbar_demux_007_src0_data;                                                                                   // cmd_xbar_demux_007:src0_data -> width_adapter_001:in_data
	wire    [5:0] cmd_xbar_demux_007_src0_channel;                                                                                // cmd_xbar_demux_007:src0_channel -> width_adapter_001:in_channel
	wire          cmd_xbar_demux_007_src0_ready;                                                                                  // width_adapter_001:in_ready -> cmd_xbar_demux_007:src0_ready
	wire          width_adapter_001_src_endofpacket;                                                                              // width_adapter_001:out_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire          width_adapter_001_src_valid;                                                                                    // width_adapter_001:out_valid -> cmd_xbar_mux_010:sink1_valid
	wire          width_adapter_001_src_startofpacket;                                                                            // width_adapter_001:out_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [124:0] width_adapter_001_src_data;                                                                                     // width_adapter_001:out_data -> cmd_xbar_mux_010:sink1_data
	wire          width_adapter_001_src_ready;                                                                                    // cmd_xbar_mux_010:sink1_ready -> width_adapter_001:out_ready
	wire    [5:0] width_adapter_001_src_channel;                                                                                  // width_adapter_001:out_channel -> cmd_xbar_mux_010:sink1_channel
	wire          cmd_xbar_demux_010_src0_endofpacket;                                                                            // cmd_xbar_demux_010:src0_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_010_src0_valid;                                                                                  // cmd_xbar_demux_010:src0_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_010_src0_startofpacket;                                                                          // cmd_xbar_demux_010:src0_startofpacket -> width_adapter_002:in_startofpacket
	wire   [88:0] cmd_xbar_demux_010_src0_data;                                                                                   // cmd_xbar_demux_010:src0_data -> width_adapter_002:in_data
	wire    [5:0] cmd_xbar_demux_010_src0_channel;                                                                                // cmd_xbar_demux_010:src0_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_010_src0_ready;                                                                                  // width_adapter_002:in_ready -> cmd_xbar_demux_010:src0_ready
	wire          width_adapter_002_src_endofpacket;                                                                              // width_adapter_002:out_endofpacket -> cmd_xbar_mux_010:sink4_endofpacket
	wire          width_adapter_002_src_valid;                                                                                    // width_adapter_002:out_valid -> cmd_xbar_mux_010:sink4_valid
	wire          width_adapter_002_src_startofpacket;                                                                            // width_adapter_002:out_startofpacket -> cmd_xbar_mux_010:sink4_startofpacket
	wire  [124:0] width_adapter_002_src_data;                                                                                     // width_adapter_002:out_data -> cmd_xbar_mux_010:sink4_data
	wire          width_adapter_002_src_ready;                                                                                    // cmd_xbar_mux_010:sink4_ready -> width_adapter_002:out_ready
	wire    [5:0] width_adapter_002_src_channel;                                                                                  // width_adapter_002:out_channel -> cmd_xbar_mux_010:sink4_channel
	wire          cmd_xbar_demux_011_src0_endofpacket;                                                                            // cmd_xbar_demux_011:src0_endofpacket -> width_adapter_003:in_endofpacket
	wire          cmd_xbar_demux_011_src0_valid;                                                                                  // cmd_xbar_demux_011:src0_valid -> width_adapter_003:in_valid
	wire          cmd_xbar_demux_011_src0_startofpacket;                                                                          // cmd_xbar_demux_011:src0_startofpacket -> width_adapter_003:in_startofpacket
	wire   [88:0] cmd_xbar_demux_011_src0_data;                                                                                   // cmd_xbar_demux_011:src0_data -> width_adapter_003:in_data
	wire    [5:0] cmd_xbar_demux_011_src0_channel;                                                                                // cmd_xbar_demux_011:src0_channel -> width_adapter_003:in_channel
	wire          cmd_xbar_demux_011_src0_ready;                                                                                  // width_adapter_003:in_ready -> cmd_xbar_demux_011:src0_ready
	wire          width_adapter_003_src_endofpacket;                                                                              // width_adapter_003:out_endofpacket -> cmd_xbar_mux_010:sink5_endofpacket
	wire          width_adapter_003_src_valid;                                                                                    // width_adapter_003:out_valid -> cmd_xbar_mux_010:sink5_valid
	wire          width_adapter_003_src_startofpacket;                                                                            // width_adapter_003:out_startofpacket -> cmd_xbar_mux_010:sink5_startofpacket
	wire  [124:0] width_adapter_003_src_data;                                                                                     // width_adapter_003:out_data -> cmd_xbar_mux_010:sink5_data
	wire          width_adapter_003_src_ready;                                                                                    // cmd_xbar_mux_010:sink5_ready -> width_adapter_003:out_ready
	wire    [5:0] width_adapter_003_src_channel;                                                                                  // width_adapter_003:out_channel -> cmd_xbar_mux_010:sink5_channel
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                            // rsp_xbar_demux_010:src0_endofpacket -> width_adapter_004:in_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                  // rsp_xbar_demux_010:src0_valid -> width_adapter_004:in_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                          // rsp_xbar_demux_010:src0_startofpacket -> width_adapter_004:in_startofpacket
	wire  [124:0] rsp_xbar_demux_010_src0_data;                                                                                   // rsp_xbar_demux_010:src0_data -> width_adapter_004:in_data
	wire    [5:0] rsp_xbar_demux_010_src0_channel;                                                                                // rsp_xbar_demux_010:src0_channel -> width_adapter_004:in_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                  // width_adapter_004:in_ready -> rsp_xbar_demux_010:src0_ready
	wire          width_adapter_004_src_endofpacket;                                                                              // width_adapter_004:out_endofpacket -> limiter_006:rsp_sink_endofpacket
	wire          width_adapter_004_src_valid;                                                                                    // width_adapter_004:out_valid -> limiter_006:rsp_sink_valid
	wire          width_adapter_004_src_startofpacket;                                                                            // width_adapter_004:out_startofpacket -> limiter_006:rsp_sink_startofpacket
	wire   [88:0] width_adapter_004_src_data;                                                                                     // width_adapter_004:out_data -> limiter_006:rsp_sink_data
	wire    [5:0] width_adapter_004_src_channel;                                                                                  // width_adapter_004:out_channel -> limiter_006:rsp_sink_channel
	wire          rsp_xbar_demux_010_src1_endofpacket;                                                                            // rsp_xbar_demux_010:src1_endofpacket -> width_adapter_005:in_endofpacket
	wire          rsp_xbar_demux_010_src1_valid;                                                                                  // rsp_xbar_demux_010:src1_valid -> width_adapter_005:in_valid
	wire          rsp_xbar_demux_010_src1_startofpacket;                                                                          // rsp_xbar_demux_010:src1_startofpacket -> width_adapter_005:in_startofpacket
	wire  [124:0] rsp_xbar_demux_010_src1_data;                                                                                   // rsp_xbar_demux_010:src1_data -> width_adapter_005:in_data
	wire    [5:0] rsp_xbar_demux_010_src1_channel;                                                                                // rsp_xbar_demux_010:src1_channel -> width_adapter_005:in_channel
	wire          rsp_xbar_demux_010_src1_ready;                                                                                  // width_adapter_005:in_ready -> rsp_xbar_demux_010:src1_ready
	wire          width_adapter_005_src_endofpacket;                                                                              // width_adapter_005:out_endofpacket -> limiter_007:rsp_sink_endofpacket
	wire          width_adapter_005_src_valid;                                                                                    // width_adapter_005:out_valid -> limiter_007:rsp_sink_valid
	wire          width_adapter_005_src_startofpacket;                                                                            // width_adapter_005:out_startofpacket -> limiter_007:rsp_sink_startofpacket
	wire   [88:0] width_adapter_005_src_data;                                                                                     // width_adapter_005:out_data -> limiter_007:rsp_sink_data
	wire    [5:0] width_adapter_005_src_channel;                                                                                  // width_adapter_005:out_channel -> limiter_007:rsp_sink_channel
	wire          rsp_xbar_demux_010_src4_endofpacket;                                                                            // rsp_xbar_demux_010:src4_endofpacket -> width_adapter_006:in_endofpacket
	wire          rsp_xbar_demux_010_src4_valid;                                                                                  // rsp_xbar_demux_010:src4_valid -> width_adapter_006:in_valid
	wire          rsp_xbar_demux_010_src4_startofpacket;                                                                          // rsp_xbar_demux_010:src4_startofpacket -> width_adapter_006:in_startofpacket
	wire  [124:0] rsp_xbar_demux_010_src4_data;                                                                                   // rsp_xbar_demux_010:src4_data -> width_adapter_006:in_data
	wire    [5:0] rsp_xbar_demux_010_src4_channel;                                                                                // rsp_xbar_demux_010:src4_channel -> width_adapter_006:in_channel
	wire          rsp_xbar_demux_010_src4_ready;                                                                                  // width_adapter_006:in_ready -> rsp_xbar_demux_010:src4_ready
	wire          width_adapter_006_src_endofpacket;                                                                              // width_adapter_006:out_endofpacket -> rsp_xbar_mux_010:sink0_endofpacket
	wire          width_adapter_006_src_valid;                                                                                    // width_adapter_006:out_valid -> rsp_xbar_mux_010:sink0_valid
	wire          width_adapter_006_src_startofpacket;                                                                            // width_adapter_006:out_startofpacket -> rsp_xbar_mux_010:sink0_startofpacket
	wire   [88:0] width_adapter_006_src_data;                                                                                     // width_adapter_006:out_data -> rsp_xbar_mux_010:sink0_data
	wire          width_adapter_006_src_ready;                                                                                    // rsp_xbar_mux_010:sink0_ready -> width_adapter_006:out_ready
	wire    [5:0] width_adapter_006_src_channel;                                                                                  // width_adapter_006:out_channel -> rsp_xbar_mux_010:sink0_channel
	wire          rsp_xbar_demux_010_src5_endofpacket;                                                                            // rsp_xbar_demux_010:src5_endofpacket -> width_adapter_007:in_endofpacket
	wire          rsp_xbar_demux_010_src5_valid;                                                                                  // rsp_xbar_demux_010:src5_valid -> width_adapter_007:in_valid
	wire          rsp_xbar_demux_010_src5_startofpacket;                                                                          // rsp_xbar_demux_010:src5_startofpacket -> width_adapter_007:in_startofpacket
	wire  [124:0] rsp_xbar_demux_010_src5_data;                                                                                   // rsp_xbar_demux_010:src5_data -> width_adapter_007:in_data
	wire    [5:0] rsp_xbar_demux_010_src5_channel;                                                                                // rsp_xbar_demux_010:src5_channel -> width_adapter_007:in_channel
	wire          rsp_xbar_demux_010_src5_ready;                                                                                  // width_adapter_007:in_ready -> rsp_xbar_demux_010:src5_ready
	wire          width_adapter_007_src_endofpacket;                                                                              // width_adapter_007:out_endofpacket -> limiter_011:rsp_sink_endofpacket
	wire          width_adapter_007_src_valid;                                                                                    // width_adapter_007:out_valid -> limiter_011:rsp_sink_valid
	wire          width_adapter_007_src_startofpacket;                                                                            // width_adapter_007:out_startofpacket -> limiter_011:rsp_sink_startofpacket
	wire   [88:0] width_adapter_007_src_data;                                                                                     // width_adapter_007:out_data -> limiter_011:rsp_sink_data
	wire    [5:0] width_adapter_007_src_channel;                                                                                  // width_adapter_007:out_channel -> limiter_011:rsp_sink_channel
	wire          cmd_xbar_mux_012_src_endofpacket;                                                                               // cmd_xbar_mux_012:src_endofpacket -> width_adapter_008:in_endofpacket
	wire          cmd_xbar_mux_012_src_valid;                                                                                     // cmd_xbar_mux_012:src_valid -> width_adapter_008:in_valid
	wire          cmd_xbar_mux_012_src_startofpacket;                                                                             // cmd_xbar_mux_012:src_startofpacket -> width_adapter_008:in_startofpacket
	wire   [86:0] cmd_xbar_mux_012_src_data;                                                                                      // cmd_xbar_mux_012:src_data -> width_adapter_008:in_data
	wire    [1:0] cmd_xbar_mux_012_src_channel;                                                                                   // cmd_xbar_mux_012:src_channel -> width_adapter_008:in_channel
	wire          cmd_xbar_mux_012_src_ready;                                                                                     // width_adapter_008:in_ready -> cmd_xbar_mux_012:src_ready
	wire          width_adapter_008_src_endofpacket;                                                                              // width_adapter_008:out_endofpacket -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          width_adapter_008_src_valid;                                                                                    // width_adapter_008:out_valid -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          width_adapter_008_src_startofpacket;                                                                            // width_adapter_008:out_startofpacket -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [122:0] width_adapter_008_src_data;                                                                                     // width_adapter_008:out_data -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire          width_adapter_008_src_ready;                                                                                    // sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_008:out_ready
	wire    [1:0] width_adapter_008_src_channel;                                                                                  // width_adapter_008:out_channel -> sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          id_router_012_src_endofpacket;                                                                                  // id_router_012:src_endofpacket -> width_adapter_009:in_endofpacket
	wire          id_router_012_src_valid;                                                                                        // id_router_012:src_valid -> width_adapter_009:in_valid
	wire          id_router_012_src_startofpacket;                                                                                // id_router_012:src_startofpacket -> width_adapter_009:in_startofpacket
	wire  [122:0] id_router_012_src_data;                                                                                         // id_router_012:src_data -> width_adapter_009:in_data
	wire    [1:0] id_router_012_src_channel;                                                                                      // id_router_012:src_channel -> width_adapter_009:in_channel
	wire          id_router_012_src_ready;                                                                                        // width_adapter_009:in_ready -> id_router_012:src_ready
	wire          width_adapter_009_src_endofpacket;                                                                              // width_adapter_009:out_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          width_adapter_009_src_valid;                                                                                    // width_adapter_009:out_valid -> rsp_xbar_demux_012:sink_valid
	wire          width_adapter_009_src_startofpacket;                                                                            // width_adapter_009:out_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire   [86:0] width_adapter_009_src_data;                                                                                     // width_adapter_009:out_data -> rsp_xbar_demux_012:sink_data
	wire          width_adapter_009_src_ready;                                                                                    // rsp_xbar_demux_012:sink_ready -> width_adapter_009:out_ready
	wire    [1:0] width_adapter_009_src_channel;                                                                                  // width_adapter_009:out_channel -> rsp_xbar_demux_012:sink_channel
	wire          cmd_xbar_demux_018_src0_ready;                                                                                  // width_adapter_010:in_ready -> cmd_xbar_demux_018:src0_ready
	wire          width_adapter_010_src_endofpacket;                                                                              // width_adapter_010:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_010_src_valid;                                                                                    // width_adapter_010:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_010_src_startofpacket;                                                                            // width_adapter_010:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [61:0] width_adapter_010_src_data;                                                                                     // width_adapter_010:out_data -> burst_adapter:sink0_data
	wire          width_adapter_010_src_ready;                                                                                    // burst_adapter:sink0_ready -> width_adapter_010:out_ready
	wire    [1:0] width_adapter_010_src_channel;                                                                                  // width_adapter_010:out_channel -> burst_adapter:sink0_channel
	wire          id_router_031_src_endofpacket;                                                                                  // id_router_031:src_endofpacket -> width_adapter_011:in_endofpacket
	wire          id_router_031_src_valid;                                                                                        // id_router_031:src_valid -> width_adapter_011:in_valid
	wire          id_router_031_src_startofpacket;                                                                                // id_router_031:src_startofpacket -> width_adapter_011:in_startofpacket
	wire   [61:0] id_router_031_src_data;                                                                                         // id_router_031:src_data -> width_adapter_011:in_data
	wire    [1:0] id_router_031_src_channel;                                                                                      // id_router_031:src_channel -> width_adapter_011:in_channel
	wire          id_router_031_src_ready;                                                                                        // width_adapter_011:in_ready -> id_router_031:src_ready
	wire          width_adapter_011_src_endofpacket;                                                                              // width_adapter_011:out_endofpacket -> rsp_xbar_demux_031:sink_endofpacket
	wire          width_adapter_011_src_valid;                                                                                    // width_adapter_011:out_valid -> rsp_xbar_demux_031:sink_valid
	wire          width_adapter_011_src_startofpacket;                                                                            // width_adapter_011:out_startofpacket -> rsp_xbar_demux_031:sink_startofpacket
	wire   [79:0] width_adapter_011_src_data;                                                                                     // width_adapter_011:out_data -> rsp_xbar_demux_031:sink_data
	wire          width_adapter_011_src_ready;                                                                                    // rsp_xbar_demux_031:sink_ready -> width_adapter_011:out_ready
	wire    [1:0] width_adapter_011_src_channel;                                                                                  // width_adapter_011:out_channel -> rsp_xbar_demux_031:sink_channel
	wire          crosser_out_endofpacket;                                                                                        // crosser:out_endofpacket -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                              // crosser:out_valid -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                                      // crosser:out_startofpacket -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] crosser_out_data;                                                                                               // crosser:out_data -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:cp_data
	wire    [9:0] crosser_out_channel;                                                                                            // crosser:out_channel -> sls_sdhc_control_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src5_endofpacket;                                                                                // cmd_xbar_demux:src5_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_src5_valid;                                                                                      // cmd_xbar_demux:src5_valid -> crosser:in_valid
	wire          cmd_xbar_demux_src5_startofpacket;                                                                              // cmd_xbar_demux:src5_startofpacket -> crosser:in_startofpacket
	wire   [88:0] cmd_xbar_demux_src5_data;                                                                                       // cmd_xbar_demux:src5_data -> crosser:in_data
	wire    [9:0] cmd_xbar_demux_src5_channel;                                                                                    // cmd_xbar_demux:src5_channel -> crosser:in_channel
	wire          cmd_xbar_demux_src5_ready;                                                                                      // crosser:in_ready -> cmd_xbar_demux:src5_ready
	wire          crosser_001_out_endofpacket;                                                                                    // crosser_001:out_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire          crosser_001_out_valid;                                                                                          // crosser_001:out_valid -> rsp_xbar_mux:sink5_valid
	wire          crosser_001_out_startofpacket;                                                                                  // crosser_001:out_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire   [88:0] crosser_001_out_data;                                                                                           // crosser_001:out_data -> rsp_xbar_mux:sink5_data
	wire    [9:0] crosser_001_out_channel;                                                                                        // crosser_001:out_channel -> rsp_xbar_mux:sink5_channel
	wire          crosser_001_out_ready;                                                                                          // rsp_xbar_mux:sink5_ready -> crosser_001:out_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                            // rsp_xbar_demux_005:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                  // rsp_xbar_demux_005:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                          // rsp_xbar_demux_005:src0_startofpacket -> crosser_001:in_startofpacket
	wire   [88:0] rsp_xbar_demux_005_src0_data;                                                                                   // rsp_xbar_demux_005:src0_data -> crosser_001:in_data
	wire    [9:0] rsp_xbar_demux_005_src0_channel;                                                                                // rsp_xbar_demux_005:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                  // crosser_001:in_ready -> rsp_xbar_demux_005:src0_ready
	wire          crosser_002_out_endofpacket;                                                                                    // crosser_002:out_endofpacket -> cmd_xbar_mux_012:sink0_endofpacket
	wire          crosser_002_out_valid;                                                                                          // crosser_002:out_valid -> cmd_xbar_mux_012:sink0_valid
	wire          crosser_002_out_startofpacket;                                                                                  // crosser_002:out_startofpacket -> cmd_xbar_mux_012:sink0_startofpacket
	wire   [86:0] crosser_002_out_data;                                                                                           // crosser_002:out_data -> cmd_xbar_mux_012:sink0_data
	wire    [1:0] crosser_002_out_channel;                                                                                        // crosser_002:out_channel -> cmd_xbar_mux_012:sink0_channel
	wire          crosser_002_out_ready;                                                                                          // cmd_xbar_mux_012:sink0_ready -> crosser_002:out_ready
	wire          cmd_xbar_demux_012_src0_endofpacket;                                                                            // cmd_xbar_demux_012:src0_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_012_src0_valid;                                                                                  // cmd_xbar_demux_012:src0_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_012_src0_startofpacket;                                                                          // cmd_xbar_demux_012:src0_startofpacket -> crosser_002:in_startofpacket
	wire   [86:0] cmd_xbar_demux_012_src0_data;                                                                                   // cmd_xbar_demux_012:src0_data -> crosser_002:in_data
	wire    [1:0] cmd_xbar_demux_012_src0_channel;                                                                                // cmd_xbar_demux_012:src0_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_012_src0_ready;                                                                                  // crosser_002:in_ready -> cmd_xbar_demux_012:src0_ready
	wire          crosser_003_out_endofpacket;                                                                                    // crosser_003:out_endofpacket -> cmd_xbar_mux_012:sink1_endofpacket
	wire          crosser_003_out_valid;                                                                                          // crosser_003:out_valid -> cmd_xbar_mux_012:sink1_valid
	wire          crosser_003_out_startofpacket;                                                                                  // crosser_003:out_startofpacket -> cmd_xbar_mux_012:sink1_startofpacket
	wire   [86:0] crosser_003_out_data;                                                                                           // crosser_003:out_data -> cmd_xbar_mux_012:sink1_data
	wire    [1:0] crosser_003_out_channel;                                                                                        // crosser_003:out_channel -> cmd_xbar_mux_012:sink1_channel
	wire          crosser_003_out_ready;                                                                                          // cmd_xbar_mux_012:sink1_ready -> crosser_003:out_ready
	wire          cmd_xbar_demux_013_src0_endofpacket;                                                                            // cmd_xbar_demux_013:src0_endofpacket -> crosser_003:in_endofpacket
	wire          cmd_xbar_demux_013_src0_valid;                                                                                  // cmd_xbar_demux_013:src0_valid -> crosser_003:in_valid
	wire          cmd_xbar_demux_013_src0_startofpacket;                                                                          // cmd_xbar_demux_013:src0_startofpacket -> crosser_003:in_startofpacket
	wire   [86:0] cmd_xbar_demux_013_src0_data;                                                                                   // cmd_xbar_demux_013:src0_data -> crosser_003:in_data
	wire    [1:0] cmd_xbar_demux_013_src0_channel;                                                                                // cmd_xbar_demux_013:src0_channel -> crosser_003:in_channel
	wire          cmd_xbar_demux_013_src0_ready;                                                                                  // crosser_003:in_ready -> cmd_xbar_demux_013:src0_ready
	wire          crosser_004_out_endofpacket;                                                                                    // crosser_004:out_endofpacket -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_004_out_valid;                                                                                          // crosser_004:out_valid -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_004_out_startofpacket;                                                                                  // crosser_004:out_startofpacket -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [86:0] crosser_004_out_data;                                                                                           // crosser_004:out_data -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] crosser_004_out_channel;                                                                                        // crosser_004:out_channel -> sls_sdhc_read_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                            // rsp_xbar_demux_012:src0_endofpacket -> crosser_004:in_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                  // rsp_xbar_demux_012:src0_valid -> crosser_004:in_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                          // rsp_xbar_demux_012:src0_startofpacket -> crosser_004:in_startofpacket
	wire   [86:0] rsp_xbar_demux_012_src0_data;                                                                                   // rsp_xbar_demux_012:src0_data -> crosser_004:in_data
	wire    [1:0] rsp_xbar_demux_012_src0_channel;                                                                                // rsp_xbar_demux_012:src0_channel -> crosser_004:in_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                                  // crosser_004:in_ready -> rsp_xbar_demux_012:src0_ready
	wire          crosser_005_out_endofpacket;                                                                                    // crosser_005:out_endofpacket -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_005_out_valid;                                                                                          // crosser_005:out_valid -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_005_out_startofpacket;                                                                                  // crosser_005:out_startofpacket -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [86:0] crosser_005_out_data;                                                                                           // crosser_005:out_data -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] crosser_005_out_channel;                                                                                        // crosser_005:out_channel -> sls_sdhc_write_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_012_src1_endofpacket;                                                                            // rsp_xbar_demux_012:src1_endofpacket -> crosser_005:in_endofpacket
	wire          rsp_xbar_demux_012_src1_valid;                                                                                  // rsp_xbar_demux_012:src1_valid -> crosser_005:in_valid
	wire          rsp_xbar_demux_012_src1_startofpacket;                                                                          // rsp_xbar_demux_012:src1_startofpacket -> crosser_005:in_startofpacket
	wire   [86:0] rsp_xbar_demux_012_src1_data;                                                                                   // rsp_xbar_demux_012:src1_data -> crosser_005:in_data
	wire    [1:0] rsp_xbar_demux_012_src1_channel;                                                                                // rsp_xbar_demux_012:src1_channel -> crosser_005:in_channel
	wire          rsp_xbar_demux_012_src1_ready;                                                                                  // crosser_005:in_ready -> rsp_xbar_demux_012:src1_ready
	wire          crosser_006_out_endofpacket;                                                                                    // crosser_006:out_endofpacket -> pll_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_006_out_valid;                                                                                          // crosser_006:out_valid -> pll_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_006_out_startofpacket;                                                                                  // crosser_006:out_startofpacket -> pll_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [68:0] crosser_006_out_data;                                                                                           // crosser_006:out_data -> pll_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_006_out_channel;                                                                                        // crosser_006:out_channel -> pll_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_015_src6_endofpacket;                                                                            // cmd_xbar_demux_015:src6_endofpacket -> crosser_006:in_endofpacket
	wire          cmd_xbar_demux_015_src6_valid;                                                                                  // cmd_xbar_demux_015:src6_valid -> crosser_006:in_valid
	wire          cmd_xbar_demux_015_src6_startofpacket;                                                                          // cmd_xbar_demux_015:src6_startofpacket -> crosser_006:in_startofpacket
	wire   [68:0] cmd_xbar_demux_015_src6_data;                                                                                   // cmd_xbar_demux_015:src6_data -> crosser_006:in_data
	wire   [15:0] cmd_xbar_demux_015_src6_channel;                                                                                // cmd_xbar_demux_015:src6_channel -> crosser_006:in_channel
	wire          cmd_xbar_demux_015_src6_ready;                                                                                  // crosser_006:in_ready -> cmd_xbar_demux_015:src6_ready
	wire          crosser_007_out_endofpacket;                                                                                    // crosser_007:out_endofpacket -> rsp_xbar_mux_015:sink6_endofpacket
	wire          crosser_007_out_valid;                                                                                          // crosser_007:out_valid -> rsp_xbar_mux_015:sink6_valid
	wire          crosser_007_out_startofpacket;                                                                                  // crosser_007:out_startofpacket -> rsp_xbar_mux_015:sink6_startofpacket
	wire   [68:0] crosser_007_out_data;                                                                                           // crosser_007:out_data -> rsp_xbar_mux_015:sink6_data
	wire   [15:0] crosser_007_out_channel;                                                                                        // crosser_007:out_channel -> rsp_xbar_mux_015:sink6_channel
	wire          crosser_007_out_ready;                                                                                          // rsp_xbar_mux_015:sink6_ready -> crosser_007:out_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                                            // rsp_xbar_demux_020:src0_endofpacket -> crosser_007:in_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                                  // rsp_xbar_demux_020:src0_valid -> crosser_007:in_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                                          // rsp_xbar_demux_020:src0_startofpacket -> crosser_007:in_startofpacket
	wire   [68:0] rsp_xbar_demux_020_src0_data;                                                                                   // rsp_xbar_demux_020:src0_data -> crosser_007:in_data
	wire   [15:0] rsp_xbar_demux_020_src0_channel;                                                                                // rsp_xbar_demux_020:src0_channel -> crosser_007:in_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                                  // crosser_007:in_ready -> rsp_xbar_demux_020:src0_ready
	wire    [9:0] limiter_cmd_valid_data;                                                                                         // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire    [9:0] limiter_001_cmd_valid_data;                                                                                     // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire    [9:0] limiter_002_cmd_valid_data;                                                                                     // limiter_002:cmd_src_valid -> cmd_xbar_demux_002:sink_valid
	wire    [9:0] limiter_003_cmd_valid_data;                                                                                     // limiter_003:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire    [9:0] limiter_004_cmd_valid_data;                                                                                     // limiter_004:cmd_src_valid -> cmd_xbar_demux_004:sink_valid
	wire    [9:0] limiter_005_cmd_valid_data;                                                                                     // limiter_005:cmd_src_valid -> cmd_xbar_demux_005:sink_valid
	wire    [5:0] limiter_006_cmd_valid_data;                                                                                     // limiter_006:cmd_src_valid -> cmd_xbar_demux_006:sink_valid
	wire    [5:0] limiter_007_cmd_valid_data;                                                                                     // limiter_007:cmd_src_valid -> cmd_xbar_demux_007:sink_valid
	wire    [5:0] limiter_008_cmd_valid_data;                                                                                     // limiter_008:cmd_src_valid -> cmd_xbar_demux_008:sink_valid
	wire    [5:0] limiter_009_cmd_valid_data;                                                                                     // limiter_009:cmd_src_valid -> cmd_xbar_demux_009:sink_valid
	wire    [5:0] limiter_010_cmd_valid_data;                                                                                     // limiter_010:cmd_src_valid -> cmd_xbar_demux_010:sink_valid
	wire    [5:0] limiter_011_cmd_valid_data;                                                                                     // limiter_011:cmd_src_valid -> cmd_xbar_demux_011:sink_valid
	wire   [15:0] limiter_012_cmd_valid_data;                                                                                     // limiter_012:cmd_src_valid -> cmd_xbar_demux_015:sink_valid
	wire    [1:0] limiter_013_cmd_valid_data;                                                                                     // limiter_013:cmd_src_valid -> cmd_xbar_demux_018:sink_valid
	wire          irq_mapper_receiver4_irq;                                                                                       // sgdma_rx:csr_irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                                                       // sgdma_tx:csr_irq -> irq_mapper:receiver5_irq
	wire   [31:0] cpu_d_irq_irq;                                                                                                  // irq_mapper:sender_irq -> cpu:d_irq
	wire          irq_mapper_receiver0_irq;                                                                                       // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                                  // button_pio:irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver1_irq;                                                                                       // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                                              // high_res_timer:irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver2_irq;                                                                                       // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                                                                              // jtag_uart:av_irq -> irq_synchronizer_002:receiver_irq
	wire          irq_mapper_receiver3_irq;                                                                                       // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_003_receiver_irq;                                                                              // lcd_sgdma:csr_irq -> irq_synchronizer_003:receiver_irq
	wire          irq_mapper_receiver6_irq;                                                                                       // irq_synchronizer_004:sender_irq -> irq_mapper:receiver6_irq
	wire    [0:0] irq_synchronizer_004_receiver_irq;                                                                              // sys_clk_timer:irq -> irq_synchronizer_004:receiver_irq
	wire          irq_mapper_receiver7_irq;                                                                                       // irq_synchronizer_005:sender_irq -> irq_mapper:receiver7_irq
	wire    [0:0] irq_synchronizer_005_receiver_irq;                                                                              // touch_panel_pen_irq_n:irq -> irq_synchronizer_005:receiver_irq
	wire          irq_mapper_receiver8_irq;                                                                                       // irq_synchronizer_006:sender_irq -> irq_mapper:receiver8_irq
	wire    [0:0] irq_synchronizer_006_receiver_irq;                                                                              // touch_panel_spi:irq -> irq_synchronizer_006:receiver_irq
	wire          irq_mapper_receiver9_irq;                                                                                       // irq_synchronizer_007:sender_irq -> irq_mapper:receiver9_irq
	wire    [0:0] irq_synchronizer_007_receiver_irq;                                                                              // uart1:irq -> irq_synchronizer_007:receiver_irq
	wire          irq_mapper_receiver10_irq;                                                                                      // irq_synchronizer_008:sender_irq -> irq_mapper:receiver10_irq
	wire    [0:0] irq_synchronizer_008_receiver_irq;                                                                              // sls_sdhc:AvS_irq -> irq_synchronizer_008:receiver_irq

	application_selector_pll pll (
		.address      (pll_s1_translator_avalon_anti_slave_0_address),    //           s1.address
		.chipselect   (pll_s1_translator_avalon_anti_slave_0_chipselect), //             .chipselect
		.read         (pll_s1_translator_avalon_anti_slave_0_read),       //             .read
		.readdata     (pll_s1_translator_avalon_anti_slave_0_readdata),   //             .readdata
		.write        (pll_s1_translator_avalon_anti_slave_0_write),      //             .write
		.writedata    (pll_s1_translator_avalon_anti_slave_0_writedata),  //             .writedata
		.clk          (clk),                                              //       inclk0.clk
		.reset_n      (~rst_controller_reset_out_reset),                  //        reset.reset_n
		.resetrequest (pll_resetrequest_reset),                           // resetrequest.reset
		.c0           (pll_c0_out),                                       //           c0.clk
		.c2           (pll_c2_out)                                        //           c2.clk
	);

	application_selector_descriptor_memory descriptor_memory (
		.clk        (pll_c0_out),                                                     //   clk1.clk
		.address    (descriptor_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (descriptor_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset)                              // reset1.reset
	);

	application_selector_ddr2_sdram ddr2_sdram (
		.local_address     (ddr2_sdram_s1_translator_avalon_anti_slave_0_address),            //                  s1.address
		.local_write_req   (ddr2_sdram_s1_translator_avalon_anti_slave_0_write),              //                    .write
		.local_read_req    (ddr2_sdram_s1_translator_avalon_anti_slave_0_read),               //                    .read
		.local_burstbegin  (ddr2_sdram_s1_translator_avalon_anti_slave_0_beginbursttransfer), //                    .beginbursttransfer
		.local_ready       (ddr2_sdram_s1_translator_avalon_anti_slave_0_waitrequest),        //                    .waitrequest_n
		.local_rdata       (ddr2_sdram_s1_translator_avalon_anti_slave_0_readdata),           //                    .readdata
		.local_rdata_valid (ddr2_sdram_s1_translator_avalon_anti_slave_0_readdatavalid),      //                    .readdatavalid
		.local_wdata       (ddr2_sdram_s1_translator_avalon_anti_slave_0_writedata),          //                    .writedata
		.local_be          (ddr2_sdram_s1_translator_avalon_anti_slave_0_byteenable),         //                    .byteenable
		.local_size        (ddr2_sdram_s1_translator_avalon_anti_slave_0_burstcount),         //                    .burstcount
		.local_refresh_ack (local_refresh_ack_from_the_ddr2_sdram),                           // external_connection.export
		.local_wdata_req   (local_wdata_req_from_the_ddr2_sdram),                             //                    .export
		.local_init_done   (local_init_done_from_the_ddr2_sdram),                             //                    .export
		.reset_phy_clk_n   (reset_phy_clk_n_from_the_ddr2_sdram),                             //                    .export
		.mem_odt           (mem_odt_from_the_ddr2_sdram),                                     //              memory.mem_odt
		.mem_clk           (mem_clk_to_and_from_the_ddr2_sdram),                              //                    .mem_clk
		.mem_clk_n         (mem_clk_n_to_and_from_the_ddr2_sdram),                            //                    .mem_clk_n
		.mem_cs_n          (mem_cs_n_from_the_ddr2_sdram),                                    //                    .mem_cs_n
		.mem_cke           (mem_cke_from_the_ddr2_sdram),                                     //                    .mem_cke
		.mem_addr          (mem_addr_from_the_ddr2_sdram),                                    //                    .mem_addr
		.mem_ba            (mem_ba_from_the_ddr2_sdram),                                      //                    .mem_ba
		.mem_ras_n         (mem_ras_n_from_the_ddr2_sdram),                                   //                    .mem_ras_n
		.mem_cas_n         (mem_cas_n_from_the_ddr2_sdram),                                   //                    .mem_cas_n
		.mem_we_n          (mem_we_n_from_the_ddr2_sdram),                                    //                    .mem_we_n
		.mem_dq            (mem_dq_to_and_from_the_ddr2_sdram),                               //                    .mem_dq
		.mem_dqs           (mem_dqs_to_and_from_the_ddr2_sdram),                              //                    .mem_dqs
		.mem_dm            (mem_dm_from_the_ddr2_sdram),                                      //                    .mem_dm
		.pll_ref_clk       (clk),                                                             //              refclk.clk
		.soft_reset_n      (~rst_controller_reset_out_reset),                                 //        soft_reset_n.reset_n
		.global_reset_n    (ddr2_sdram_reset_n),                                              //      global_reset_n.reset_n
		.reset_request_n   (ddr2_sdram_reset_request_n_reset),                                //     reset_request_n.reset_n
		.phy_clk           (ddr2_sdram_phy_clk_out),                                          //              sysclk.clk
		.aux_full_rate_clk (ddr2_sdram_aux_full_rate_clk_out),                                //             auxfull.clk
		.aux_half_rate_clk (ddr2_sdram_aux_half_rate_clk_out)                                 //             auxhalf.clk
	);

	application_selector_ddr2_sdram_1 ddr2_sdram_1 (
		.local_address     (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_address),            //                  s1.address
		.local_write_req   (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_write),              //                    .write
		.local_read_req    (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_read),               //                    .read
		.local_burstbegin  (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_beginbursttransfer), //                    .beginbursttransfer
		.local_ready       (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_waitrequest),        //                    .waitrequest_n
		.local_rdata       (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_readdata),           //                    .readdata
		.local_rdata_valid (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_readdatavalid),      //                    .readdatavalid
		.local_wdata       (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_writedata),          //                    .writedata
		.local_be          (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_byteenable),         //                    .byteenable
		.local_size        (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_burstcount),         //                    .burstcount
		.local_refresh_ack (local_refresh_ack_from_the_ddr2_sdram_1),                           // external_connection.export
		.local_wdata_req   (local_wdata_req_from_the_ddr2_sdram_1),                             //                    .export
		.local_init_done   (local_init_done_from_the_ddr2_sdram_1),                             //                    .export
		.reset_phy_clk_n   (reset_phy_clk_n_from_the_ddr2_sdram_1),                             //                    .export
		.mem_odt           (mem_odt_from_the_ddr2_sdram_1),                                     //              memory.mem_odt
		.mem_clk           (mem_clk_to_and_from_the_ddr2_sdram_1),                              //                    .mem_clk
		.mem_clk_n         (mem_clk_n_to_and_from_the_ddr2_sdram_1),                            //                    .mem_clk_n
		.mem_cs_n          (mem_cs_n_from_the_ddr2_sdram_1),                                    //                    .mem_cs_n
		.mem_cke           (mem_cke_from_the_ddr2_sdram_1),                                     //                    .mem_cke
		.mem_addr          (mem_addr_from_the_ddr2_sdram_1),                                    //                    .mem_addr
		.mem_ba            (mem_ba_from_the_ddr2_sdram_1),                                      //                    .mem_ba
		.mem_ras_n         (mem_ras_n_from_the_ddr2_sdram_1),                                   //                    .mem_ras_n
		.mem_cas_n         (mem_cas_n_from_the_ddr2_sdram_1),                                   //                    .mem_cas_n
		.mem_we_n          (mem_we_n_from_the_ddr2_sdram_1),                                    //                    .mem_we_n
		.mem_dq            (mem_dq_to_and_from_the_ddr2_sdram_1),                               //                    .mem_dq
		.mem_dqs           (mem_dqs_to_and_from_the_ddr2_sdram_1),                              //                    .mem_dqs
		.mem_dm            (mem_dm_from_the_ddr2_sdram_1),                                      //                    .mem_dm
		.pll_ref_clk       (clk_125),                                                           //              refclk.clk
		.soft_reset_n      (~rst_controller_002_reset_out_reset),                               //        soft_reset_n.reset_n
		.global_reset_n    (ddr2_sdram_1_reset_n),                                              //      global_reset_n.reset_n
		.reset_request_n   (ddr2_sdram_1_reset_request_n_reset),                                //     reset_request_n.reset_n
		.phy_clk           (ddr2_sdram_1_phy_clk_out),                                          //              sysclk.clk
		.aux_full_rate_clk (ddr2_sdram_1_aux_full_rate_clk_out),                                //             auxfull.clk
		.aux_half_rate_clk (ddr2_sdram_1_aux_half_rate_clk_out)                                 //             auxhalf.clk
	);

	application_selector_sgdma_tx sgdma_tx (
		.clk                           (pll_c0_out),                                             //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),                    //            reset.reset_n
		.csr_chipselect                (sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_tx_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_tx_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_tx_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_tx_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_tx_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_mapper_receiver5_irq),                               //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                               //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),                          //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),                            //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                                //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                                   //                 .read
		.out_data                      (sgdma_tx_out_data),                                      //              out.data
		.out_valid                     (sgdma_tx_out_valid),                                     //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                                     //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                               //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                             //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                                     //                 .empty
		.out_error                     (sgdma_tx_out_error)                                      //                 .error
	);

	application_selector_sgdma_rx sgdma_rx (
		.clk                           (pll_c0_out),                                             //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),                    //            reset.reset_n
		.csr_chipselect                (sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_rx_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_rx_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_rx_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_rx_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_rx_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_mapper_receiver4_irq),                               //          csr_irq.irq
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),                           //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                               //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                                 //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                             //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable),                            //                 .byteenable
		.in_startofpacket              (tse_mac_receive_startofpacket),                          //               in.startofpacket
		.in_endofpacket                (tse_mac_receive_endofpacket),                            //                 .endofpacket
		.in_empty                      (tse_mac_receive_empty),                                  //                 .empty
		.in_data                       (tse_mac_receive_data),                                   //                 .data
		.in_valid                      (tse_mac_receive_valid),                                  //                 .valid
		.in_ready                      (tse_mac_receive_ready),                                  //                 .ready
		.in_error                      (tse_mac_receive_error)                                   //                 .error
	);

	application_selector_lcd_sgdma lcd_sgdma (
		.clk                           (ddr2_sdram_phy_clk_out),                                  //              clk.clk
		.system_reset_n                (~rst_controller_003_reset_out_reset),                     //            reset.reset_n
		.csr_chipselect                (lcd_sgdma_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (lcd_sgdma_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (lcd_sgdma_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (lcd_sgdma_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (lcd_sgdma_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (lcd_sgdma_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (lcd_sgdma_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (lcd_sgdma_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (lcd_sgdma_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (lcd_sgdma_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (lcd_sgdma_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (lcd_sgdma_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (lcd_sgdma_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (lcd_sgdma_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (lcd_sgdma_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_synchronizer_003_receiver_irq),                       //          csr_irq.irq
		.m_read_readdata               (lcd_sgdma_m_read_readdata),                               //           m_read.readdata
		.m_read_readdatavalid          (lcd_sgdma_m_read_readdatavalid),                          //                 .readdatavalid
		.m_read_waitrequest            (lcd_sgdma_m_read_waitrequest),                            //                 .waitrequest
		.m_read_address                (lcd_sgdma_m_read_address),                                //                 .address
		.m_read_read                   (lcd_sgdma_m_read_read),                                   //                 .read
		.out_data                      (lcd_sgdma_out_data),                                      //              out.data
		.out_valid                     (lcd_sgdma_out_valid),                                     //                 .valid
		.out_ready                     (lcd_sgdma_out_ready),                                     //                 .ready
		.out_endofpacket               (lcd_sgdma_out_endofpacket),                               //                 .endofpacket
		.out_startofpacket             (lcd_sgdma_out_startofpacket),                             //                 .startofpacket
		.out_empty                     (lcd_sgdma_out_empty)                                      //                 .empty
	);

	application_selector_tse_mac tse_mac (
		.ff_tx_data  (sgdma_tx_out_data),                                               //                      transmit.data
		.ff_tx_eop   (sgdma_tx_out_endofpacket),                                        //                              .endofpacket
		.ff_tx_err   (sgdma_tx_out_error),                                              //                              .error
		.ff_tx_mod   (sgdma_tx_out_empty),                                              //                              .empty
		.ff_tx_rdy   (sgdma_tx_out_ready),                                              //                              .ready
		.ff_tx_sop   (sgdma_tx_out_startofpacket),                                      //                              .startofpacket
		.ff_tx_wren  (sgdma_tx_out_valid),                                              //                              .valid
		.ff_tx_clk   (pll_c0_out),                                                      //      receive_clock_connection.clk
		.ff_rx_data  (tse_mac_receive_data),                                            //                       receive.data
		.ff_rx_dval  (tse_mac_receive_valid),                                           //                              .valid
		.ff_rx_eop   (tse_mac_receive_endofpacket),                                     //                              .endofpacket
		.ff_rx_mod   (tse_mac_receive_empty),                                           //                              .empty
		.ff_rx_rdy   (tse_mac_receive_ready),                                           //                              .ready
		.ff_rx_sop   (tse_mac_receive_startofpacket),                                   //                              .startofpacket
		.rx_err      (tse_mac_receive_error),                                           //                              .error
		.ff_rx_clk   (pll_c0_out),                                                      //     transmit_clock_connection.clk
		.address     (tse_mac_control_port_translator_avalon_anti_slave_0_address),     //                  control_port.address
		.readdata    (tse_mac_control_port_translator_avalon_anti_slave_0_readdata),    //                              .readdata
		.read        (tse_mac_control_port_translator_avalon_anti_slave_0_read),        //                              .read
		.writedata   (tse_mac_control_port_translator_avalon_anti_slave_0_writedata),   //                              .writedata
		.write       (tse_mac_control_port_translator_avalon_anti_slave_0_write),       //                              .write
		.waitrequest (tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest), //                              .waitrequest
		.clk         (pll_c0_out),                                                      // control_port_clock_connection.clk
		.reset       (rst_controller_001_reset_out_reset),                              //              reset_connection.reset
		.gm_rx_d     (gm_rx_d_to_the_tse_mac),                                          //            conduit_connection.export
		.gm_rx_dv    (gm_rx_dv_to_the_tse_mac),                                         //                              .export
		.gm_rx_err   (gm_rx_err_to_the_tse_mac),                                        //                              .export
		.gm_tx_d     (gm_tx_d_from_the_tse_mac),                                        //                              .export
		.gm_tx_en    (gm_tx_en_from_the_tse_mac),                                       //                              .export
		.gm_tx_err   (gm_tx_err_from_the_tse_mac),                                      //                              .export
		.m_rx_d      (m_rx_d_to_the_tse_mac),                                           //                              .export
		.m_rx_en     (m_rx_en_to_the_tse_mac),                                          //                              .export
		.m_rx_err    (m_rx_err_to_the_tse_mac),                                         //                              .export
		.m_tx_d      (m_tx_d_from_the_tse_mac),                                         //                              .export
		.m_tx_en     (m_tx_en_from_the_tse_mac),                                        //                              .export
		.m_tx_err    (m_tx_err_from_the_tse_mac),                                       //                              .export
		.m_rx_col    (m_rx_col_to_the_tse_mac),                                         //                              .export
		.m_rx_crs    (m_rx_crs_to_the_tse_mac),                                         //                              .export
		.tx_clk      (tx_clk_to_the_tse_mac),                                           //                              .export
		.rx_clk      (rx_clk_to_the_tse_mac),                                           //                              .export
		.set_10      (set_10_to_the_tse_mac),                                           //                              .export
		.set_1000    (set_1000_to_the_tse_mac),                                         //                              .export
		.ena_10      (ena_10_from_the_tse_mac),                                         //                              .export
		.eth_mode    (eth_mode_from_the_tse_mac),                                       //                              .export
		.mdio_out    (mdio_out_from_the_tse_mac),                                       //                              .export
		.mdio_oen    (mdio_oen_from_the_tse_mac),                                       //                              .export
		.mdio_in     (mdio_in_to_the_tse_mac),                                          //                              .export
		.mdc         (mdc_from_the_tse_mac)                                             //                              .export
	);

	application_selector_sys_clk_timer sys_clk_timer (
		.clk        (pll_c2_out),                                                 //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                        // reset.reset_n
		.address    (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~sys_clk_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_004_receiver_irq)                           //   irq.irq
	);

	application_selector_high_res_timer high_res_timer (
		.clk        (pll_c2_out),                                                  //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                         // reset.reset_n
		.address    (high_res_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_res_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_res_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_res_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_res_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)                            //   irq.irq
	);

	application_selector_performance_counter performance_counter (
		.clk           (pll_c2_out),                                                                     //           clk.clk
		.reset_n       (~rst_controller_004_reset_out_reset),                                            //         reset.reset_n
		.address       (performance_counter_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.readdata      (performance_counter_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (performance_counter_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (performance_counter_control_slave_translator_avalon_anti_slave_0_writedata)      //              .writedata
	);

	application_selector_jtag_uart jtag_uart (
		.clk            (pll_c2_out),                                                             //               clk.clk
		.rst_n          (~rst_controller_004_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.dataavailable  (),                                                                       //                  .dataavailable
		.readyfordata   (),                                                                       //                  .readyfordata
		.av_irq         (irq_synchronizer_002_receiver_irq)                                       //               irq.irq
	);

	application_selector_uart1 uart1 (
		.clk           (pll_c2_out),                                            //                 clk.clk
		.reset_n       (~rst_controller_004_reset_out_reset),                   //               reset.reset_n
		.address       (uart1_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart1_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart1_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart1_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart1_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart1_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart1_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                      //                    .dataavailable
		.readyfordata  (),                                                      //                    .readyfordata
		.rxd           (rxd_to_the_uart1),                                      // external_connection.export
		.txd           (txd_from_the_uart1),                                    //                    .export
		.irq           (irq_synchronizer_007_receiver_irq)                      //                 irq.irq
	);

	application_selector_button_pio button_pio (
		.clk        (pll_c2_out),                                              //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                     //               reset.reset_n
		.address    (button_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~button_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (button_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (button_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (button_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (in_port_to_the_button_pio),                               // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)                            //                 irq.irq
	);

	application_selector_led_pio led_pio (
		.clk        (pll_c2_out),                                           //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                  //               reset.reset_n
		.address    (led_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_led_pio)                             // external_connection.export
	);

	application_selector_pio_id_eeprom_scl pio_id_eeprom_scl (
		.clk        (pll_c2_out),                                                     //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                            //               reset.reset_n
		.address    (pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_pio_id_eeprom_scl)                             // external_connection.export
	);

	application_selector_pio_id_eeprom_scl lcd_i2c_scl (
		.clk        (pll_c2_out),                                               //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                      //               reset.reset_n
		.address    (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_i2c_scl_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_lcd_i2c_scl)                             // external_connection.export
	);

	application_selector_pio_id_eeprom_scl lcd_i2c_en (
		.clk        (pll_c2_out),                                              //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                     //               reset.reset_n
		.address    (lcd_i2c_en_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_i2c_en_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_i2c_en_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_i2c_en_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_i2c_en_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_lcd_i2c_en)                             // external_connection.export
	);

	application_selector_pio_id_eeprom_dat pio_id_eeprom_dat (
		.clk        (pll_c2_out),                                                     //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                            //               reset.reset_n
		.address    (pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (bidir_port_to_and_from_the_pio_id_eeprom_dat)                    // external_connection.export
	);

	application_selector_pio_id_eeprom_dat lcd_i2c_sdat (
		.clk        (pll_c2_out),                                                //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                       //               reset.reset_n
		.address    (lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (bidir_port_to_and_from_the_lcd_i2c_sdat)                    // external_connection.export
	);

	application_selector_touch_panel_pen_irq_n touch_panel_pen_irq_n (
		.clk        (pll_c2_out),                                                         //                 clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),                                //               reset.reset_n
		.address    (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (in_port_to_the_touch_panel_pen_irq_n),                               // external_connection.export
		.irq        (irq_synchronizer_005_receiver_irq)                                   //                 irq.irq
	);

	application_selector_touch_panel_spi touch_panel_spi (
		.clk           (pll_c2_out),                                                                 //              clk.clk
		.reset_n       (~rst_controller_004_reset_out_reset),                                        //            reset.reset_n
		.data_from_cpu (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_writedata),  // spi_control_port.writedata
		.data_to_cpu   (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.mem_addr      (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_address),    //                 .address
		.read_n        (~touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_read),      //                 .read_n
		.spi_select    (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_chipselect), //                 .chipselect
		.write_n       (~touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_write),     //                 .write_n
		.dataavailable (),                                                                           //                 .dataavailable
		.endofpacket   (),                                                                           //                 .endofpacket
		.readyfordata  (),                                                                           //                 .readyfordata
		.irq           (irq_synchronizer_006_receiver_irq),                                          //              irq.irq
		.MISO          (MISO_to_the_touch_panel_spi),                                                //         external.export
		.MOSI          (MOSI_from_the_touch_panel_spi),                                              //                 .export
		.SCLK          (SCLK_from_the_touch_panel_spi),                                              //                 .export
		.SS_n          (SS_n_from_the_touch_panel_spi)                                               //                 .export
	);

	application_selector_lcd_ta_sgdma_to_fifo lcd_ta_sgdma_to_fifo (
		.clk               (ddr2_sdram_phy_clk_out),                 //   clk.clk
		.reset_n           (~rst_controller_003_reset_out_reset),    // reset.reset_n
		.in_ready          (lcd_sgdma_out_ready),                    //    in.ready
		.in_valid          (lcd_sgdma_out_valid),                    //      .valid
		.in_data           (lcd_sgdma_out_data),                     //      .data
		.in_startofpacket  (lcd_sgdma_out_startofpacket),            //      .startofpacket
		.in_endofpacket    (lcd_sgdma_out_endofpacket),              //      .endofpacket
		.in_empty          (lcd_sgdma_out_empty),                    //      .empty
		.out_ready         (lcd_ta_sgdma_to_fifo_out_ready),         //   out.ready
		.out_valid         (lcd_ta_sgdma_to_fifo_out_valid),         //      .valid
		.out_data          (lcd_ta_sgdma_to_fifo_out_data),          //      .data
		.out_startofpacket (lcd_ta_sgdma_to_fifo_out_startofpacket), //      .startofpacket
		.out_endofpacket   (lcd_ta_sgdma_to_fifo_out_endofpacket),   //      .endofpacket
		.out_empty         (lcd_ta_sgdma_to_fifo_out_empty)          //      .empty
	);

	application_selector_lcd_pixel_fifo lcd_pixel_fifo (
		.wrclock                       (ddr2_sdram_phy_clk_out),                 //    clk_in.clk
		.wrreset_n                     (~rst_controller_003_reset_out_reset),    //  reset_in.reset_n
		.avalonst_sink_valid           (lcd_ta_sgdma_to_fifo_out_valid),         //        in.valid
		.avalonst_sink_data            (lcd_ta_sgdma_to_fifo_out_data),          //          .data
		.avalonst_sink_startofpacket   (lcd_ta_sgdma_to_fifo_out_startofpacket), //          .startofpacket
		.avalonst_sink_endofpacket     (lcd_ta_sgdma_to_fifo_out_endofpacket),   //          .endofpacket
		.avalonst_sink_empty           (lcd_ta_sgdma_to_fifo_out_empty),         //          .empty
		.avalonst_sink_ready           (lcd_ta_sgdma_to_fifo_out_ready),         //          .ready
		.rdclock                       (pll_c0_out),                             //   clk_out.clk
		.rdreset_n                     (~rst_controller_001_reset_out_reset),    // reset_out.reset_n
		.avalonst_source_valid         (lcd_pixel_fifo_out_valid),               //       out.valid
		.avalonst_source_data          (lcd_pixel_fifo_out_data),                //          .data
		.avalonst_source_startofpacket (lcd_pixel_fifo_out_startofpacket),       //          .startofpacket
		.avalonst_source_endofpacket   (lcd_pixel_fifo_out_endofpacket),         //          .endofpacket
		.avalonst_source_empty         (lcd_pixel_fifo_out_empty),               //          .empty
		.avalonst_source_ready         (lcd_pixel_fifo_out_ready)                //          .ready
	);

	application_selector_lcd_ta_fifo_to_dfa lcd_ta_fifo_to_dfa (
		.clk               (pll_c0_out),                           //   clk.clk
		.reset_n           (~rst_controller_001_reset_out_reset),  // reset.reset_n
		.in_ready          (lcd_pixel_fifo_out_ready),             //    in.ready
		.in_valid          (lcd_pixel_fifo_out_valid),             //      .valid
		.in_data           (lcd_pixel_fifo_out_data),              //      .data
		.in_startofpacket  (lcd_pixel_fifo_out_startofpacket),     //      .startofpacket
		.in_endofpacket    (lcd_pixel_fifo_out_endofpacket),       //      .endofpacket
		.in_empty          (lcd_pixel_fifo_out_empty),             //      .empty
		.out_ready         (lcd_ta_fifo_to_dfa_out_ready),         //   out.ready
		.out_valid         (lcd_ta_fifo_to_dfa_out_valid),         //      .valid
		.out_data          (lcd_ta_fifo_to_dfa_out_data),          //      .data
		.out_startofpacket (lcd_ta_fifo_to_dfa_out_startofpacket), //      .startofpacket
		.out_endofpacket   (lcd_ta_fifo_to_dfa_out_endofpacket),   //      .endofpacket
		.out_empty         (lcd_ta_fifo_to_dfa_out_empty)          //      .empty
	);

	application_selector_lcd_64_to_32_bits_dfa lcd_64_to_32_bits_dfa (
		.clk               (pll_c0_out),                              //   clk.clk
		.reset_n           (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.in_ready          (lcd_ta_fifo_to_dfa_out_ready),            //    in.ready
		.in_valid          (lcd_ta_fifo_to_dfa_out_valid),            //      .valid
		.in_data           (lcd_ta_fifo_to_dfa_out_data),             //      .data
		.in_startofpacket  (lcd_ta_fifo_to_dfa_out_startofpacket),    //      .startofpacket
		.in_endofpacket    (lcd_ta_fifo_to_dfa_out_endofpacket),      //      .endofpacket
		.in_empty          (lcd_ta_fifo_to_dfa_out_empty),            //      .empty
		.out_ready         (lcd_64_to_32_bits_dfa_out_ready),         //   out.ready
		.out_valid         (lcd_64_to_32_bits_dfa_out_valid),         //      .valid
		.out_data          (lcd_64_to_32_bits_dfa_out_data),          //      .data
		.out_startofpacket (lcd_64_to_32_bits_dfa_out_startofpacket), //      .startofpacket
		.out_endofpacket   (lcd_64_to_32_bits_dfa_out_endofpacket),   //      .endofpacket
		.out_empty         (lcd_64_to_32_bits_dfa_out_empty)          //      .empty
	);

	altera_avalon_pixel_converter #(
		.SOURCE_SYMBOLS_PER_BEAT (3)
	) lcd_pixel_converter (
		.clk       (pll_c0_out),                              //       clk.clk
		.reset_n   (~rst_controller_001_reset_out_reset),     // clk_reset.reset_n
		.ready_out (lcd_64_to_32_bits_dfa_out_ready),         //        in.ready
		.valid_in  (lcd_64_to_32_bits_dfa_out_valid),         //          .valid
		.data_in   (lcd_64_to_32_bits_dfa_out_data),          //          .data
		.eop_in    (lcd_64_to_32_bits_dfa_out_endofpacket),   //          .endofpacket
		.sop_in    (lcd_64_to_32_bits_dfa_out_startofpacket), //          .startofpacket
		.empty_in  (lcd_64_to_32_bits_dfa_out_empty),         //          .empty
		.ready_in  (lcd_pixel_converter_out_ready),           //       out.ready
		.valid_out (lcd_pixel_converter_out_valid),           //          .valid
		.data_out  (lcd_pixel_converter_out_data),            //          .data
		.eop_out   (lcd_pixel_converter_out_endofpacket),     //          .endofpacket
		.sop_out   (lcd_pixel_converter_out_startofpacket),   //          .startofpacket
		.empty_out (lcd_pixel_converter_out_empty)            //          .empty
	);

	application_selector_lcd_32_to_8_bits_dfa lcd_32_to_8_bits_dfa (
		.clk               (pll_c0_out),                             //   clk.clk
		.reset_n           (~rst_controller_001_reset_out_reset),    // reset.reset_n
		.in_ready          (lcd_pixel_converter_out_ready),          //    in.ready
		.in_valid          (lcd_pixel_converter_out_valid),          //      .valid
		.in_data           (lcd_pixel_converter_out_data),           //      .data
		.in_startofpacket  (lcd_pixel_converter_out_startofpacket),  //      .startofpacket
		.in_endofpacket    (lcd_pixel_converter_out_endofpacket),    //      .endofpacket
		.in_empty          (lcd_pixel_converter_out_empty),          //      .empty
		.out_ready         (lcd_32_to_8_bits_dfa_out_ready),         //   out.ready
		.out_valid         (lcd_32_to_8_bits_dfa_out_valid),         //      .valid
		.out_data          (lcd_32_to_8_bits_dfa_out_data),          //      .data
		.out_startofpacket (lcd_32_to_8_bits_dfa_out_startofpacket), //      .startofpacket
		.out_endofpacket   (lcd_32_to_8_bits_dfa_out_endofpacket),   //      .endofpacket
		.out_empty         (lcd_32_to_8_bits_dfa_out_empty)          //      .empty
	);

	altera_avalon_video_sync_generator #(
		.DATA_STREAM_BIT_WIDTH (8),
		.BEATS_PER_PIXEL       (3),
		.NUM_COLUMNS           (800),
		.NUM_ROWS              (480),
		.H_BLANK_PIXELS        (216),
		.H_FRONT_PORCH_PIXELS  (40),
		.H_SYNC_PULSE_PIXELS   (1),
		.H_SYNC_PULSE_POLARITY (0),
		.V_BLANK_LINES         (35),
		.V_FRONT_PORCH_LINES   (10),
		.V_SYNC_PULSE_LINES    (1),
		.V_SYNC_PULSE_POLARITY (0),
		.TOTAL_HSCAN_PIXELS    (1056),
		.TOTAL_VSCAN_LINES     (525)
	) lcd_sync_generator (
		.clk     (pll_c0_out),                             //       clk.clk
		.reset_n (~rst_controller_001_reset_out_reset),    // clk_reset.reset_n
		.ready   (lcd_32_to_8_bits_dfa_out_ready),         //        in.ready
		.valid   (lcd_32_to_8_bits_dfa_out_valid),         //          .valid
		.data    (lcd_32_to_8_bits_dfa_out_data),          //          .data
		.eop     (lcd_32_to_8_bits_dfa_out_endofpacket),   //          .endofpacket
		.sop     (lcd_32_to_8_bits_dfa_out_startofpacket), //          .startofpacket
		.empty   (lcd_32_to_8_bits_dfa_out_empty),         //          .empty
		.RGB_OUT (RGB_OUT_from_the_lcd_sync_generator),    //      sync.export
		.HD      (HD_from_the_lcd_sync_generator),         //          .export
		.VD      (VD_from_the_lcd_sync_generator),         //          .export
		.DEN     (DEN_from_the_lcd_sync_generator)         //          .export
	);

	sls_sdhc_top #(
		.tx_buffer_depth (2048),
		.tx_buffer_add   (11),
		.rx_buffer_depth (2048),
		.rx_buffer_add   (11)
	) sls_sdhc (
		.clk                  (clk),                                                         //            clock.clk
		.reset_n              (~rst_controller_reset_out_reset),                             //      clock_reset.reset_n
		.AvS_address          (sls_sdhc_control_translator_avalon_anti_slave_0_address),     //          control.address
		.AvS_chipselect       (sls_sdhc_control_translator_avalon_anti_slave_0_chipselect),  //                 .chipselect
		.AvS_write_n          (~sls_sdhc_control_translator_avalon_anti_slave_0_write),      //                 .write_n
		.AvS_read_n           (~sls_sdhc_control_translator_avalon_anti_slave_0_read),       //                 .read_n
		.AvS_writedata        (sls_sdhc_control_translator_avalon_anti_slave_0_writedata),   //                 .writedata
		.AvS_readdata         (sls_sdhc_control_translator_avalon_anti_slave_0_readdata),    //                 .readdata
		.AvS_waitrequest      (sls_sdhc_control_translator_avalon_anti_slave_0_waitrequest), //                 .waitrequest
		.AvM_wr_address       (sls_sdhc_write_master_address),                               //     write_master.address
		.AvM_wr_writedata     (sls_sdhc_write_master_writedata),                             //                 .writedata
		.AvM_wr_write_n       (sls_sdhc_write_master_write),                                 //                 .write_n
		.AvM_wr_chipselect    (sls_sdhc_write_master_chipselect),                            //                 .chipselect
		.AvM_wr_waitrequest   (sls_sdhc_write_master_waitrequest),                           //                 .waitrequest
		.AvM_wr_byteenable    (sls_sdhc_write_master_byteenable),                            //                 .byteenable
		.AvM_rd_readdata      (sls_sdhc_read_master_readdata),                               //      read_master.readdata
		.AvM_rd_read_n        (sls_sdhc_read_master_read),                                   //                 .read_n
		.AvM_rd_address       (sls_sdhc_read_master_address),                                //                 .address
		.AvM_rd_waitrequest   (sls_sdhc_read_master_waitrequest),                            //                 .waitrequest
		.AvM_rd_readdatavalid (sls_sdhc_read_master_readdatavalid),                          //                 .readdatavalid
		.AvM_rd_byteenable    (sls_sdhc_read_master_byteenable),                             //                 .byteenable
		.AvS_irq              (irq_synchronizer_008_receiver_irq),                           // interrupt_sender.irq
		.SD_CLK               (SD_CLK_from_the_sls_sdhc),                                    //      conduit_end.export
		.SD_CMD               (SD_CMD_to_and_from_the_sls_sdhc),                             //                 .export
		.SD_DAT0              (SD_DAT0_to_and_from_the_sls_sdhc),                            //                 .export
		.SD_DAT1              (SD_DAT1_to_and_from_the_sls_sdhc),                            //                 .export
		.SD_DAT2              (SD_DAT2_to_and_from_the_sls_sdhc),                            //                 .export
		.SD_DAT3              (SD_DAT3_to_and_from_the_sls_sdhc),                            //                 .export
		.SD_In                (SD_In_to_the_sls_sdhc),                                       //                 .export
		.SD_Wp                (SD_Wp_to_the_sls_sdhc),                                       //                 .export
		.SD_Busy              (SD_Busy_from_the_sls_sdhc)                                    //                 .export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (27),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipeline_bridge_before_tristate_bridge (
		.clk              (pll_c0_out),                                                                             //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                     // reset.reset
		.s0_waitrequest   (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.s0_readdatavalid (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.s0_writedata     (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.s0_address       (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_address),       //      .address
		.s0_write         (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_write),         //      .write
		.s0_read          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_read),          //      .read
		.s0_byteenable    (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.s0_debugaccess   (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pipeline_bridge_before_tristate_bridge_m0_waitrequest),                                  //    m0.waitrequest
		.m0_readdata      (pipeline_bridge_before_tristate_bridge_m0_readdata),                                     //      .readdata
		.m0_readdatavalid (pipeline_bridge_before_tristate_bridge_m0_readdatavalid),                                //      .readdatavalid
		.m0_burstcount    (pipeline_bridge_before_tristate_bridge_m0_burstcount),                                   //      .burstcount
		.m0_writedata     (pipeline_bridge_before_tristate_bridge_m0_writedata),                                    //      .writedata
		.m0_address       (pipeline_bridge_before_tristate_bridge_m0_address),                                      //      .address
		.m0_write         (pipeline_bridge_before_tristate_bridge_m0_write),                                        //      .write
		.m0_read          (pipeline_bridge_before_tristate_bridge_m0_read),                                         //      .read
		.m0_byteenable    (pipeline_bridge_before_tristate_bridge_m0_byteenable),                                   //      .byteenable
		.m0_debugaccess   (pipeline_bridge_before_tristate_bridge_m0_debugaccess)                                   //      .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (64),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (26),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) sdhc_ddr_clock_bridge (
		.m0_clk           (ddr2_sdram_phy_clk_out),                                                //   m0_clk.clk
		.m0_reset         (rst_controller_003_reset_out_reset),                                    // m0_reset.reset
		.s0_clk           (pll_c0_out),                                                            //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                                    // s0_reset.reset
		.s0_waitrequest   (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (sdhc_ddr_clock_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (sdhc_ddr_clock_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (sdhc_ddr_clock_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (sdhc_ddr_clock_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (sdhc_ddr_clock_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (sdhc_ddr_clock_bridge_m0_address),                                      //         .address
		.m0_write         (sdhc_ddr_clock_bridge_m0_write),                                        //         .write
		.m0_read          (sdhc_ddr_clock_bridge_m0_read),                                         //         .read
		.m0_byteenable    (sdhc_ddr_clock_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (sdhc_ddr_clock_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (27),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) cpu_ddr_clock_bridge (
		.m0_clk           (ddr2_sdram_phy_clk_out),                                               //   m0_clk.clk
		.m0_reset         (rst_controller_003_reset_out_reset),                                   // m0_reset.reset
		.s0_clk           (pll_c0_out),                                                           //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                                   // s0_reset.reset
		.s0_waitrequest   (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (cpu_ddr_clock_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (cpu_ddr_clock_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (cpu_ddr_clock_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (cpu_ddr_clock_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (cpu_ddr_clock_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (cpu_ddr_clock_bridge_m0_address),                                      //         .address
		.m0_write         (cpu_ddr_clock_bridge_m0_write),                                        //         .write
		.m0_read          (cpu_ddr_clock_bridge_m0_read),                                         //         .read
		.m0_byteenable    (cpu_ddr_clock_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (cpu_ddr_clock_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (26),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) cpu_ddr_1_clock_bridge (
		.m0_clk           (ddr2_sdram_1_phy_clk_out),                                               //   m0_clk.clk
		.m0_reset         (rst_controller_005_reset_out_reset),                                     // m0_reset.reset
		.s0_clk           (pll_c0_out),                                                             //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                                     // s0_reset.reset
		.s0_waitrequest   (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (cpu_ddr_1_clock_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (cpu_ddr_1_clock_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (cpu_ddr_1_clock_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (cpu_ddr_1_clock_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (cpu_ddr_1_clock_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (cpu_ddr_1_clock_bridge_m0_address),                                      //         .address
		.m0_write         (cpu_ddr_1_clock_bridge_m0_write),                                        //         .write
		.m0_read          (cpu_ddr_1_clock_bridge_m0_read),                                         //         .read
		.m0_byteenable    (cpu_ddr_1_clock_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (cpu_ddr_1_clock_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) slow_peripheral_bridge (
		.m0_clk           (pll_c2_out),                                                             //   m0_clk.clk
		.m0_reset         (rst_controller_004_reset_out_reset),                                     // m0_reset.reset
		.s0_clk           (pll_c0_out),                                                             //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                                     // s0_reset.reset
		.s0_waitrequest   (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (slow_peripheral_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (slow_peripheral_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (slow_peripheral_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (slow_peripheral_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (slow_peripheral_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (slow_peripheral_bridge_m0_address),                                      //         .address
		.m0_write         (slow_peripheral_bridge_m0_write),                                        //         .write
		.m0_read          (slow_peripheral_bridge_m0_read),                                         //         .read
		.m0_byteenable    (slow_peripheral_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (slow_peripheral_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (26),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) tse_ddr_clock_bridge (
		.m0_clk           (ddr2_sdram_phy_clk_out),                                               //   m0_clk.clk
		.m0_reset         (rst_controller_003_reset_out_reset),                                   // m0_reset.reset
		.s0_clk           (pll_c0_out),                                                           //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                                   // s0_reset.reset
		.s0_waitrequest   (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (tse_ddr_clock_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (tse_ddr_clock_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (tse_ddr_clock_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (tse_ddr_clock_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (tse_ddr_clock_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (tse_ddr_clock_bridge_m0_address),                                      //         .address
		.m0_write         (tse_ddr_clock_bridge_m0_write),                                        //         .write
		.m0_read          (tse_ddr_clock_bridge_m0_read),                                         //         .read
		.m0_byteenable    (tse_ddr_clock_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (tse_ddr_clock_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	application_selector_cpu cpu (
		.clk                                   (pll_c0_out),                                                         //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                                //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	application_selector_sysid sysid (
		.clock    (pll_c2_out),                                                  //           clk.clk
		.reset_n  (~rst_controller_004_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	application_selector_flash_tristate_bridge_bridge_0 flash_tristate_bridge_bridge_0 (
		.clk                                  (pll_c0_out),                                                              //   clk.clk
		.reset                                (rst_controller_001_reset_out_reset),                                      // reset.reset
		.request                              (flash_tristate_bridge_pinsharer_0_tcm_request),                           //   tcs.request
		.grant                                (flash_tristate_bridge_pinsharer_0_tcm_grant),                             //      .grant
		.tcs_read_n_to_the_ext_flash          (flash_tristate_bridge_pinsharer_0_tcm_read_n_to_the_ext_flash_out),       //      .read_n_to_the_ext_flash_out
		.tcs_select_n_to_the_ext_flash        (flash_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out),     //      .select_n_to_the_ext_flash_out
		.tcs_oe_n_to_the_max2                 (flash_tristate_bridge_pinsharer_0_tcm_oe_n_to_the_max2_out),              //      .oe_n_to_the_max2_out
		.tcs_cs_n_to_the_max2                 (flash_tristate_bridge_pinsharer_0_tcm_cs_n_to_the_max2_out),              //      .cs_n_to_the_max2_out
		.tcs_flash_tristate_bridge_data       (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_out),    //      .flash_tristate_bridge_data_out
		.tcs_flash_tristate_bridge_data_outen (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_outen),  //      .flash_tristate_bridge_data_outen
		.tcs_flash_tristate_bridge_data_in    (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_in),     //      .flash_tristate_bridge_data_in
		.tcs_write_n_to_the_ext_flash         (flash_tristate_bridge_pinsharer_0_tcm_write_n_to_the_ext_flash_out),      //      .write_n_to_the_ext_flash_out
		.tcs_flash_tristate_bridge_address    (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_address_out), //      .flash_tristate_bridge_address_out
		.tcs_we_n_to_the_max2                 (flash_tristate_bridge_pinsharer_0_tcm_we_n_to_the_max2_out),              //      .we_n_to_the_max2_out
		.read_n_to_the_ext_flash              (read_n_to_the_ext_flash),                                                 //   out.read_n_to_the_ext_flash
		.select_n_to_the_ext_flash            (select_n_to_the_ext_flash),                                               //      .select_n_to_the_ext_flash
		.oe_n_to_the_max2                     (oe_n_to_the_max2),                                                        //      .oe_n_to_the_max2
		.cs_n_to_the_max2                     (cs_n_to_the_max2),                                                        //      .cs_n_to_the_max2
		.flash_tristate_bridge_data           (flash_tristate_bridge_data),                                              //      .flash_tristate_bridge_data
		.write_n_to_the_ext_flash             (write_n_to_the_ext_flash),                                                //      .write_n_to_the_ext_flash
		.flash_tristate_bridge_address        (flash_tristate_bridge_address),                                           //      .flash_tristate_bridge_address
		.we_n_to_the_max2                     (we_n_to_the_max2)                                                         //      .we_n_to_the_max2
	);

	application_selector_flash_tristate_bridge_pinSharer_0 flash_tristate_bridge_pinsharer_0 (
		.clk_clk                          (pll_c0_out),                                                              //   clk.clk
		.reset_reset                      (rst_controller_001_reset_out_reset),                                      // reset.reset
		.request                          (flash_tristate_bridge_pinsharer_0_tcm_request),                           //   tcm.request
		.grant                            (flash_tristate_bridge_pinsharer_0_tcm_grant),                             //      .grant
		.oe_n_to_the_max2                 (flash_tristate_bridge_pinsharer_0_tcm_oe_n_to_the_max2_out),              //      .oe_n_to_the_max2_out
		.we_n_to_the_max2                 (flash_tristate_bridge_pinsharer_0_tcm_we_n_to_the_max2_out),              //      .we_n_to_the_max2_out
		.cs_n_to_the_max2                 (flash_tristate_bridge_pinsharer_0_tcm_cs_n_to_the_max2_out),              //      .cs_n_to_the_max2_out
		.flash_tristate_bridge_address    (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_address_out), //      .flash_tristate_bridge_address_out
		.read_n_to_the_ext_flash          (flash_tristate_bridge_pinsharer_0_tcm_read_n_to_the_ext_flash_out),       //      .read_n_to_the_ext_flash_out
		.write_n_to_the_ext_flash         (flash_tristate_bridge_pinsharer_0_tcm_write_n_to_the_ext_flash_out),      //      .write_n_to_the_ext_flash_out
		.flash_tristate_bridge_data       (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_out),    //      .flash_tristate_bridge_data_out
		.flash_tristate_bridge_data_in    (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_in),     //      .flash_tristate_bridge_data_in
		.flash_tristate_bridge_data_outen (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_outen),  //      .flash_tristate_bridge_data_outen
		.select_n_to_the_ext_flash        (flash_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out),     //      .select_n_to_the_ext_flash_out
		.tcs0_request                     (ext_flash_tcm_request),                                                   //  tcs0.request
		.tcs0_grant                       (ext_flash_tcm_grant),                                                     //      .grant
		.tcs0_address_out                 (ext_flash_tcm_address_out),                                               //      .address_out
		.tcs0_read_n_out                  (ext_flash_tcm_read_n_out),                                                //      .read_n_out
		.tcs0_write_n_out                 (ext_flash_tcm_write_n_out),                                               //      .write_n_out
		.tcs0_data_out                    (ext_flash_tcm_data_out),                                                  //      .data_out
		.tcs0_data_in                     (ext_flash_tcm_data_in),                                                   //      .data_in
		.tcs0_data_outen                  (ext_flash_tcm_data_outen),                                                //      .data_outen
		.tcs0_chipselect_n_out            (ext_flash_tcm_chipselect_n_out),                                          //      .chipselect_n_out
		.tcs1_request                     (max2_tcm_request),                                                        //  tcs1.request
		.tcs1_grant                       (max2_tcm_grant),                                                          //      .grant
		.tcs1_address_out                 (max2_tcm_address_out),                                                    //      .address_out
		.tcs1_read_n_out                  (max2_tcm_read_n_out),                                                     //      .read_n_out
		.tcs1_write_n_out                 (max2_tcm_write_n_out),                                                    //      .write_n_out
		.tcs1_data_out                    (max2_tcm_data_out),                                                       //      .data_out
		.tcs1_data_in                     (max2_tcm_data_in),                                                        //      .data_in
		.tcs1_data_outen                  (max2_tcm_data_outen),                                                     //      .data_outen
		.tcs1_chipselect_n_out            (max2_tcm_chipselect_n_out)                                                //      .chipselect_n_out
	);

	application_selector_ext_flash #(
		.TCM_ADDRESS_W                  (26),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (40),
		.TCM_WRITE_WAIT                 (40),
		.TCM_SETUP_WAIT                 (80),
		.TCM_DATA_HOLD                  (20),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) ext_flash (
		.clk_clk              (pll_c0_out),                                                 //   clk.clk
		.reset_reset          (rst_controller_001_reset_out_reset),                         // reset.reset
		.uas_address          (ext_flash_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (ext_flash_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (ext_flash_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (ext_flash_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (ext_flash_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (ext_flash_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (ext_flash_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (ext_flash_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (ext_flash_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (ext_flash_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (ext_flash_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (ext_flash_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (ext_flash_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (ext_flash_tcm_request),                                      //      .request
		.tcm_grant            (ext_flash_tcm_grant),                                        //      .grant
		.tcm_address_out      (ext_flash_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (ext_flash_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (ext_flash_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (ext_flash_tcm_data_in)                                       //      .data_in
	);

	application_selector_max2 #(
		.TCM_ADDRESS_W                  (5),
		.TCM_DATA_W                     (32),
		.TCM_BYTEENABLE_W               (4),
		.TCM_READ_WAIT                  (100),
		.TCM_WRITE_WAIT                 (100),
		.TCM_SETUP_WAIT                 (0),
		.TCM_DATA_HOLD                  (0),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (4),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) max2 (
		.clk_clk              (pll_c0_out),                                            //   clk.clk
		.reset_reset          (rst_controller_001_reset_out_reset),                    // reset.reset
		.uas_address          (max2_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (max2_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (max2_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (max2_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (max2_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (max2_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (max2_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (max2_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (max2_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (max2_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (max2_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (max2_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (max2_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (max2_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (max2_tcm_request),                                      //      .request
		.tcm_grant            (max2_tcm_grant),                                        //      .grant
		.tcm_address_out      (max2_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (max2_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (max2_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (max2_tcm_data_in)                                       //      .data_in
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (29),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                   (pll_c0_out),                                                         //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                 //                     reset.reset
		.uav_address           (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_data_master_read),                                               //                          .read
		.av_readdata           (cpu_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cpu_data_master_write),                                              //                          .write
		.av_writedata          (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (29),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                   (pll_c0_out),                                                                //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                        //                     reset.reset
		.uav_address           (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_byteenable         (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_write              (1'b0),                                                                      //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_descriptor_read_translator (
		.clk                   (pll_c0_out),                                                                  //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                     reset.reset
		.uav_address           (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_rx_descriptor_read_read),                                               //                          .read
		.av_readdata           (sgdma_rx_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_rx_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_descriptor_write_translator (
		.clk                   (pll_c0_out),                                                                   //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                           //                     reset.reset
		.uav_address           (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (sgdma_rx_descriptor_write_write),                                              //                          .write
		.av_writedata          (sgdma_rx_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_descriptor_read_translator (
		.clk                   (pll_c0_out),                                                                  //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                     reset.reset
		.uav_address           (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_tx_descriptor_read_read),                                               //                          .read
		.av_readdata           (sgdma_tx_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_tx_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_descriptor_write_translator (
		.clk                   (pll_c0_out),                                                                   //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                           //                     reset.reset
		.uav_address           (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (sgdma_tx_descriptor_write_write),                                              //                          .write
		.av_writedata          (sgdma_tx_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                   (pll_c0_out),                                                                       //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                               //                    reset.reset
		.uav_address           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) descriptor_memory_s1_translator (
		.clk                   (pll_c0_out),                                                                      //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                              //                    reset.reset
		.uav_address           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (descriptor_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (descriptor_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_rx_csr_translator (
		.clk                   (pll_c0_out),                                                              //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sgdma_rx_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sgdma_rx_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sgdma_rx_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sgdma_rx_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sgdma_rx_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_tx_csr_translator (
		.clk                   (pll_c0_out),                                                              //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sgdma_tx_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sgdma_tx_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sgdma_tx_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sgdma_tx_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sgdma_tx_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tse_mac_control_port_translator (
		.clk                   (pll_c0_out),                                                                      //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                              //                    reset.reset
		.uav_address           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (tse_mac_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (tse_mac_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (tse_mac_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (tse_mac_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (tse_mac_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sls_sdhc_control_translator (
		.clk                   (clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sls_sdhc_control_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sls_sdhc_control_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sls_sdhc_control_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sls_sdhc_control_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sls_sdhc_control_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (sls_sdhc_control_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sls_sdhc_control_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (27),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pipeline_bridge_before_tristate_bridge_s0_translator (
		.clk                   (pll_c0_out),                                                                                           //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                                   //                    reset.reset
		.uav_address           (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                                     //              (terminated)
		.av_lock               (),                                                                                                     //              (terminated)
		.av_chipselect         (),                                                                                                     //              (terminated)
		.av_clken              (),                                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (27),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_ddr_clock_bridge_s0_translator (
		.clk                   (pll_c0_out),                                                                         //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (cpu_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (26),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_ddr_1_clock_bridge_s0_translator (
		.clk                   (pll_c0_out),                                                                           //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (cpu_ddr_1_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_chipselect         (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) slow_peripheral_bridge_s0_translator (
		.clk                   (pll_c0_out),                                                                           //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_chipselect         (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) lcd_sgdma_descriptor_read_translator (
		.clk                   (ddr2_sdram_phy_clk_out),                                                       //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                           //                     reset.reset
		.uav_address           (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (lcd_sgdma_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (lcd_sgdma_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (lcd_sgdma_descriptor_read_read),                                               //                          .read
		.av_readdata           (lcd_sgdma_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (lcd_sgdma_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_write              (1'b0),                                                                         //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                         //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) lcd_sgdma_descriptor_write_translator (
		.clk                   (ddr2_sdram_phy_clk_out),                                                        //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                            //                     reset.reset
		.uav_address           (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (lcd_sgdma_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (lcd_sgdma_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (lcd_sgdma_descriptor_write_write),                                              //                          .write
		.av_writedata          (lcd_sgdma_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                          //               (terminated)
		.av_byteenable         (4'b1111),                                                                       //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                          //               (terminated)
		.av_begintransfer      (1'b0),                                                                          //               (terminated)
		.av_chipselect         (1'b0),                                                                          //               (terminated)
		.av_read               (1'b0),                                                                          //               (terminated)
		.av_readdata           (),                                                                              //               (terminated)
		.av_readdatavalid      (),                                                                              //               (terminated)
		.av_lock               (1'b0),                                                                          //               (terminated)
		.av_debugaccess        (1'b0),                                                                          //               (terminated)
		.uav_clken             (),                                                                              //               (terminated)
		.av_clken              (1'b1)                                                                           //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (64),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (8),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (4),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (8),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) lcd_sgdma_m_read_translator (
		.clk                   (ddr2_sdram_phy_clk_out),                                               //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                   //                     reset.reset
		.uav_address           (lcd_sgdma_m_read_translator_avalon_universal_master_0_address),        // avalon_universal_master_0.address
		.uav_burstcount        (lcd_sgdma_m_read_translator_avalon_universal_master_0_burstcount),     //                          .burstcount
		.uav_read              (lcd_sgdma_m_read_translator_avalon_universal_master_0_read),           //                          .read
		.uav_write             (lcd_sgdma_m_read_translator_avalon_universal_master_0_write),          //                          .write
		.uav_waitrequest       (lcd_sgdma_m_read_translator_avalon_universal_master_0_waitrequest),    //                          .waitrequest
		.uav_readdatavalid     (lcd_sgdma_m_read_translator_avalon_universal_master_0_readdatavalid),  //                          .readdatavalid
		.uav_byteenable        (lcd_sgdma_m_read_translator_avalon_universal_master_0_byteenable),     //                          .byteenable
		.uav_readdata          (lcd_sgdma_m_read_translator_avalon_universal_master_0_readdata),       //                          .readdata
		.uav_writedata         (lcd_sgdma_m_read_translator_avalon_universal_master_0_writedata),      //                          .writedata
		.uav_lock              (lcd_sgdma_m_read_translator_avalon_universal_master_0_lock),           //                          .lock
		.uav_debugaccess       (lcd_sgdma_m_read_translator_avalon_universal_master_0_debugaccess),    //                          .debugaccess
		.av_address            (lcd_sgdma_m_read_address),                                             //      avalon_anti_master_0.address
		.av_waitrequest        (lcd_sgdma_m_read_waitrequest),                                         //                          .waitrequest
		.av_read               (lcd_sgdma_m_read_read),                                                //                          .read
		.av_readdata           (lcd_sgdma_m_read_readdata),                                            //                          .readdata
		.av_readdatavalid      (lcd_sgdma_m_read_readdatavalid),                                       //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_byteenable         (8'b11111111),                                                          //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_write              (1'b0),                                                                 //               (terminated)
		.av_writedata          (64'b0000000000000000000000000000000000000000000000000000000000000000), //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.av_debugaccess        (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (64),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (8),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (4),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (8),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sdhc_ddr_clock_bridge_m0_translator (
		.clk                   (ddr2_sdram_phy_clk_out),                                                      //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                          //                     reset.reset
		.uav_address           (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sdhc_ddr_clock_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sdhc_ddr_clock_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (sdhc_ddr_clock_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (sdhc_ddr_clock_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (sdhc_ddr_clock_bridge_m0_read),                                               //                          .read
		.av_readdata           (sdhc_ddr_clock_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (sdhc_ddr_clock_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (sdhc_ddr_clock_bridge_m0_write),                                              //                          .write
		.av_writedata          (sdhc_ddr_clock_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (sdhc_ddr_clock_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_ddr_clock_bridge_m0_translator (
		.clk                   (ddr2_sdram_phy_clk_out),                                                     //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                         //                     reset.reset
		.uav_address           (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_ddr_clock_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_ddr_clock_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (cpu_ddr_clock_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (cpu_ddr_clock_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (cpu_ddr_clock_bridge_m0_read),                                               //                          .read
		.av_readdata           (cpu_ddr_clock_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_ddr_clock_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cpu_ddr_clock_bridge_m0_write),                                              //                          .write
		.av_writedata          (cpu_ddr_clock_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_ddr_clock_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                       //               (terminated)
		.av_begintransfer      (1'b0),                                                                       //               (terminated)
		.av_chipselect         (1'b0),                                                                       //               (terminated)
		.av_lock               (1'b0),                                                                       //               (terminated)
		.uav_clken             (),                                                                           //               (terminated)
		.av_clken              (1'b1)                                                                        //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) tse_ddr_clock_bridge_m0_translator (
		.clk                   (ddr2_sdram_phy_clk_out),                                                     //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                         //                     reset.reset
		.uav_address           (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (tse_ddr_clock_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (tse_ddr_clock_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (tse_ddr_clock_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (tse_ddr_clock_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (tse_ddr_clock_bridge_m0_read),                                               //                          .read
		.av_readdata           (tse_ddr_clock_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (tse_ddr_clock_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (tse_ddr_clock_bridge_m0_write),                                              //                          .write
		.av_writedata          (tse_ddr_clock_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (tse_ddr_clock_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                       //               (terminated)
		.av_begintransfer      (1'b0),                                                                       //               (terminated)
		.av_chipselect         (1'b0),                                                                       //               (terminated)
		.av_lock               (1'b0),                                                                       //               (terminated)
		.uav_clken             (),                                                                           //               (terminated)
		.av_clken              (1'b1)                                                                        //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (23),
		.AV_DATA_W                      (64),
		.UAV_DATA_W                     (64),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (8),
		.UAV_BYTEENABLE_W               (8),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (4),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (8),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_sdram_s1_translator (
		.clk                   (ddr2_sdram_phy_clk_out),                                                   //                      clk.clk
		.reset                 (~ddr2_sdram_reset_request_n_reset),                                        //                    reset.reset
		.uav_address           (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ddr2_sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ddr2_sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ddr2_sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ddr2_sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ddr2_sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer (ddr2_sdram_s1_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount         (ddr2_sdram_s1_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (ddr2_sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (ddr2_sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (~ddr2_sdram_s1_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_sgdma_csr_translator (
		.clk                   (ddr2_sdram_phy_clk_out),                                                   //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                       //                    reset.reset
		.uav_address           (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (lcd_sgdma_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (lcd_sgdma_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (lcd_sgdma_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (lcd_sgdma_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (lcd_sgdma_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (lcd_sgdma_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sls_sdhc_read_master_translator (
		.clk                   (clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                     reset.reset
		.uav_address           (sls_sdhc_read_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sls_sdhc_read_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sls_sdhc_read_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sls_sdhc_read_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sls_sdhc_read_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sls_sdhc_read_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sls_sdhc_read_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sls_sdhc_read_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sls_sdhc_read_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sls_sdhc_read_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sls_sdhc_read_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sls_sdhc_read_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sls_sdhc_read_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (sls_sdhc_read_master_byteenable),                                         //                          .byteenable
		.av_read               (~sls_sdhc_read_master_read),                                              //                          .read
		.av_readdata           (sls_sdhc_read_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (sls_sdhc_read_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                    //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                    //               (terminated)
		.av_begintransfer      (1'b0),                                                                    //               (terminated)
		.av_chipselect         (1'b0),                                                                    //               (terminated)
		.av_write              (1'b0),                                                                    //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                    //               (terminated)
		.av_lock               (1'b0),                                                                    //               (terminated)
		.av_debugaccess        (1'b0),                                                                    //               (terminated)
		.uav_clken             (),                                                                        //               (terminated)
		.av_clken              (1'b1)                                                                     //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sls_sdhc_write_master_translator (
		.clk                   (clk),                                                                      //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                     reset.reset
		.uav_address           (sls_sdhc_write_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sls_sdhc_write_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sls_sdhc_write_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sls_sdhc_write_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sls_sdhc_write_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sls_sdhc_write_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sls_sdhc_write_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sls_sdhc_write_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sls_sdhc_write_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sls_sdhc_write_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sls_sdhc_write_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sls_sdhc_write_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sls_sdhc_write_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (sls_sdhc_write_master_byteenable),                                         //                          .byteenable
		.av_chipselect         (sls_sdhc_write_master_chipselect),                                         //                          .chipselect
		.av_write              (~sls_sdhc_write_master_write),                                             //                          .write
		.av_writedata          (sls_sdhc_write_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                     //               (terminated)
		.av_begintransfer      (1'b0),                                                                     //               (terminated)
		.av_read               (1'b0),                                                                     //               (terminated)
		.av_readdata           (),                                                                         //               (terminated)
		.av_readdatavalid      (),                                                                         //               (terminated)
		.av_lock               (1'b0),                                                                     //               (terminated)
		.av_debugaccess        (1'b0),                                                                     //               (terminated)
		.uav_clken             (),                                                                         //               (terminated)
		.av_clken              (1'b1)                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (26),
		.AV_DATA_W                      (64),
		.UAV_DATA_W                     (64),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (8),
		.UAV_BYTEENABLE_W               (8),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (4),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (8),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdhc_ddr_clock_bridge_s0_translator (
		.clk                   (pll_c0_out),                                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (sdhc_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_chipselect         (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_ddr_1_clock_bridge_m0_translator (
		.clk                   (ddr2_sdram_1_phy_clk_out),                                                     //                       clk.clk
		.reset                 (rst_controller_005_reset_out_reset),                                           //                     reset.reset
		.uav_address           (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_ddr_1_clock_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_ddr_1_clock_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (cpu_ddr_1_clock_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (cpu_ddr_1_clock_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (cpu_ddr_1_clock_bridge_m0_read),                                               //                          .read
		.av_readdata           (cpu_ddr_1_clock_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_ddr_1_clock_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cpu_ddr_1_clock_bridge_m0_write),                                              //                          .write
		.av_writedata          (cpu_ddr_1_clock_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_ddr_1_clock_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (2),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (4),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (1),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_sdram_1_s1_translator (
		.clk                   (ddr2_sdram_1_phy_clk_out),                                                   //                      clk.clk
		.reset                 (~ddr2_sdram_1_reset_request_n_reset),                                        //                    reset.reset
		.uav_address           (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount         (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (ddr2_sdram_1_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (~ddr2_sdram_1_s1_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_chipselect         (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (10),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) slow_peripheral_bridge_m0_translator (
		.clk                   (pll_c2_out),                                                                   //                       clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                           //                     reset.reset
		.uav_address           (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (slow_peripheral_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (slow_peripheral_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (slow_peripheral_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (slow_peripheral_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (slow_peripheral_bridge_m0_read),                                               //                          .read
		.av_readdata           (slow_peripheral_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (slow_peripheral_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (slow_peripheral_bridge_m0_write),                                              //                          .write
		.av_writedata          (slow_peripheral_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (slow_peripheral_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button_pio_s1_translator (
		.clk                   (pll_c2_out),                                                               //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                       //                    reset.reset
		.uav_address           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (button_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (button_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (button_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (button_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (button_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_res_timer_s1_translator (
		.clk                   (pll_c2_out),                                                                   //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                           //                    reset.reset
		.uav_address           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (high_res_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (high_res_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (high_res_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (high_res_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (high_res_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                   (pll_c2_out),                                                                             //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart1_s1_translator (
		.clk                   (pll_c2_out),                                                          //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                  //                    reset.reset
		.uav_address           (uart1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (uart1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (uart1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (uart1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (uart1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (uart1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (uart1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (uart1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (uart1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (uart1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (uart1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (uart1_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (uart1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (uart1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (uart1_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect         (uart1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_byteenable         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_pio_s1_translator (
		.clk                   (pll_c2_out),                                                            //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                    //                    reset.reset
		.uav_address           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (led_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (led_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (led_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (led_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (led_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) performance_counter_control_slave_translator (
		.clk                   (pll_c2_out),                                                                                   //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (performance_counter_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (performance_counter_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (performance_counter_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (performance_counter_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_read               (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                             //              (terminated)
		.av_byteenable         (),                                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_lock               (),                                                                                             //              (terminated)
		.av_chipselect         (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_debugaccess        (),                                                                                             //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pll_s1_translator (
		.clk                   (clk),                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address           (pll_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pll_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pll_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pll_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pll_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pll_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pll_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pll_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pll_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pll_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pll_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pll_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pll_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pll_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pll_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pll_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pll_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                  //              (terminated)
		.av_burstcount         (),                                                                  //              (terminated)
		.av_byteenable         (),                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                              //              (terminated)
		.av_writebyteenable    (),                                                                  //              (terminated)
		.av_lock               (),                                                                  //              (terminated)
		.av_clken              (),                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                              //              (terminated)
		.av_debugaccess        (),                                                                  //              (terminated)
		.av_outputenable       ()                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sys_clk_timer_s1_translator (
		.clk                   (pll_c2_out),                                                                  //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                          //                    reset.reset
		.uav_address           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sys_clk_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                   (pll_c2_out),                                                                     //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                             //                    reset.reset
		.uav_address           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_writedata          (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_i2c_en_s1_translator (
		.clk                   (pll_c2_out),                                                               //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                       //                    reset.reset
		.uav_address           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (lcd_i2c_en_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (lcd_i2c_en_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (lcd_i2c_en_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (lcd_i2c_en_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (lcd_i2c_en_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_i2c_scl_s1_translator (
		.clk                   (pll_c2_out),                                                                //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                        //                    reset.reset
		.uav_address           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_byteenable         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_i2c_sdat_s1_translator (
		.clk                   (pll_c2_out),                                                                 //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                         //                    reset.reset
		.uav_address           (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (lcd_i2c_sdat_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                           //              (terminated)
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_burstcount         (),                                                                           //              (terminated)
		.av_byteenable         (),                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                       //              (terminated)
		.av_waitrequest        (1'b0),                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_id_eeprom_dat_s1_translator (
		.clk                   (pll_c2_out),                                                                      //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                              //                    reset.reset
		.uav_address           (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pio_id_eeprom_dat_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_id_eeprom_scl_s1_translator (
		.clk                   (pll_c2_out),                                                                      //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                              //                    reset.reset
		.uav_address           (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pio_id_eeprom_scl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) touch_panel_pen_irq_n_s1_translator (
		.clk                   (pll_c2_out),                                                                          //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                    //              (terminated)
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_byteenable         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) touch_panel_spi_spi_control_port_translator (
		.clk                   (pll_c2_out),                                                                                  //                      clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                                                          //                    reset.reset
		.uav_address           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                                            //              (terminated)
		.av_burstcount         (),                                                                                            //              (terminated)
		.av_byteenable         (),                                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                                            //              (terminated)
		.av_lock               (),                                                                                            //              (terminated)
		.av_clken              (),                                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                                        //              (terminated)
		.av_debugaccess        (),                                                                                            //              (terminated)
		.av_outputenable       ()                                                                                             //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_m_write_translator (
		.clk                   (pll_c0_out),                                                          //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                  //                     reset.reset
		.uav_address           (sgdma_rx_m_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_m_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_m_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_m_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_m_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_m_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_m_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_m_write_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (sgdma_rx_m_write_byteenable),                                         //                          .byteenable
		.av_write              (sgdma_rx_m_write_write),                                              //                          .write
		.av_writedata          (sgdma_rx_m_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                //               (terminated)
		.av_begintransfer      (1'b0),                                                                //               (terminated)
		.av_chipselect         (1'b0),                                                                //               (terminated)
		.av_read               (1'b0),                                                                //               (terminated)
		.av_readdata           (),                                                                    //               (terminated)
		.av_readdatavalid      (),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                //               (terminated)
		.av_debugaccess        (1'b0),                                                                //               (terminated)
		.uav_clken             (),                                                                    //               (terminated)
		.av_clken              (1'b1)                                                                 //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_m_read_translator (
		.clk                   (pll_c0_out),                                                         //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                 //                     reset.reset
		.uav_address           (sgdma_tx_m_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_m_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_m_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_m_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_m_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_m_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_m_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_m_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_tx_m_read_read),                                               //                          .read
		.av_readdata           (sgdma_tx_m_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_tx_m_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_write              (1'b0),                                                               //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (26),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tse_ddr_clock_bridge_s0_translator (
		.clk                   (pll_c0_out),                                                                         //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (tse_ddr_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (27),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) pipeline_bridge_before_tristate_bridge_m0_translator (
		.clk                   (pll_c0_out),                                                                                   //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                           //                     reset.reset
		.uav_address           (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (pipeline_bridge_before_tristate_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (pipeline_bridge_before_tristate_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (pipeline_bridge_before_tristate_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (pipeline_bridge_before_tristate_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read               (pipeline_bridge_before_tristate_bridge_m0_read),                                               //                          .read
		.av_readdata           (pipeline_bridge_before_tristate_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (pipeline_bridge_before_tristate_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (pipeline_bridge_before_tristate_bridge_m0_write),                                              //                          .write
		.av_writedata          (pipeline_bridge_before_tristate_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (pipeline_bridge_before_tristate_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                                         //               (terminated)
		.av_lock               (1'b0),                                                                                         //               (terminated)
		.uav_clken             (),                                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                                          //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (26),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (2),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ext_flash_uas_translator (
		.clk                   (pll_c0_out),                                                               //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ext_flash_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ext_flash_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ext_flash_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ext_flash_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ext_flash_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (ext_flash_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (ext_flash_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (ext_flash_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (ext_flash_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (ext_flash_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (3),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) max2_uas_translator (
		.clk                   (pll_c0_out),                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address           (max2_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (max2_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (max2_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (max2_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (max2_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (max2_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (max2_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (max2_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (max2_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (max2_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (max2_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (max2_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (max2_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (max2_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (max2_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (max2_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (max2_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (max2_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (max2_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (max2_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (max2_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (max2_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_chipselect         (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                  //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.av_address       (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                       //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                        //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                     //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                 //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                        //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (3)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                         //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.av_address       (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                          //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                           //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                        //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                    //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                           //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7)
	) sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                           //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_002_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_002_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_002_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_002_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_002_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_002_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7)
	) sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                            //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_003_rsp_src_valid),                                                             //        rp.valid
		.rp_data          (limiter_003_rsp_src_data),                                                              //          .data
		.rp_channel       (limiter_003_rsp_src_channel),                                                           //          .channel
		.rp_startofpacket (limiter_003_rsp_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (limiter_003_rsp_src_endofpacket),                                                       //          .endofpacket
		.rp_ready         (limiter_003_rsp_src_ready)                                                              //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (5),
		.BURSTWRAP_VALUE           (7)
	) sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                           //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_004_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_004_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_004_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_004_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_004_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_004_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (6),
		.BURSTWRAP_VALUE           (7)
	) sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                            //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_005_rsp_src_valid),                                                             //        rp.valid
		.rp_data          (limiter_005_rsp_src_data),                                                              //          .data
		.rp_channel       (limiter_005_rsp_src_channel),                                                           //          .channel
		.rp_startofpacket (limiter_005_rsp_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (limiter_005_rsp_src_endofpacket),                                                       //          .endofpacket
		.rp_ready         (limiter_005_rsp_src_ready)                                                              //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                              //                .channel
		.rf_sink_ready           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sgdma_rx_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                       //                .channel
		.rf_sink_ready           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sgdma_tx_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src3_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_src3_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_src3_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_src3_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src3_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src3_channel),                                                       //                .channel
		.rf_sink_ready           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) tse_mac_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src4_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_src4_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_src4_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_src4_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src4_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src4_channel),                                                               //                .channel
		.rf_sink_ready           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sls_sdhc_control_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sls_sdhc_control_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                     //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                     //                .valid
		.cp_data                 (crosser_out_data),                                                                      //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                               //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                   //                .channel
		.rf_sink_ready           (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_startofpacket  (1'b0),                                                                            // (terminated)
		.in_endofpacket    (1'b0),                                                                            // (terminated)
		.out_startofpacket (),                                                                                // (terminated)
		.out_endofpacket   (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_006_src_ready),                                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_006_src_valid),                                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_006_src_data),                                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_006_src_startofpacket),                                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_006_src_endofpacket),                                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_006_src_channel),                                                                                   //                .channel
		.rf_sink_ready           (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (6),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                                           // (terminated)
		.csr_readdata      (),                                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                           // (terminated)
		.almost_full_data  (),                                                                                                               // (terminated)
		.almost_empty_data (),                                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                                           // (terminated)
		.out_empty         (),                                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                                           // (terminated)
		.out_error         (),                                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                                           // (terminated)
		.out_channel       ()                                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src7_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_src7_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_src7_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_src7_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src7_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src7_channel),                                                                  //                .channel
		.rf_sink_ready           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (73),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (73),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src9_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_src9_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_src9_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_src9_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src9_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src9_channel),                                                                    //                .channel
		.rf_sink_ready           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (81),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (1),
		.BURSTWRAP_VALUE           (15)
	) lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (ddr2_sdram_phy_clk_out),                                                                //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_006_rsp_src_valid),                                                             //        rp.valid
		.rp_data          (limiter_006_rsp_src_data),                                                              //          .data
		.rp_channel       (limiter_006_rsp_src_channel),                                                           //          .channel
		.rp_startofpacket (limiter_006_rsp_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (limiter_006_rsp_src_endofpacket),                                                       //          .endofpacket
		.rp_ready         (limiter_006_rsp_src_ready)                                                              //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (2),
		.BURSTWRAP_VALUE           (15)
	) lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (ddr2_sdram_phy_clk_out),                                                                 //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.av_address       (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_007_rsp_src_valid),                                                              //        rp.valid
		.rp_data          (limiter_007_rsp_src_data),                                                               //          .data
		.rp_channel       (limiter_007_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket (limiter_007_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket   (limiter_007_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready         (limiter_007_rsp_src_ready)                                                               //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (124),
		.PKT_PROTECTION_L          (124),
		.PKT_BEGIN_BURST           (117),
		.PKT_BURSTWRAP_H           (116),
		.PKT_BURSTWRAP_L           (113),
		.PKT_BYTE_CNT_H            (112),
		.PKT_BYTE_CNT_L            (109),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (120),
		.PKT_SRC_ID_L              (118),
		.PKT_DEST_ID_H             (123),
		.PKT_DEST_ID_L             (121),
		.ST_DATA_W                 (125),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (4),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (15)
	) lcd_sgdma_m_read_translator_avalon_universal_master_0_agent (
		.clk              (ddr2_sdram_phy_clk_out),                                                       //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                           // clk_reset.reset
		.av_address       (lcd_sgdma_m_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (lcd_sgdma_m_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (lcd_sgdma_m_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (lcd_sgdma_m_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (lcd_sgdma_m_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (lcd_sgdma_m_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (lcd_sgdma_m_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (lcd_sgdma_m_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (lcd_sgdma_m_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (lcd_sgdma_m_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (lcd_sgdma_m_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_008_rsp_src_valid),                                                    //        rp.valid
		.rp_data          (limiter_008_rsp_src_data),                                                     //          .data
		.rp_channel       (limiter_008_rsp_src_channel),                                                  //          .channel
		.rp_startofpacket (limiter_008_rsp_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (limiter_008_rsp_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (limiter_008_rsp_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (124),
		.PKT_PROTECTION_L          (124),
		.PKT_BEGIN_BURST           (117),
		.PKT_BURSTWRAP_H           (116),
		.PKT_BURSTWRAP_L           (113),
		.PKT_BYTE_CNT_H            (112),
		.PKT_BYTE_CNT_L            (109),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (120),
		.PKT_SRC_ID_L              (118),
		.PKT_DEST_ID_H             (123),
		.PKT_DEST_ID_L             (121),
		.ST_DATA_W                 (125),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (4),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (15)
	) sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (ddr2_sdram_phy_clk_out),                                                               //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_009_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_009_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_009_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_009_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_009_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_009_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (5),
		.BURSTWRAP_VALUE           (15)
	) cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (ddr2_sdram_phy_clk_out),                                                              //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.av_address       (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_010_rsp_src_valid),                                                           //        rp.valid
		.rp_data          (limiter_010_rsp_src_data),                                                            //          .data
		.rp_channel       (limiter_010_rsp_src_channel),                                                         //          .channel
		.rp_startofpacket (limiter_010_rsp_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket   (limiter_010_rsp_src_endofpacket),                                                     //          .endofpacket
		.rp_ready         (limiter_010_rsp_src_ready)                                                            //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (6),
		.BURSTWRAP_VALUE           (15)
	) tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (ddr2_sdram_phy_clk_out),                                                              //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.av_address       (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_011_rsp_src_valid),                                                           //        rp.valid
		.rp_data          (limiter_011_rsp_src_data),                                                            //          .data
		.rp_channel       (limiter_011_rsp_src_channel),                                                         //          .channel
		.rp_startofpacket (limiter_011_rsp_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket   (limiter_011_rsp_src_endofpacket),                                                     //          .endofpacket
		.rp_ready         (limiter_011_rsp_src_ready)                                                            //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (117),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_SRC_ID_H              (120),
		.PKT_SRC_ID_L              (118),
		.PKT_DEST_ID_H             (123),
		.PKT_DEST_ID_L             (121),
		.PKT_BURSTWRAP_H           (116),
		.PKT_BURSTWRAP_L           (113),
		.PKT_BYTE_CNT_H            (112),
		.PKT_BYTE_CNT_L            (109),
		.PKT_PROTECTION_H          (124),
		.PKT_PROTECTION_L          (124),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (125),
		.AVS_BURSTCOUNT_W          (4),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ddr2_sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (ddr2_sdram_phy_clk_out),                                                             //             clk.clk
		.reset                   (~ddr2_sdram_reset_request_n_reset),                                                  //       clk_reset.reset
		.m0_address              (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_010_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_010_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_010_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_010_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_010_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_010_src_channel),                                                       //                .channel
		.rf_sink_ready           (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (126),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ddr2_sdram_phy_clk_out),                                                             //       clk.clk
		.reset             (~ddr2_sdram_reset_request_n_reset),                                                  // clk_reset.reset
		.in_data           (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) lcd_sgdma_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (ddr2_sdram_phy_clk_out),                                                             //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_010_src1_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_010_src1_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_010_src1_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_010_src1_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_010_src1_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_010_src1_channel),                                                    //                .channel
		.rf_sink_ready           (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ddr2_sdram_phy_clk_out),                                                             //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (1),
		.BURSTWRAP_VALUE           (15)
	) sls_sdhc_read_master_translator_avalon_universal_master_0_agent (
		.clk              (clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (sls_sdhc_read_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sls_sdhc_read_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sls_sdhc_read_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sls_sdhc_read_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sls_sdhc_read_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sls_sdhc_read_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sls_sdhc_read_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sls_sdhc_read_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sls_sdhc_read_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sls_sdhc_read_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sls_sdhc_read_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (crosser_004_out_valid),                                                            //        rp.valid
		.rp_data          (crosser_004_out_data),                                                             //          .data
		.rp_channel       (crosser_004_out_channel),                                                          //          .channel
		.rp_startofpacket (crosser_004_out_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (crosser_004_out_endofpacket),                                                      //          .endofpacket
		.rp_ready         (crosser_004_out_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (2),
		.BURSTWRAP_VALUE           (15)
	) sls_sdhc_write_master_translator_avalon_universal_master_0_agent (
		.clk              (clk),                                                                               //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (sls_sdhc_write_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sls_sdhc_write_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sls_sdhc_write_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sls_sdhc_write_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sls_sdhc_write_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sls_sdhc_write_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sls_sdhc_write_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sls_sdhc_write_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sls_sdhc_write_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sls_sdhc_write_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sls_sdhc_write_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (crosser_005_out_valid),                                                             //        rp.valid
		.rp_data          (crosser_005_out_data),                                                              //          .data
		.rp_channel       (crosser_005_out_channel),                                                           //          .channel
		.rp_startofpacket (crosser_005_out_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (crosser_005_out_endofpacket),                                                       //          .endofpacket
		.rp_ready         (crosser_005_out_ready)                                                              //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (117),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_SRC_ID_H              (119),
		.PKT_SRC_ID_L              (118),
		.PKT_DEST_ID_H             (121),
		.PKT_DEST_ID_L             (120),
		.PKT_BURSTWRAP_H           (116),
		.PKT_BURSTWRAP_L           (113),
		.PKT_BYTE_CNT_H            (112),
		.PKT_BYTE_CNT_L            (109),
		.PKT_PROTECTION_H          (122),
		.PKT_PROTECTION_L          (122),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (123),
		.AVS_BURSTCOUNT_W          (4),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (width_adapter_008_src_ready),                                                                   //              cp.ready
		.cp_valid                (width_adapter_008_src_valid),                                                                   //                .valid
		.cp_data                 (width_adapter_008_src_data),                                                                    //                .data
		.cp_startofpacket        (width_adapter_008_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (width_adapter_008_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (width_adapter_008_src_channel),                                                                 //                .channel
		.rf_sink_ready           (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (124),
		.FIFO_DEPTH          (73),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (64),
		.FIFO_DEPTH          (128),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c0_out),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                                    // (terminated)
		.out_startofpacket (),                                                                                        // (terminated)
		.out_endofpacket   (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (78),
		.PKT_BEGIN_BURST           (75),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (77),
		.PKT_DEST_ID_L             (77),
		.ST_DATA_W                 (79),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (15)
	) cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (ddr2_sdram_1_phy_clk_out),                                                              //       clk.clk
		.reset            (rst_controller_005_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_013_src0_valid),                                                         //        rp.valid
		.rp_data          (rsp_xbar_demux_013_src0_data),                                                          //          .data
		.rp_channel       (rsp_xbar_demux_013_src0_channel),                                                       //          .channel
		.rp_startofpacket (rsp_xbar_demux_013_src0_startofpacket),                                                 //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),                                                   //          .endofpacket
		.rp_ready         (rsp_xbar_demux_013_src0_ready)                                                          //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (77),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (78),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (79),
		.AVS_BURSTCOUNT_W          (4),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (ddr2_sdram_1_phy_clk_out),                                                             //             clk.clk
		.reset                   (~ddr2_sdram_1_reset_request_n_reset),                                                  //       clk_reset.reset
		.m0_address              (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_014_src0_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_014_src0_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_014_src0_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_014_src0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_014_src0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_014_src0_channel),                                                      //                .channel
		.rf_sink_ready           (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (80),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ddr2_sdram_1_phy_clk_out),                                                             //       clk.clk
		.reset             (~ddr2_sdram_1_reset_request_n_reset),                                                  // clk_reset.reset
		.in_data           (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.PKT_BEGIN_BURST           (57),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.ST_DATA_W                 (69),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7)
	) slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (pll_c2_out),                                                                            //       clk.clk
		.reset            (rst_controller_004_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_012_rsp_src_valid),                                                             //        rp.valid
		.rp_data          (limiter_012_rsp_src_data),                                                              //          .data
		.rp_channel       (limiter_012_rsp_src_channel),                                                           //          .channel
		.rp_startofpacket (limiter_012_rsp_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (limiter_012_rsp_src_endofpacket),                                                       //          .endofpacket
		.rp_ready         (limiter_012_rsp_src_ready)                                                              //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) button_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                         //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src0_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src0_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_015_src0_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src0_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src0_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src0_channel),                                                    //                .channel
		.rf_sink_ready           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                         //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) high_res_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                             //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src1_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src1_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_015_src1_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src1_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src1_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src1_channel),                                                        //                .channel
		.rf_sink_ready           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                             //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                       //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src2_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src2_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_015_src2_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src2_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src2_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src2_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                       //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) uart1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                    //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (uart1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src3_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src3_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_015_src3_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src3_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src3_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src3_channel),                                               //                .channel
		.rf_sink_ready           (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                    //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                            // clk_reset.reset
		.in_data           (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) led_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                      //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src4_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src4_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_015_src4_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src4_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src4_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src4_channel),                                                 //                .channel
		.rf_sink_ready           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                      //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                              // clk_reset.reset
		.in_data           (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) performance_counter_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                             //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src5_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src5_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_015_src5_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src5_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src5_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src5_channel),                                                                        //                .channel
		.rf_sink_ready           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                             //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pll_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (pll_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pll_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pll_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pll_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pll_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pll_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pll_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pll_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pll_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pll_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pll_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pll_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pll_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pll_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pll_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pll_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_006_out_ready),                                                       //              cp.ready
		.cp_valid                (crosser_006_out_valid),                                                       //                .valid
		.cp_data                 (crosser_006_out_data),                                                        //                .data
		.cp_startofpacket        (crosser_006_out_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (crosser_006_out_endofpacket),                                                 //                .endofpacket
		.cp_channel              (crosser_006_out_channel),                                                     //                .channel
		.rf_sink_ready           (pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pll_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pll_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pll_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pll_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pll_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (pll_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pll_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pll_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pll_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pll_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pll_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.in_data           (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (pll_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                 // (terminated)
		.csr_read          (1'b0),                                                                  // (terminated)
		.csr_write         (1'b0),                                                                  // (terminated)
		.csr_readdata      (),                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                  // (terminated)
		.almost_full_data  (),                                                                      // (terminated)
		.almost_empty_data (),                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                  // (terminated)
		.out_startofpacket (),                                                                      // (terminated)
		.out_endofpacket   (),                                                                      // (terminated)
		.in_empty          (1'b0),                                                                  // (terminated)
		.out_empty         (),                                                                      // (terminated)
		.in_error          (1'b0),                                                                  // (terminated)
		.out_error         (),                                                                      // (terminated)
		.in_channel        (1'b0),                                                                  // (terminated)
		.out_channel       ()                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                            //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src7_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src7_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_015_src7_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src7_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src7_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src7_channel),                                                       //                .channel
		.rf_sink_ready           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                            //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                               //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src8_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src8_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_015_src8_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src8_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src8_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src8_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                               //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                         //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src9_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src9_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_015_src9_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src9_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src9_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src9_channel),                                                    //                .channel
		.rf_sink_ready           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                         //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                          //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src10_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src10_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_015_src10_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src10_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src10_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src10_channel),                                                    //                .channel
		.rf_sink_ready           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                          //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                           //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src11_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src11_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_015_src11_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src11_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src11_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src11_channel),                                                     //                .channel
		.rf_sink_ready           (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                           //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src12_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src12_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_015_src12_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src12_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src12_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src12_channel),                                                          //                .channel
		.rf_sink_ready           (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src13_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src13_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_015_src13_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src13_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src13_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src13_channel),                                                          //                .channel
		.rf_sink_ready           (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                    //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src14_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src14_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_015_src14_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src14_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src14_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src14_channel),                                                              //                .channel
		.rf_sink_ready           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                    //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (62),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                            //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_015_src15_ready),                                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_015_src15_valid),                                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_015_src15_data),                                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_015_src15_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_015_src15_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_015_src15_channel),                                                                      //                .channel
		.rf_sink_ready           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                            //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (82),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7)
	) sgdma_rx_m_write_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                   //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.av_address       (sgdma_rx_m_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_m_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_m_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_m_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_m_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_m_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_030_src0_valid),                                                //        rp.valid
		.rp_data          (rsp_xbar_demux_030_src0_data),                                                 //          .data
		.rp_channel       (rsp_xbar_demux_030_src0_channel),                                              //          .channel
		.rp_startofpacket (rsp_xbar_demux_030_src0_startofpacket),                                        //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_030_src0_endofpacket),                                          //          .endofpacket
		.rp_ready         (rsp_xbar_demux_030_src0_ready)                                                 //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (82),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7)
	) sgdma_tx_m_read_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                  //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.av_address       (sgdma_tx_m_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_m_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_m_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_m_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_m_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_m_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_030_src1_valid),                                               //        rp.valid
		.rp_data          (rsp_xbar_demux_030_src1_data),                                                //          .data
		.rp_channel       (rsp_xbar_demux_030_src1_channel),                                             //          .channel
		.rp_startofpacket (rsp_xbar_demux_030_src1_startofpacket),                                       //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_030_src1_endofpacket),                                         //          .endofpacket
		.rp_ready         (rsp_xbar_demux_030_src1_ready)                                                //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (84),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_030_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_030_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_030_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_030_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_030_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_030_src_channel),                                                                 //                .channel
		.rf_sink_ready           (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (73),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (79),
		.PKT_PROTECTION_L          (79),
		.PKT_BEGIN_BURST           (74),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (77),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7)
	) pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk              (pll_c0_out),                                                                                            //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                                    // clk_reset.reset
		.av_address       (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_013_rsp_src_valid),                                                                             //        rp.valid
		.rp_data          (limiter_013_rsp_src_data),                                                                              //          .data
		.rp_channel       (limiter_013_rsp_src_channel),                                                                           //          .channel
		.rp_startofpacket (limiter_013_rsp_src_startofpacket),                                                                     //          .startofpacket
		.rp_endofpacket   (limiter_013_rsp_src_endofpacket),                                                                       //          .endofpacket
		.rp_ready         (limiter_013_rsp_src_ready)                                                                              //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (56),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (57),
		.PKT_DEST_ID_H             (60),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (53),
		.PKT_BYTE_CNT_H            (52),
		.PKT_BYTE_CNT_L            (50),
		.PKT_PROTECTION_H          (61),
		.PKT_PROTECTION_L          (61),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (62),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ext_flash_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                      //                .channel
		.rf_sink_ready           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (63),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (75),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (79),
		.PKT_PROTECTION_L          (79),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) max2_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (max2_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (max2_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (max2_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (max2_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (max2_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (max2_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (max2_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (max2_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (max2_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (max2_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (max2_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (max2_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (max2_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (max2_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (max2_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (max2_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_018_src1_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_018_src1_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_018_src1_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_018_src1_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_018_src1_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_018_src1_channel),                                               //                .channel
		.rf_sink_ready           (max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (max2_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (max2_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (max2_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (max2_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (max2_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (max2_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (max2_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (max2_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (max2_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (max2_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (max2_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (max2_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (max2_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (max2_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (max2_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (max2_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (max2_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	application_selector_addr_router addr_router (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                       //          .valid
		.src_data           (addr_router_src_data),                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                  //          .endofpacket
	);

	application_selector_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                          //          .valid
		.src_data           (addr_router_001_src_data),                                                           //          .data
		.src_channel        (addr_router_001_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                     //          .endofpacket
	);

	application_selector_addr_router_002 addr_router_002 (
		.sink_ready         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                            //          .valid
		.src_data           (addr_router_002_src_data),                                                             //          .data
		.src_channel        (addr_router_002_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                       //          .endofpacket
	);

	application_selector_addr_router_002 addr_router_003 (
		.sink_ready         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                             //          .valid
		.src_data           (addr_router_003_src_data),                                                              //          .data
		.src_channel        (addr_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	application_selector_addr_router_002 addr_router_004 (
		.sink_ready         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                            //          .valid
		.src_data           (addr_router_004_src_data),                                                             //          .data
		.src_channel        (addr_router_004_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                       //          .endofpacket
	);

	application_selector_addr_router_002 addr_router_005 (
		.sink_ready         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                             //          .valid
		.src_data           (addr_router_005_src_data),                                                              //          .data
		.src_channel        (addr_router_005_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                        //          .endofpacket
	);

	application_selector_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	application_selector_id_router_001 id_router_001 (
		.sink_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                         //       src.ready
		.src_valid          (id_router_001_src_valid),                                                         //          .valid
		.src_data           (id_router_001_src_data),                                                          //          .data
		.src_channel        (id_router_001_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                    //          .endofpacket
	);

	application_selector_id_router_002 id_router_002 (
		.sink_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                 //       src.ready
		.src_valid          (id_router_002_src_valid),                                                 //          .valid
		.src_data           (id_router_002_src_data),                                                  //          .data
		.src_channel        (id_router_002_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                            //          .endofpacket
	);

	application_selector_id_router_002 id_router_003 (
		.sink_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                 //       src.ready
		.src_valid          (id_router_003_src_valid),                                                 //          .valid
		.src_data           (id_router_003_src_data),                                                  //          .data
		.src_channel        (id_router_003_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                            //          .endofpacket
	);

	application_selector_id_router_002 id_router_004 (
		.sink_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                         //       src.ready
		.src_valid          (id_router_004_src_valid),                                                         //          .valid
		.src_data           (id_router_004_src_data),                                                          //          .data
		.src_channel        (id_router_004_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                    //          .endofpacket
	);

	application_selector_id_router_002 id_router_005 (
		.sink_ready         (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sls_sdhc_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                     //       src.ready
		.src_valid          (id_router_005_src_valid),                                                     //          .valid
		.src_data           (id_router_005_src_data),                                                      //          .data
		.src_channel        (id_router_005_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                //          .endofpacket
	);

	application_selector_id_router id_router_006 (
		.sink_ready         (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pipeline_bridge_before_tristate_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                              //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                              //          .valid
		.src_data           (id_router_006_src_data),                                                                               //          .data
		.src_channel        (id_router_006_src_channel),                                                                            //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                                         //          .endofpacket
	);

	application_selector_id_router_002 id_router_007 (
		.sink_ready         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                            //       src.ready
		.src_valid          (id_router_007_src_valid),                                                            //          .valid
		.src_data           (id_router_007_src_data),                                                             //          .data
		.src_channel        (id_router_007_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                       //          .endofpacket
	);

	application_selector_id_router id_router_008 (
		.sink_ready         (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_ddr_1_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                              //       src.ready
		.src_valid          (id_router_008_src_valid),                                                              //          .valid
		.src_data           (id_router_008_src_data),                                                               //          .data
		.src_channel        (id_router_008_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                         //          .endofpacket
	);

	application_selector_id_router_002 id_router_009 (
		.sink_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                              //       src.ready
		.src_valid          (id_router_009_src_valid),                                                              //          .valid
		.src_data           (id_router_009_src_data),                                                               //          .data
		.src_channel        (id_router_009_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                         //          .endofpacket
	);

	application_selector_addr_router_006 addr_router_006 (
		.sink_ready         (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sdram_phy_clk_out),                                                                //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_006_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_006_src_valid),                                                             //          .valid
		.src_data           (addr_router_006_src_data),                                                              //          .data
		.src_channel        (addr_router_006_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_006_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_006_src_endofpacket)                                                        //          .endofpacket
	);

	application_selector_addr_router_006 addr_router_007 (
		.sink_ready         (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sdram_phy_clk_out),                                                                 //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_007_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_007_src_valid),                                                              //          .valid
		.src_data           (addr_router_007_src_data),                                                               //          .data
		.src_channel        (addr_router_007_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_007_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_007_src_endofpacket)                                                         //          .endofpacket
	);

	application_selector_addr_router_008 addr_router_008 (
		.sink_ready         (lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_sgdma_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sdram_phy_clk_out),                                                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (addr_router_008_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_008_src_valid),                                                    //          .valid
		.src_data           (addr_router_008_src_data),                                                     //          .data
		.src_channel        (addr_router_008_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_008_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_008_src_endofpacket)                                               //          .endofpacket
	);

	application_selector_addr_router_008 addr_router_009 (
		.sink_ready         (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdhc_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sdram_phy_clk_out),                                                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_009_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_009_src_valid),                                                            //          .valid
		.src_data           (addr_router_009_src_data),                                                             //          .data
		.src_channel        (addr_router_009_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_009_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_009_src_endofpacket)                                                       //          .endofpacket
	);

	application_selector_addr_router_010 addr_router_010 (
		.sink_ready         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sdram_phy_clk_out),                                                              //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (addr_router_010_src_ready),                                                           //       src.ready
		.src_valid          (addr_router_010_src_valid),                                                           //          .valid
		.src_data           (addr_router_010_src_data),                                                            //          .data
		.src_channel        (addr_router_010_src_channel),                                                         //          .channel
		.src_startofpacket  (addr_router_010_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (addr_router_010_src_endofpacket)                                                      //          .endofpacket
	);

	application_selector_addr_router_006 addr_router_011 (
		.sink_ready         (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tse_ddr_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sdram_phy_clk_out),                                                              //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (addr_router_011_src_ready),                                                           //       src.ready
		.src_valid          (addr_router_011_src_valid),                                                           //          .valid
		.src_data           (addr_router_011_src_data),                                                            //          .data
		.src_channel        (addr_router_011_src_channel),                                                         //          .channel
		.src_startofpacket  (addr_router_011_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (addr_router_011_src_endofpacket)                                                      //          .endofpacket
	);

	application_selector_id_router_010 id_router_010 (
		.sink_ready         (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sdram_phy_clk_out),                                                   //       clk.clk
		.reset              (~ddr2_sdram_reset_request_n_reset),                                        // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                  //       src.ready
		.src_valid          (id_router_010_src_valid),                                                  //          .valid
		.src_data           (id_router_010_src_data),                                                   //          .data
		.src_channel        (id_router_010_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                             //          .endofpacket
	);

	application_selector_id_router_011 id_router_011 (
		.sink_ready         (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_sgdma_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sdram_phy_clk_out),                                                   //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                  //       src.ready
		.src_valid          (id_router_011_src_valid),                                                  //          .valid
		.src_data           (id_router_011_src_data),                                                   //          .data
		.src_channel        (id_router_011_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                             //          .endofpacket
	);

	application_selector_addr_router_012 addr_router_012 (
		.sink_ready         (sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sls_sdhc_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_012_src_ready),                                                        //       src.ready
		.src_valid          (addr_router_012_src_valid),                                                        //          .valid
		.src_data           (addr_router_012_src_data),                                                         //          .data
		.src_channel        (addr_router_012_src_channel),                                                      //          .channel
		.src_startofpacket  (addr_router_012_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (addr_router_012_src_endofpacket)                                                   //          .endofpacket
	);

	application_selector_addr_router_012 addr_router_013 (
		.sink_ready         (sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sls_sdhc_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_013_src_ready),                                                         //       src.ready
		.src_valid          (addr_router_013_src_valid),                                                         //          .valid
		.src_data           (addr_router_013_src_data),                                                          //          .data
		.src_channel        (addr_router_013_src_channel),                                                       //          .channel
		.src_startofpacket  (addr_router_013_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (addr_router_013_src_endofpacket)                                                    //          .endofpacket
	);

	application_selector_id_router_012 id_router_012 (
		.sink_ready         (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdhc_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                             //       src.ready
		.src_valid          (id_router_012_src_valid),                                                             //          .valid
		.src_data           (id_router_012_src_data),                                                              //          .data
		.src_channel        (id_router_012_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                        //          .endofpacket
	);

	application_selector_addr_router_014 addr_router_014 (
		.sink_ready         (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_ddr_1_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sdram_1_phy_clk_out),                                                              //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_014_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_014_src_valid),                                                             //          .valid
		.src_data           (addr_router_014_src_data),                                                              //          .data
		.src_channel        (addr_router_014_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_014_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_014_src_endofpacket)                                                        //          .endofpacket
	);

	application_selector_id_router_013 id_router_013 (
		.sink_ready         (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_sdram_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sdram_1_phy_clk_out),                                                   //       clk.clk
		.reset              (~ddr2_sdram_1_reset_request_n_reset),                                        // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                    //       src.ready
		.src_valid          (id_router_013_src_valid),                                                    //          .valid
		.src_data           (id_router_013_src_data),                                                     //          .data
		.src_channel        (id_router_013_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                               //          .endofpacket
	);

	application_selector_addr_router_015 addr_router_015 (
		.sink_ready         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_015_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_015_src_valid),                                                             //          .valid
		.src_data           (addr_router_015_src_data),                                                              //          .data
		.src_channel        (addr_router_015_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_015_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_015_src_endofpacket)                                                        //          .endofpacket
	);

	application_selector_id_router_014 id_router_014 (
		.sink_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                  //       src.ready
		.src_valid          (id_router_014_src_valid),                                                  //          .valid
		.src_data           (id_router_014_src_data),                                                   //          .data
		.src_channel        (id_router_014_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                             //          .endofpacket
	);

	application_selector_id_router_014 id_router_015 (
		.sink_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                   //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                      //       src.ready
		.src_valid          (id_router_015_src_valid),                                                      //          .valid
		.src_data           (id_router_015_src_data),                                                       //          .data
		.src_channel        (id_router_015_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                 //          .endofpacket
	);

	application_selector_id_router_014 id_router_016 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                             //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                                //       src.ready
		.src_valid          (id_router_016_src_valid),                                                                //          .valid
		.src_data           (id_router_016_src_data),                                                                 //          .data
		.src_channel        (id_router_016_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                           //          .endofpacket
	);

	application_selector_id_router_014 id_router_017 (
		.sink_ready         (uart1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                          //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                             //       src.ready
		.src_valid          (id_router_017_src_valid),                                             //          .valid
		.src_data           (id_router_017_src_data),                                              //          .data
		.src_channel        (id_router_017_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                        //          .endofpacket
	);

	application_selector_id_router_014 id_router_018 (
		.sink_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                               //       src.ready
		.src_valid          (id_router_018_src_valid),                                               //          .valid
		.src_data           (id_router_018_src_data),                                                //          .data
		.src_channel        (id_router_018_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                          //          .endofpacket
	);

	application_selector_id_router_014 id_router_019 (
		.sink_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                                   //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_019_src_valid),                                                                      //          .valid
		.src_data           (id_router_019_src_data),                                                                       //          .data
		.src_channel        (id_router_019_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                                                 //          .endofpacket
	);

	application_selector_id_router_014 id_router_020 (
		.sink_ready         (pll_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pll_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pll_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pll_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pll_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                           //       src.ready
		.src_valid          (id_router_020_src_valid),                                           //          .valid
		.src_data           (id_router_020_src_data),                                            //          .data
		.src_channel        (id_router_020_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                      //          .endofpacket
	);

	application_selector_id_router_014 id_router_021 (
		.sink_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                  //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                     //       src.ready
		.src_valid          (id_router_021_src_valid),                                                     //          .valid
		.src_data           (id_router_021_src_data),                                                      //          .data
		.src_channel        (id_router_021_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                                //          .endofpacket
	);

	application_selector_id_router_014 id_router_022 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                     //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                                        //       src.ready
		.src_valid          (id_router_022_src_valid),                                                        //          .valid
		.src_data           (id_router_022_src_data),                                                         //          .data
		.src_channel        (id_router_022_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                                   //          .endofpacket
	);

	application_selector_id_router_014 id_router_023 (
		.sink_ready         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                                  //       src.ready
		.src_valid          (id_router_023_src_valid),                                                  //          .valid
		.src_data           (id_router_023_src_data),                                                   //          .data
		.src_channel        (id_router_023_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                             //          .endofpacket
	);

	application_selector_id_router_014 id_router_024 (
		.sink_ready         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                                   //       src.ready
		.src_valid          (id_router_024_src_valid),                                                   //          .valid
		.src_data           (id_router_024_src_data),                                                    //          .data
		.src_channel        (id_router_024_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                              //          .endofpacket
	);

	application_selector_id_router_014 id_router_025 (
		.sink_ready         (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_i2c_sdat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                 //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                    //       src.ready
		.src_valid          (id_router_025_src_valid),                                                    //          .valid
		.src_data           (id_router_025_src_data),                                                     //          .data
		.src_channel        (id_router_025_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                               //          .endofpacket
	);

	application_selector_id_router_014 id_router_026 (
		.sink_ready         (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_id_eeprom_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                      //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                                         //       src.ready
		.src_valid          (id_router_026_src_valid),                                                         //          .valid
		.src_data           (id_router_026_src_data),                                                          //          .data
		.src_channel        (id_router_026_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                                    //          .endofpacket
	);

	application_selector_id_router_014 id_router_027 (
		.sink_ready         (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_id_eeprom_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                      //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                                         //       src.ready
		.src_valid          (id_router_027_src_valid),                                                         //          .valid
		.src_data           (id_router_027_src_data),                                                          //          .data
		.src_channel        (id_router_027_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                                    //          .endofpacket
	);

	application_selector_id_router_014 id_router_028 (
		.sink_ready         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                          //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                                             //       src.ready
		.src_valid          (id_router_028_src_valid),                                                             //          .valid
		.src_data           (id_router_028_src_data),                                                              //          .data
		.src_channel        (id_router_028_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                                        //          .endofpacket
	);

	application_selector_id_router_014 id_router_029 (
		.sink_ready         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                                  //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_029_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_029_src_valid),                                                                     //          .valid
		.src_data           (id_router_029_src_data),                                                                      //          .data
		.src_channel        (id_router_029_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_029_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_029_src_endofpacket)                                                                //          .endofpacket
	);

	application_selector_addr_router_016 addr_router_016 (
		.sink_ready         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (addr_router_016_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_016_src_valid),                                                    //          .valid
		.src_data           (addr_router_016_src_data),                                                     //          .data
		.src_channel        (addr_router_016_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_016_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_016_src_endofpacket)                                               //          .endofpacket
	);

	application_selector_addr_router_016 addr_router_017 (
		.sink_ready         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_017_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_017_src_valid),                                                   //          .valid
		.src_data           (addr_router_017_src_data),                                                    //          .data
		.src_channel        (addr_router_017_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_017_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_017_src_endofpacket)                                              //          .endofpacket
	);

	application_selector_id_router_030 id_router_030 (
		.sink_ready         (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tse_ddr_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_030_src_ready),                                                            //       src.ready
		.src_valid          (id_router_030_src_valid),                                                            //          .valid
		.src_data           (id_router_030_src_data),                                                             //          .data
		.src_channel        (id_router_030_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_030_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_030_src_endofpacket)                                                       //          .endofpacket
	);

	application_selector_addr_router_018 addr_router_018 (
		.sink_ready         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pipeline_bridge_before_tristate_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                                    // clk_reset.reset
		.src_ready          (addr_router_018_src_ready),                                                                             //       src.ready
		.src_valid          (addr_router_018_src_valid),                                                                             //          .valid
		.src_data           (addr_router_018_src_data),                                                                              //          .data
		.src_channel        (addr_router_018_src_channel),                                                                           //          .channel
		.src_startofpacket  (addr_router_018_src_startofpacket),                                                                     //          .startofpacket
		.src_endofpacket    (addr_router_018_src_endofpacket)                                                                        //          .endofpacket
	);

	application_selector_id_router_031 id_router_031 (
		.sink_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_031_src_ready),                                                  //       src.ready
		.src_valid          (id_router_031_src_valid),                                                  //          .valid
		.src_data           (id_router_031_src_data),                                                   //          .data
		.src_channel        (id_router_031_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_031_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_031_src_endofpacket)                                             //          .endofpacket
	);

	application_selector_id_router_032 id_router_032 (
		.sink_ready         (max2_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (max2_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (max2_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (max2_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (max2_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_032_src_ready),                                             //       src.ready
		.src_valid          (id_router_032_src_valid),                                             //          .valid
		.src_data           (id_router_032_src_data),                                              //          .data
		.src_channel        (id_router_032_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_032_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_032_src_endofpacket)                                        //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (84),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.VALID_WIDTH               (10),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (pll_c0_out),                         //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),              //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),              //          .valid
		.cmd_sink_data          (addr_router_src_data),               //          .data
		.cmd_sink_channel       (addr_router_src_channel),            //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),             //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),             //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),           //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),              //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket),     //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),       //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (76),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.VALID_WIDTH               (10),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (pll_c0_out),                         //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.VALID_WIDTH               (10),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (pll_c0_out),                            //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.cmd_sink_ready         (addr_router_002_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_002_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_002_src_data),              //          .data
		.cmd_sink_channel       (addr_router_002_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_001_src1_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.VALID_WIDTH               (10),
		.ENFORCE_ORDER             (0),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_003 (
		.clk                    (pll_c0_out),                            //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_003_src_data),              //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_003_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_003_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_003_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_003_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_003_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_001_src2_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_003_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_003_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_003_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_003_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_003_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_003_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_003_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.VALID_WIDTH               (10),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_004 (
		.clk                    (pll_c0_out),                            //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.cmd_sink_ready         (addr_router_004_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_004_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_004_src_data),              //          .data
		.cmd_sink_channel       (addr_router_004_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_004_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_004_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_004_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_004_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_004_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_001_src3_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_004_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_004_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_004_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_004_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_004_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_004_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_004_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (10),
		.VALID_WIDTH               (10),
		.ENFORCE_ORDER             (0),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_005 (
		.clk                    (pll_c0_out),                            //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.cmd_sink_ready         (addr_router_005_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_005_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_005_src_data),              //          .data
		.cmd_sink_channel       (addr_router_005_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_005_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_005_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_005_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_005_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_005_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_001_src4_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_001_src4_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_001_src4_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_001_src4_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_005_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_005_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_005_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_005_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_005_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_005_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_005_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (36),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_006 (
		.clk                    (ddr2_sdram_phy_clk_out),              //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset),  // clk_reset.reset
		.cmd_sink_ready         (addr_router_006_src_ready),           //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_006_src_valid),           //          .valid
		.cmd_sink_data          (addr_router_006_src_data),            //          .data
		.cmd_sink_channel       (addr_router_006_src_channel),         //          .channel
		.cmd_sink_startofpacket (addr_router_006_src_startofpacket),   //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_006_src_endofpacket),     //          .endofpacket
		.cmd_src_ready          (limiter_006_cmd_src_ready),           //   cmd_src.ready
		.cmd_src_data           (limiter_006_cmd_src_data),            //          .data
		.cmd_src_channel        (limiter_006_cmd_src_channel),         //          .channel
		.cmd_src_startofpacket  (limiter_006_cmd_src_startofpacket),   //          .startofpacket
		.cmd_src_endofpacket    (limiter_006_cmd_src_endofpacket),     //          .endofpacket
		.rsp_sink_ready         (width_adapter_004_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (width_adapter_004_src_valid),         //          .valid
		.rsp_sink_channel       (width_adapter_004_src_channel),       //          .channel
		.rsp_sink_data          (width_adapter_004_src_data),          //          .data
		.rsp_sink_startofpacket (width_adapter_004_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (width_adapter_004_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_006_rsp_src_ready),           //   rsp_src.ready
		.rsp_src_valid          (limiter_006_rsp_src_valid),           //          .valid
		.rsp_src_data           (limiter_006_rsp_src_data),            //          .data
		.rsp_src_channel        (limiter_006_rsp_src_channel),         //          .channel
		.rsp_src_startofpacket  (limiter_006_rsp_src_startofpacket),   //          .startofpacket
		.rsp_src_endofpacket    (limiter_006_rsp_src_endofpacket),     //          .endofpacket
		.cmd_src_valid          (limiter_006_cmd_valid_data)           // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (36),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_007 (
		.clk                    (ddr2_sdram_phy_clk_out),              //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset),  // clk_reset.reset
		.cmd_sink_ready         (addr_router_007_src_ready),           //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_007_src_valid),           //          .valid
		.cmd_sink_data          (addr_router_007_src_data),            //          .data
		.cmd_sink_channel       (addr_router_007_src_channel),         //          .channel
		.cmd_sink_startofpacket (addr_router_007_src_startofpacket),   //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_007_src_endofpacket),     //          .endofpacket
		.cmd_src_ready          (limiter_007_cmd_src_ready),           //   cmd_src.ready
		.cmd_src_data           (limiter_007_cmd_src_data),            //          .data
		.cmd_src_channel        (limiter_007_cmd_src_channel),         //          .channel
		.cmd_src_startofpacket  (limiter_007_cmd_src_startofpacket),   //          .startofpacket
		.cmd_src_endofpacket    (limiter_007_cmd_src_endofpacket),     //          .endofpacket
		.rsp_sink_ready         (width_adapter_005_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (width_adapter_005_src_valid),         //          .valid
		.rsp_sink_channel       (width_adapter_005_src_channel),       //          .channel
		.rsp_sink_data          (width_adapter_005_src_data),          //          .data
		.rsp_sink_startofpacket (width_adapter_005_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (width_adapter_005_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_007_rsp_src_ready),           //   rsp_src.ready
		.rsp_src_valid          (limiter_007_rsp_src_valid),           //          .valid
		.rsp_src_data           (limiter_007_rsp_src_data),            //          .data
		.rsp_src_channel        (limiter_007_rsp_src_channel),         //          .channel
		.rsp_src_startofpacket  (limiter_007_rsp_src_startofpacket),   //          .startofpacket
		.rsp_src_endofpacket    (limiter_007_rsp_src_endofpacket),     //          .endofpacket
		.cmd_src_valid          (limiter_007_cmd_valid_data)           // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (123),
		.PKT_DEST_ID_L             (121),
		.PKT_TRANS_POSTED          (105),
		.MAX_OUTSTANDING_RESPONSES (36),
		.PIPELINED                 (0),
		.ST_DATA_W                 (125),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (112),
		.PKT_BYTE_CNT_L            (109),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64)
	) limiter_008 (
		.clk                    (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.cmd_sink_ready         (addr_router_008_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_008_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_008_src_data),              //          .data
		.cmd_sink_channel       (addr_router_008_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_008_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_008_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_008_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_008_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_008_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_008_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_008_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_010_src2_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_010_src2_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_010_src2_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_010_src2_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_010_src2_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_010_src2_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_008_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_008_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_008_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_008_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_008_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_008_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_008_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (123),
		.PKT_DEST_ID_L             (121),
		.PKT_TRANS_POSTED          (105),
		.MAX_OUTSTANDING_RESPONSES (36),
		.PIPELINED                 (0),
		.ST_DATA_W                 (125),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (112),
		.PKT_BYTE_CNT_L            (109),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64)
	) limiter_009 (
		.clk                    (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.cmd_sink_ready         (addr_router_009_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_009_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_009_src_data),              //          .data
		.cmd_sink_channel       (addr_router_009_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_009_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_009_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_009_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_009_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_009_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_009_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_009_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_010_src3_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_010_src3_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_010_src3_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_010_src3_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_010_src3_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_010_src3_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_009_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_009_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_009_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_009_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_009_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_009_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_009_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (36),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_010 (
		.clk                    (ddr2_sdram_phy_clk_out),             //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_010_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_010_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_010_src_data),           //          .data
		.cmd_sink_channel       (addr_router_010_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_010_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_010_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_010_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_010_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_010_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_010_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_010_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_010_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_010_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_010_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_010_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_010_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_010_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_010_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_010_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_010_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_010_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_010_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_010_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_010_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (36),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_011 (
		.clk                    (ddr2_sdram_phy_clk_out),              //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset),  // clk_reset.reset
		.cmd_sink_ready         (addr_router_011_src_ready),           //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_011_src_valid),           //          .valid
		.cmd_sink_data          (addr_router_011_src_data),            //          .data
		.cmd_sink_channel       (addr_router_011_src_channel),         //          .channel
		.cmd_sink_startofpacket (addr_router_011_src_startofpacket),   //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_011_src_endofpacket),     //          .endofpacket
		.cmd_src_ready          (limiter_011_cmd_src_ready),           //   cmd_src.ready
		.cmd_src_data           (limiter_011_cmd_src_data),            //          .data
		.cmd_src_channel        (limiter_011_cmd_src_channel),         //          .channel
		.cmd_src_startofpacket  (limiter_011_cmd_src_startofpacket),   //          .startofpacket
		.cmd_src_endofpacket    (limiter_011_cmd_src_endofpacket),     //          .endofpacket
		.rsp_sink_ready         (width_adapter_007_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (width_adapter_007_src_valid),         //          .valid
		.rsp_sink_channel       (width_adapter_007_src_channel),       //          .channel
		.rsp_sink_data          (width_adapter_007_src_data),          //          .data
		.rsp_sink_startofpacket (width_adapter_007_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (width_adapter_007_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_011_rsp_src_ready),           //   rsp_src.ready
		.rsp_src_valid          (limiter_011_rsp_src_valid),           //          .valid
		.rsp_src_data           (limiter_011_rsp_src_data),            //          .data
		.rsp_src_channel        (limiter_011_rsp_src_channel),         //          .channel
		.rsp_src_startofpacket  (limiter_011_rsp_src_startofpacket),   //          .startofpacket
		.rsp_src_endofpacket    (limiter_011_rsp_src_endofpacket),     //          .endofpacket
		.cmd_src_valid          (limiter_011_cmd_valid_data)           // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (63),
		.PKT_TRANS_POSTED          (47),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (69),
		.ST_CHANNEL_W              (16),
		.VALID_WIDTH               (16),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_012 (
		.clk                    (pll_c2_out),                         //       clk.clk
		.reset                  (rst_controller_004_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_015_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_015_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_015_src_data),           //          .data
		.cmd_sink_channel       (addr_router_015_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_015_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_015_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_012_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_012_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_012_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_012_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_012_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_015_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_015_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_015_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_015_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_015_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_015_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_012_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_012_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_012_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_012_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_012_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_012_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_012_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (77),
		.PKT_TRANS_POSTED          (64),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (2),
		.VALID_WIDTH               (2),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_013 (
		.clk                    (pll_c0_out),                         //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_018_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_018_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_018_src_data),           //          .data
		.cmd_sink_channel       (addr_router_018_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_018_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_018_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_013_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_013_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_013_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_013_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_013_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_018_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_018_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_018_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_018_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_018_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_018_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_013_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_013_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_013_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_013_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_013_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_013_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_013_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (56),
		.PKT_BYTE_CNT_H            (52),
		.PKT_BYTE_CNT_L            (50),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (53),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.ST_DATA_W                 (62),
		.ST_CHANNEL_W              (2),
		.OUT_BYTE_CNT_H            (51),
		.OUT_BURSTWRAP_H           (55),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter (
		.clk                   (pll_c0_out),                          //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_010_src_valid),         //     sink0.valid
		.sink0_data            (width_adapter_010_src_data),          //          .data
		.sink0_channel         (width_adapter_010_src_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_010_src_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_010_src_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_010_src_ready),         //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (6),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_n),                            // reset_in0.reset
		.reset_in1  (~reset_n),                            // reset_in1.reset
		.reset_in2  (pll_resetrequest_reset),              // reset_in2.reset
		.reset_in3  (~ddr2_sdram_reset_request_n_reset),   // reset_in3.reset
		.reset_in4  (~ddr2_sdram_1_reset_request_n_reset), // reset_in4.reset
		.reset_in5  (cpu_jtag_debug_module_reset_reset),   // reset_in5.reset
		.clk        (clk),                                 //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (6),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_n),                            // reset_in0.reset
		.reset_in1  (~reset_n),                            // reset_in1.reset
		.reset_in2  (pll_resetrequest_reset),              // reset_in2.reset
		.reset_in3  (~ddr2_sdram_reset_request_n_reset),   // reset_in3.reset
		.reset_in4  (~ddr2_sdram_1_reset_request_n_reset), // reset_in4.reset
		.reset_in5  (cpu_jtag_debug_module_reset_reset),   // reset_in5.reset
		.clk        (pll_c0_out),                          //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (6),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_n),                            // reset_in0.reset
		.reset_in1  (~reset_n),                            // reset_in1.reset
		.reset_in2  (pll_resetrequest_reset),              // reset_in2.reset
		.reset_in3  (~ddr2_sdram_reset_request_n_reset),   // reset_in3.reset
		.reset_in4  (~ddr2_sdram_1_reset_request_n_reset), // reset_in4.reset
		.reset_in5  (cpu_jtag_debug_module_reset_reset),   // reset_in5.reset
		.clk        (clk_125),                             //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),  // reset_out.reset
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (6),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_n),                            // reset_in0.reset
		.reset_in1  (~reset_n),                            // reset_in1.reset
		.reset_in2  (pll_resetrequest_reset),              // reset_in2.reset
		.reset_in3  (~ddr2_sdram_reset_request_n_reset),   // reset_in3.reset
		.reset_in4  (~ddr2_sdram_1_reset_request_n_reset), // reset_in4.reset
		.reset_in5  (cpu_jtag_debug_module_reset_reset),   // reset_in5.reset
		.clk        (ddr2_sdram_phy_clk_out),              //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset),  // reset_out.reset
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (6),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_004 (
		.reset_in0  (~reset_n),                            // reset_in0.reset
		.reset_in1  (~reset_n),                            // reset_in1.reset
		.reset_in2  (pll_resetrequest_reset),              // reset_in2.reset
		.reset_in3  (~ddr2_sdram_reset_request_n_reset),   // reset_in3.reset
		.reset_in4  (~ddr2_sdram_1_reset_request_n_reset), // reset_in4.reset
		.reset_in5  (cpu_jtag_debug_module_reset_reset),   // reset_in5.reset
		.clk        (pll_c2_out),                          //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset),  // reset_out.reset
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (6),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_005 (
		.reset_in0  (~reset_n),                            // reset_in0.reset
		.reset_in1  (~reset_n),                            // reset_in1.reset
		.reset_in2  (pll_resetrequest_reset),              // reset_in2.reset
		.reset_in3  (~ddr2_sdram_reset_request_n_reset),   // reset_in3.reset
		.reset_in4  (~ddr2_sdram_1_reset_request_n_reset), // reset_in4.reset
		.reset_in5  (cpu_jtag_debug_module_reset_reset),   // reset_in5.reset
		.clk        (ddr2_sdram_1_phy_clk_out),            //       clk.clk
		.reset_out  (rst_controller_005_reset_out_reset),  // reset_out.reset
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	application_selector_cmd_xbar_demux cmd_xbar_demux (
		.clk                (pll_c0_out),                         //        clk.clk
		.reset              (rst_controller_001_reset_out_reset), //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),            //           .channel
		.sink_data          (limiter_cmd_src_data),               //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),    //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),          //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),          //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),           //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),        //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket),    //           .endofpacket
		.src5_ready         (cmd_xbar_demux_src5_ready),          //       src5.ready
		.src5_valid         (cmd_xbar_demux_src5_valid),          //           .valid
		.src5_data          (cmd_xbar_demux_src5_data),           //           .data
		.src5_channel       (cmd_xbar_demux_src5_channel),        //           .channel
		.src5_startofpacket (cmd_xbar_demux_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_src5_endofpacket),    //           .endofpacket
		.src6_ready         (cmd_xbar_demux_src6_ready),          //       src6.ready
		.src6_valid         (cmd_xbar_demux_src6_valid),          //           .valid
		.src6_data          (cmd_xbar_demux_src6_data),           //           .data
		.src6_channel       (cmd_xbar_demux_src6_channel),        //           .channel
		.src6_startofpacket (cmd_xbar_demux_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_src6_endofpacket),    //           .endofpacket
		.src7_ready         (cmd_xbar_demux_src7_ready),          //       src7.ready
		.src7_valid         (cmd_xbar_demux_src7_valid),          //           .valid
		.src7_data          (cmd_xbar_demux_src7_data),           //           .data
		.src7_channel       (cmd_xbar_demux_src7_channel),        //           .channel
		.src7_startofpacket (cmd_xbar_demux_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_src7_endofpacket),    //           .endofpacket
		.src8_ready         (cmd_xbar_demux_src8_ready),          //       src8.ready
		.src8_valid         (cmd_xbar_demux_src8_valid),          //           .valid
		.src8_data          (cmd_xbar_demux_src8_data),           //           .data
		.src8_channel       (cmd_xbar_demux_src8_channel),        //           .channel
		.src8_startofpacket (cmd_xbar_demux_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_src8_endofpacket),    //           .endofpacket
		.src9_ready         (cmd_xbar_demux_src9_ready),          //       src9.ready
		.src9_valid         (cmd_xbar_demux_src9_valid),          //           .valid
		.src9_data          (cmd_xbar_demux_src9_data),           //           .data
		.src9_channel       (cmd_xbar_demux_src9_channel),        //           .channel
		.src9_startofpacket (cmd_xbar_demux_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket   (cmd_xbar_demux_src9_endofpacket)     //           .endofpacket
	);

	application_selector_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_002_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_002_cmd_src_channel),           //           .channel
		.sink_data          (limiter_002_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_002_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_002_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_002_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_003_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_003_cmd_src_channel),           //           .channel
		.sink_data          (limiter_003_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_003_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_003_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_003_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_demux_002 cmd_xbar_demux_004 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_004_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_004_cmd_src_channel),           //           .channel
		.sink_data          (limiter_004_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_004_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_004_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_004_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_demux_002 cmd_xbar_demux_005 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_005_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_005_cmd_src_channel),           //           .channel
		.sink_data          (limiter_005_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_005_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_005_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_005_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_004_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (cmd_xbar_demux_005_src0_ready),         //     sink4.ready
		.sink4_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.sink4_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.sink4_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.sink4_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_mux_006 cmd_xbar_mux_006 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src6_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src6_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src6_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src6_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src6_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src6_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_mux_006 cmd_xbar_mux_008 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src8_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src8_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src8_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src8_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src8_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src8_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux rsp_xbar_demux (
		.clk                (pll_c0_out),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	application_selector_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (rsp_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (rsp_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (rsp_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (rsp_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (rsp_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (rsp_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (crosser_001_out_ready),                 //     sink5.ready
		.sink5_valid         (crosser_001_out_valid),                 //          .valid
		.sink5_channel       (crosser_001_out_channel),               //          .channel
		.sink5_data          (crosser_001_out_data),                  //          .data
		.sink5_startofpacket (crosser_001_out_startofpacket),         //          .startofpacket
		.sink5_endofpacket   (crosser_001_out_endofpacket),           //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready         (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_006_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_008_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_demux_006 cmd_xbar_demux_006 (
		.clk                (ddr2_sdram_phy_clk_out),                //        clk.clk
		.reset              (rst_controller_003_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_006_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_006_cmd_src_channel),           //           .channel
		.sink_data          (limiter_006_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_006_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_006_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_006_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_006_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_006_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_006_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_006_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_006_src0_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_demux_006 cmd_xbar_demux_007 (
		.clk                (ddr2_sdram_phy_clk_out),                //        clk.clk
		.reset              (rst_controller_003_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_007_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_007_cmd_src_channel),           //           .channel
		.sink_data          (limiter_007_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_007_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_007_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_007_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_007_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_007_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_007_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_007_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_007_src0_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_demux_008 cmd_xbar_demux_008 (
		.clk                (ddr2_sdram_phy_clk_out),                //        clk.clk
		.reset              (rst_controller_003_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_008_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_008_cmd_src_channel),           //           .channel
		.sink_data          (limiter_008_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_008_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_008_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_008_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_008_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_008_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_008_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_008_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_008_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_008_src0_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_demux_008 cmd_xbar_demux_009 (
		.clk                (ddr2_sdram_phy_clk_out),                //        clk.clk
		.reset              (rst_controller_003_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_009_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_009_cmd_src_channel),           //           .channel
		.sink_data          (limiter_009_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_009_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_009_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_009_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_009_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_009_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_009_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_009_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_009_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_009_src0_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_demux_010 cmd_xbar_demux_010 (
		.clk                (ddr2_sdram_phy_clk_out),                //        clk.clk
		.reset              (rst_controller_003_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_010_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_010_cmd_src_channel),           //           .channel
		.sink_data          (limiter_010_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_010_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_010_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_010_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_010_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_010_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_010_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_010_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_010_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_010_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_010_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_010_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_010_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_010_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_010_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_010_src1_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_demux_006 cmd_xbar_demux_011 (
		.clk                (ddr2_sdram_phy_clk_out),                //        clk.clk
		.reset              (rst_controller_003_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_011_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_011_cmd_src_channel),           //           .channel
		.sink_data          (limiter_011_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_011_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_011_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_011_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_011_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_011_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_011_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_011_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_011_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_011_src0_endofpacket)    //           .endofpacket
	);

	application_selector_cmd_xbar_mux_010 cmd_xbar_mux_010 (
		.clk                 (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset               (~ddr2_sdram_reset_request_n_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_src_ready),               //     sink0.ready
		.sink0_valid         (width_adapter_src_valid),               //          .valid
		.sink0_channel       (width_adapter_src_channel),             //          .channel
		.sink0_data          (width_adapter_src_data),                //          .data
		.sink0_startofpacket (width_adapter_src_startofpacket),       //          .startofpacket
		.sink0_endofpacket   (width_adapter_src_endofpacket),         //          .endofpacket
		.sink1_ready         (width_adapter_001_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_001_src_valid),           //          .valid
		.sink1_channel       (width_adapter_001_src_channel),         //          .channel
		.sink1_data          (width_adapter_001_src_data),            //          .data
		.sink1_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_008_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_008_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_008_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_008_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_009_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_009_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_009_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_009_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (width_adapter_002_src_ready),           //     sink4.ready
		.sink4_valid         (width_adapter_002_src_valid),           //          .valid
		.sink4_channel       (width_adapter_002_src_channel),         //          .channel
		.sink4_data          (width_adapter_002_src_data),            //          .data
		.sink4_startofpacket (width_adapter_002_src_startofpacket),   //          .startofpacket
		.sink4_endofpacket   (width_adapter_002_src_endofpacket),     //          .endofpacket
		.sink5_ready         (width_adapter_003_src_ready),           //     sink5.ready
		.sink5_valid         (width_adapter_003_src_valid),           //          .valid
		.sink5_channel       (width_adapter_003_src_channel),         //          .channel
		.sink5_data          (width_adapter_003_src_data),            //          .data
		.sink5_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink5_endofpacket   (width_adapter_003_src_endofpacket)      //          .endofpacket
	);

	application_selector_rsp_xbar_demux_010 rsp_xbar_demux_010 (
		.clk                (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset              (~ddr2_sdram_reset_request_n_reset),     // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_010_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_010_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_010_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_010_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_010_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_010_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_010_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_010_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_010_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_010_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_010_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_010_src3_endofpacket),   //          .endofpacket
		.src4_ready         (rsp_xbar_demux_010_src4_ready),         //      src4.ready
		.src4_valid         (rsp_xbar_demux_010_src4_valid),         //          .valid
		.src4_data          (rsp_xbar_demux_010_src4_data),          //          .data
		.src4_channel       (rsp_xbar_demux_010_src4_channel),       //          .channel
		.src4_startofpacket (rsp_xbar_demux_010_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (rsp_xbar_demux_010_src4_endofpacket),   //          .endofpacket
		.src5_ready         (rsp_xbar_demux_010_src5_ready),         //      src5.ready
		.src5_valid         (rsp_xbar_demux_010_src5_valid),         //          .valid
		.src5_data          (rsp_xbar_demux_010_src5_data),          //          .data
		.src5_channel       (rsp_xbar_demux_010_src5_channel),       //          .channel
		.src5_startofpacket (rsp_xbar_demux_010_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (rsp_xbar_demux_010_src5_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_011 rsp_xbar_demux_011 (
		.clk                (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_mux_010 rsp_xbar_mux_010 (
		.clk                 (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_010_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_010_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_010_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_010_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_010_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_010_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_006_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_006_src_valid),           //          .valid
		.sink0_channel       (width_adapter_006_src_channel),         //          .channel
		.sink0_data          (width_adapter_006_src_data),            //          .data
		.sink0_startofpacket (width_adapter_006_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_006_src_endofpacket),     //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_011_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_demux_012 cmd_xbar_demux_012 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_012_src_ready),             //      sink.ready
		.sink_channel       (addr_router_012_src_channel),           //          .channel
		.sink_data          (addr_router_012_src_data),              //          .data
		.sink_startofpacket (addr_router_012_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_012_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_012_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_demux_012 cmd_xbar_demux_013 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_013_src_ready),             //      sink.ready
		.sink_channel       (addr_router_013_src_channel),           //          .channel
		.sink_data          (addr_router_013_src_data),              //          .data
		.sink_startofpacket (addr_router_013_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_013_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_013_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_mux_012 cmd_xbar_mux_012 (
		.clk                 (pll_c0_out),                         //       clk.clk
		.reset               (rst_controller_001_reset_out_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_012_src_ready),         //       src.ready
		.src_valid           (cmd_xbar_mux_012_src_valid),         //          .valid
		.src_data            (cmd_xbar_mux_012_src_data),          //          .data
		.src_channel         (cmd_xbar_mux_012_src_channel),       //          .channel
		.src_startofpacket   (cmd_xbar_mux_012_src_startofpacket), //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_012_src_endofpacket),   //          .endofpacket
		.sink0_ready         (crosser_002_out_ready),              //     sink0.ready
		.sink0_valid         (crosser_002_out_valid),              //          .valid
		.sink0_channel       (crosser_002_out_channel),            //          .channel
		.sink0_data          (crosser_002_out_data),               //          .data
		.sink0_startofpacket (crosser_002_out_startofpacket),      //          .startofpacket
		.sink0_endofpacket   (crosser_002_out_endofpacket),        //          .endofpacket
		.sink1_ready         (crosser_003_out_ready),              //     sink1.ready
		.sink1_valid         (crosser_003_out_valid),              //          .valid
		.sink1_channel       (crosser_003_out_channel),            //          .channel
		.sink1_data          (crosser_003_out_data),               //          .data
		.sink1_startofpacket (crosser_003_out_startofpacket),      //          .startofpacket
		.sink1_endofpacket   (crosser_003_out_endofpacket)         //          .endofpacket
	);

	application_selector_rsp_xbar_demux_012 rsp_xbar_demux_012 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_009_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_009_src_channel),         //          .channel
		.sink_data          (width_adapter_009_src_data),            //          .data
		.sink_startofpacket (width_adapter_009_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_009_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_009_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_012_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_012_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_012_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_012_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_012_src1_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_demux_014 cmd_xbar_demux_014 (
		.clk                (ddr2_sdram_1_phy_clk_out),              //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_014_src_ready),             //      sink.ready
		.sink_channel       (addr_router_014_src_channel),           //          .channel
		.sink_data          (addr_router_014_src_data),              //          .data
		.sink_startofpacket (addr_router_014_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_014_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_014_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_demux_014 rsp_xbar_demux_013 (
		.clk                (ddr2_sdram_1_phy_clk_out),              //       clk.clk
		.reset              (~ddr2_sdram_1_reset_request_n_reset),   // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_demux_015 cmd_xbar_demux_015 (
		.clk                 (pll_c2_out),                             //        clk.clk
		.reset               (rst_controller_004_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_012_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_012_cmd_src_channel),            //           .channel
		.sink_data           (limiter_012_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_012_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_012_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_012_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_015_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_015_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_015_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_015_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_015_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_015_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_015_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_015_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_015_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_015_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_015_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_015_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_015_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_015_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_015_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_015_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_015_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_015_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_015_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_015_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_015_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_015_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_015_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_015_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_015_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_015_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_015_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_015_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_015_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_015_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_015_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_015_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_015_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_015_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_015_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_015_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_015_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_015_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_015_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_015_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_015_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_015_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_015_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_015_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_015_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_015_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_015_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_015_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_015_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_015_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_015_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_015_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_015_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_015_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_015_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_015_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_015_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_015_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_015_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_015_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_015_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_015_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_015_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_015_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_015_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_015_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_015_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_015_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_015_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_015_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_015_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_015_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_015_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_015_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_015_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_015_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_015_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_015_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_015_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_015_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_015_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_015_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_015_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_015_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_015_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_015_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_015_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_015_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_015_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_015_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_015_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_015_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_015_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_015_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_015_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_015_src15_endofpacket)    //           .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_014 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_015 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_016 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_017 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_018 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_019 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_020 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_021 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_022 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_023 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_024 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_025 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_026 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_026_src_ready),               //      sink.ready
		.sink_channel       (id_router_026_src_channel),             //          .channel
		.sink_data          (id_router_026_src_data),                //          .data
		.sink_startofpacket (id_router_026_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_026_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_026_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_027 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_027_src_ready),               //      sink.ready
		.sink_channel       (id_router_027_src_channel),             //          .channel
		.sink_data          (id_router_027_src_data),                //          .data
		.sink_startofpacket (id_router_027_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_027_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_027_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_028 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_028_src_ready),               //      sink.ready
		.sink_channel       (id_router_028_src_channel),             //          .channel
		.sink_data          (id_router_028_src_data),                //          .data
		.sink_startofpacket (id_router_028_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_028_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_028_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_014 rsp_xbar_demux_029 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_029_src_ready),               //      sink.ready
		.sink_channel       (id_router_029_src_channel),             //          .channel
		.sink_data          (id_router_029_src_data),                //          .data
		.sink_startofpacket (id_router_029_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_029_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_029_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_029_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_mux_015 rsp_xbar_mux_015 (
		.clk                  (pll_c2_out),                            //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_015_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_015_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_015_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_015_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_015_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_015_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_014_src0_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_014_src0_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_015_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_015_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_016_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_016_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_017_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_017_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_018_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_018_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_019_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_019_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (crosser_007_out_ready),                 //     sink6.ready
		.sink6_valid          (crosser_007_out_valid),                 //          .valid
		.sink6_channel        (crosser_007_out_channel),               //          .channel
		.sink6_data           (crosser_007_out_data),                  //          .data
		.sink6_startofpacket  (crosser_007_out_startofpacket),         //          .startofpacket
		.sink6_endofpacket    (crosser_007_out_endofpacket),           //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_021_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_021_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_022_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_022_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_023_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_023_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_024_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_025_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_026_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_027_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_028_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_028_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_029_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_demux_016 cmd_xbar_demux_016 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_016_src_ready),             //      sink.ready
		.sink_channel       (addr_router_016_src_channel),           //          .channel
		.sink_data          (addr_router_016_src_data),              //          .data
		.sink_startofpacket (addr_router_016_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_016_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_016_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_demux_016 cmd_xbar_demux_017 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_017_src_ready),             //      sink.ready
		.sink_channel       (addr_router_017_src_channel),           //          .channel
		.sink_data          (addr_router_017_src_data),              //          .data
		.sink_startofpacket (addr_router_017_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_017_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_017_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_mux_030 cmd_xbar_mux_030 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_030_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_030_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_030_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_030_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_030_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_030_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_016_src0_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_016_src0_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_016_src0_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_016_src0_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_017_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_017_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_017_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_017_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_030 rsp_xbar_demux_030 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_030_src_ready),               //      sink.ready
		.sink_channel       (id_router_030_src_channel),             //          .channel
		.sink_data          (id_router_030_src_data),                //          .data
		.sink_startofpacket (id_router_030_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_030_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_030_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_030_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_030_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_030_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_030_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_030_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_030_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_030_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_030_src1_endofpacket)    //          .endofpacket
	);

	application_selector_cmd_xbar_demux_018 cmd_xbar_demux_018 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_013_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_013_cmd_src_channel),           //           .channel
		.sink_data          (limiter_013_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_013_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_013_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_013_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_018_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_018_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_018_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_018_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_018_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_018_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_018_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_018_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_018_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_018_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_018_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_018_src1_endofpacket)    //           .endofpacket
	);

	application_selector_rsp_xbar_demux_031 rsp_xbar_demux_031 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_011_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_011_src_channel),         //          .channel
		.sink_data          (width_adapter_011_src_data),            //          .data
		.sink_startofpacket (width_adapter_011_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_011_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_011_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_031_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_031_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_demux_031 rsp_xbar_demux_032 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_032_src_ready),               //      sink.ready
		.sink_channel       (id_router_032_src_channel),             //          .channel
		.sink_data          (id_router_032_src_data),                //          .data
		.sink_startofpacket (id_router_032_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_032_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_032_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_032_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_032_src0_endofpacket)    //          .endofpacket
	);

	application_selector_rsp_xbar_mux_018 rsp_xbar_mux_018 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_018_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_018_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_018_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_018_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_018_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_018_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_031_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_031_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_032_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_032_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (80),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (112),
		.OUT_PKT_BYTE_CNT_L            (109),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_ST_DATA_W                 (125),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk               (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.in_valid          (cmd_xbar_demux_006_src0_valid),         //      sink.valid
		.in_channel        (cmd_xbar_demux_006_src0_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_demux_006_src0_ready),         //          .ready
		.in_data           (cmd_xbar_demux_006_src0_data),          //          .data
		.out_endofpacket   (width_adapter_src_endofpacket),         //       src.endofpacket
		.out_data          (width_adapter_src_data),                //          .data
		.out_channel       (width_adapter_src_channel),             //          .channel
		.out_valid         (width_adapter_src_valid),               //          .valid
		.out_ready         (width_adapter_src_ready),               //          .ready
		.out_startofpacket (width_adapter_src_startofpacket)        //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (80),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (112),
		.OUT_PKT_BYTE_CNT_L            (109),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_ST_DATA_W                 (125),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_001 (
		.clk               (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.in_valid          (cmd_xbar_demux_007_src0_valid),         //      sink.valid
		.in_channel        (cmd_xbar_demux_007_src0_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_demux_007_src0_ready),         //          .ready
		.in_data           (cmd_xbar_demux_007_src0_data),          //          .data
		.out_endofpacket   (width_adapter_001_src_endofpacket),     //       src.endofpacket
		.out_data          (width_adapter_001_src_data),            //          .data
		.out_channel       (width_adapter_001_src_channel),         //          .channel
		.out_valid         (width_adapter_001_src_valid),           //          .valid
		.out_ready         (width_adapter_001_src_ready),           //          .ready
		.out_startofpacket (width_adapter_001_src_startofpacket)    //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (80),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (112),
		.OUT_PKT_BYTE_CNT_L            (109),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_ST_DATA_W                 (125),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk               (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.in_valid          (cmd_xbar_demux_010_src0_valid),         //      sink.valid
		.in_channel        (cmd_xbar_demux_010_src0_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_demux_010_src0_ready),         //          .ready
		.in_data           (cmd_xbar_demux_010_src0_data),          //          .data
		.out_endofpacket   (width_adapter_002_src_endofpacket),     //       src.endofpacket
		.out_data          (width_adapter_002_src_data),            //          .data
		.out_channel       (width_adapter_002_src_channel),         //          .channel
		.out_valid         (width_adapter_002_src_valid),           //          .valid
		.out_ready         (width_adapter_002_src_ready),           //          .ready
		.out_startofpacket (width_adapter_002_src_startofpacket)    //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (80),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (112),
		.OUT_PKT_BYTE_CNT_L            (109),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_ST_DATA_W                 (125),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_003 (
		.clk               (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.in_valid          (cmd_xbar_demux_011_src0_valid),         //      sink.valid
		.in_channel        (cmd_xbar_demux_011_src0_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_demux_011_src0_ready),         //          .ready
		.in_data           (cmd_xbar_demux_011_src0_data),          //          .data
		.out_endofpacket   (width_adapter_003_src_endofpacket),     //       src.endofpacket
		.out_data          (width_adapter_003_src_data),            //          .data
		.out_channel       (width_adapter_003_src_channel),         //          .channel
		.out_valid         (width_adapter_003_src_valid),           //          .valid
		.out_ready         (width_adapter_003_src_ready),           //          .ready
		.out_startofpacket (width_adapter_003_src_startofpacket)    //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (112),
		.IN_PKT_BYTE_CNT_L             (109),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (116),
		.IN_PKT_BURSTWRAP_L            (113),
		.IN_ST_DATA_W                  (125),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_004 (
		.clk               (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset             (~ddr2_sdram_reset_request_n_reset),     // clk_reset.reset
		.in_valid          (rsp_xbar_demux_010_src0_valid),         //      sink.valid
		.in_channel        (rsp_xbar_demux_010_src0_channel),       //          .channel
		.in_startofpacket  (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.in_ready          (rsp_xbar_demux_010_src0_ready),         //          .ready
		.in_data           (rsp_xbar_demux_010_src0_data),          //          .data
		.out_endofpacket   (width_adapter_004_src_endofpacket),     //       src.endofpacket
		.out_data          (width_adapter_004_src_data),            //          .data
		.out_channel       (width_adapter_004_src_channel),         //          .channel
		.out_valid         (width_adapter_004_src_valid),           //          .valid
		.out_ready         (width_adapter_004_src_ready),           //          .ready
		.out_startofpacket (width_adapter_004_src_startofpacket)    //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (112),
		.IN_PKT_BYTE_CNT_L             (109),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (116),
		.IN_PKT_BURSTWRAP_L            (113),
		.IN_ST_DATA_W                  (125),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_005 (
		.clk               (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset             (~ddr2_sdram_reset_request_n_reset),     // clk_reset.reset
		.in_valid          (rsp_xbar_demux_010_src1_valid),         //      sink.valid
		.in_channel        (rsp_xbar_demux_010_src1_channel),       //          .channel
		.in_startofpacket  (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.in_ready          (rsp_xbar_demux_010_src1_ready),         //          .ready
		.in_data           (rsp_xbar_demux_010_src1_data),          //          .data
		.out_endofpacket   (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data          (width_adapter_005_src_data),            //          .data
		.out_channel       (width_adapter_005_src_channel),         //          .channel
		.out_valid         (width_adapter_005_src_valid),           //          .valid
		.out_ready         (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket (width_adapter_005_src_startofpacket)    //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (112),
		.IN_PKT_BYTE_CNT_L             (109),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (116),
		.IN_PKT_BURSTWRAP_L            (113),
		.IN_ST_DATA_W                  (125),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_006 (
		.clk               (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset             (~ddr2_sdram_reset_request_n_reset),     // clk_reset.reset
		.in_valid          (rsp_xbar_demux_010_src4_valid),         //      sink.valid
		.in_channel        (rsp_xbar_demux_010_src4_channel),       //          .channel
		.in_startofpacket  (rsp_xbar_demux_010_src4_startofpacket), //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_010_src4_endofpacket),   //          .endofpacket
		.in_ready          (rsp_xbar_demux_010_src4_ready),         //          .ready
		.in_data           (rsp_xbar_demux_010_src4_data),          //          .data
		.out_endofpacket   (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data          (width_adapter_006_src_data),            //          .data
		.out_channel       (width_adapter_006_src_channel),         //          .channel
		.out_valid         (width_adapter_006_src_valid),           //          .valid
		.out_ready         (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket (width_adapter_006_src_startofpacket)    //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (112),
		.IN_PKT_BYTE_CNT_L             (109),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (116),
		.IN_PKT_BURSTWRAP_L            (113),
		.IN_ST_DATA_W                  (125),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_007 (
		.clk               (ddr2_sdram_phy_clk_out),                //       clk.clk
		.reset             (~ddr2_sdram_reset_request_n_reset),     // clk_reset.reset
		.in_valid          (rsp_xbar_demux_010_src5_valid),         //      sink.valid
		.in_channel        (rsp_xbar_demux_010_src5_channel),       //          .channel
		.in_startofpacket  (rsp_xbar_demux_010_src5_startofpacket), //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_010_src5_endofpacket),   //          .endofpacket
		.in_ready          (rsp_xbar_demux_010_src5_ready),         //          .ready
		.in_data           (rsp_xbar_demux_010_src5_data),          //          .data
		.out_endofpacket   (width_adapter_007_src_endofpacket),     //       src.endofpacket
		.out_data          (width_adapter_007_src_data),            //          .data
		.out_channel       (width_adapter_007_src_channel),         //          .channel
		.out_valid         (width_adapter_007_src_valid),           //          .valid
		.out_ready         (width_adapter_007_src_ready),           //          .ready
		.out_startofpacket (width_adapter_007_src_startofpacket)    //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (80),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_ST_DATA_W                  (87),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (112),
		.OUT_PKT_BYTE_CNT_L            (109),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_ST_DATA_W                 (123),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_008 (
		.clk               (pll_c0_out),                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid          (cmd_xbar_mux_012_src_valid),          //      sink.valid
		.in_channel        (cmd_xbar_mux_012_src_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_mux_012_src_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_012_src_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_mux_012_src_ready),          //          .ready
		.in_data           (cmd_xbar_mux_012_src_data),           //          .data
		.out_endofpacket   (width_adapter_008_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_008_src_data),          //          .data
		.out_channel       (width_adapter_008_src_channel),       //          .channel
		.out_valid         (width_adapter_008_src_valid),         //          .valid
		.out_ready         (width_adapter_008_src_ready),         //          .ready
		.out_startofpacket (width_adapter_008_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (112),
		.IN_PKT_BYTE_CNT_L             (109),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (116),
		.IN_PKT_BURSTWRAP_L            (113),
		.IN_ST_DATA_W                  (123),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (87),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_009 (
		.clk               (pll_c0_out),                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid          (id_router_012_src_valid),             //      sink.valid
		.in_channel        (id_router_012_src_channel),           //          .channel
		.in_startofpacket  (id_router_012_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_012_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_012_src_ready),             //          .ready
		.in_data           (id_router_012_src_data),              //          .data
		.out_endofpacket   (width_adapter_009_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_009_src_data),          //          .data
		.out_channel       (width_adapter_009_src_channel),       //          .channel
		.out_valid         (width_adapter_009_src_valid),         //          .valid
		.out_ready         (width_adapter_009_src_ready),         //          .ready
		.out_startofpacket (width_adapter_009_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (62),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (70),
		.IN_PKT_BYTE_CNT_L             (68),
		.IN_PKT_TRANS_COMPRESSED_READ  (63),
		.IN_PKT_BURSTWRAP_H            (73),
		.IN_PKT_BURSTWRAP_L            (71),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (44),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (52),
		.OUT_PKT_BYTE_CNT_L            (50),
		.OUT_PKT_TRANS_COMPRESSED_READ (45),
		.OUT_ST_DATA_W                 (62),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_010 (
		.clk               (pll_c0_out),                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.in_valid          (cmd_xbar_demux_018_src0_valid),         //      sink.valid
		.in_channel        (cmd_xbar_demux_018_src0_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_demux_018_src0_ready),         //          .ready
		.in_data           (cmd_xbar_demux_018_src0_data),          //          .data
		.out_endofpacket   (width_adapter_010_src_endofpacket),     //       src.endofpacket
		.out_data          (width_adapter_010_src_data),            //          .data
		.out_channel       (width_adapter_010_src_channel),         //          .channel
		.out_valid         (width_adapter_010_src_valid),           //          .valid
		.out_ready         (width_adapter_010_src_ready),           //          .ready
		.out_startofpacket (width_adapter_010_src_startofpacket)    //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (44),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (52),
		.IN_PKT_BYTE_CNT_L             (50),
		.IN_PKT_TRANS_COMPRESSED_READ  (45),
		.IN_PKT_BURSTWRAP_H            (55),
		.IN_PKT_BURSTWRAP_L            (53),
		.IN_ST_DATA_W                  (62),
		.OUT_PKT_ADDR_H                (62),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (70),
		.OUT_PKT_BYTE_CNT_L            (68),
		.OUT_PKT_TRANS_COMPRESSED_READ (63),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_011 (
		.clk               (pll_c0_out),                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid          (id_router_031_src_valid),             //      sink.valid
		.in_channel        (id_router_031_src_channel),           //          .channel
		.in_startofpacket  (id_router_031_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_031_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_031_src_ready),             //          .ready
		.in_data           (id_router_031_src_data),              //          .data
		.out_endofpacket   (width_adapter_011_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_011_src_data),          //          .data
		.out_channel       (width_adapter_011_src_channel),       //          .channel
		.out_valid         (width_adapter_011_src_valid),         //          .valid
		.out_ready         (width_adapter_011_src_ready),         //          .ready
		.out_startofpacket (width_adapter_011_src_startofpacket)  //          .startofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (89),
		.BITS_PER_SYMBOL     (89),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (10),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (pll_c0_out),                         //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (clk),                                //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src5_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src5_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src5_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src5_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src5_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src5_data),           //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (89),
		.BITS_PER_SYMBOL     (89),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (10),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk),                                   //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (pll_c0_out),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_005_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_005_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_005_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_005_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (87),
		.BITS_PER_SYMBOL     (87),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (clk),                                   //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (pll_c0_out),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_012_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_012_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_012_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_012_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_012_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_012_src0_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (87),
		.BITS_PER_SYMBOL     (87),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (clk),                                   //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (pll_c0_out),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_013_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_013_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_013_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_013_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_013_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_013_src0_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (87),
		.BITS_PER_SYMBOL     (87),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (pll_c0_out),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk),                                   //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_012_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_012_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_012_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_012_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_012_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_012_src0_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (87),
		.BITS_PER_SYMBOL     (87),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (pll_c0_out),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk),                                   //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_012_src1_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_012_src1_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_012_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_012_src1_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_012_src1_channel),       //              .channel
		.in_data           (rsp_xbar_demux_012_src1_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (69),
		.BITS_PER_SYMBOL     (69),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_006 (
		.in_clk            (pll_c2_out),                            //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk),                                   //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_015_src6_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_015_src6_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_015_src6_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_015_src6_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_015_src6_channel),       //              .channel
		.in_data           (cmd_xbar_demux_015_src6_data),          //              .data
		.out_ready         (crosser_006_out_ready),                 //           out.ready
		.out_valid         (crosser_006_out_valid),                 //              .valid
		.out_startofpacket (crosser_006_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_006_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_006_out_channel),               //              .channel
		.out_data          (crosser_006_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (69),
		.BITS_PER_SYMBOL     (69),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_007 (
		.in_clk            (clk),                                   //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (pll_c2_out),                            //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_020_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_020_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_020_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_020_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_020_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_020_src0_data),          //              .data
		.out_ready         (crosser_007_out_ready),                 //           out.ready
		.out_valid         (crosser_007_out_valid),                 //              .valid
		.out_startofpacket (crosser_007_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_007_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_007_out_channel),               //              .channel
		.out_data          (crosser_007_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	application_selector_irq_mapper irq_mapper (
		.clk            (pll_c0_out),                         //        clk.clk
		.reset          (rst_controller_001_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),           //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),           //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),           //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),           //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),           //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),           //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),           //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),           //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),           //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),           //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),          // receiver10.irq
		.sender_irq     (cpu_d_irq_irq)                       //     sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_004_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_004_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_004_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (ddr2_sdram_phy_clk_out),             //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_004_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver6_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_004_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_006 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_004_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_006_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver8_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_007 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_004_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_007_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver9_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_008 (
		.receiver_clk   (clk),                                //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_008_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver10_irq)           //             sender.irq
	);

endmodule
