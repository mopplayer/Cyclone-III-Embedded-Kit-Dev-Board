��/  S����3�c�ub��_NЀP���t�,ï�!U;�P{�g��Oj*�x �*�'|�N�Q]/]	�	��"�l��.b�4;ES�����m�-�a�F���yx �7�����d8E*���뷕eu�dl���M��U[kUw'�K���hL�H����,!f��{���T�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P��dO�*���T���.+�]4�k���A�faؑPb˗�	�SD��H�"��|	��3+�:/xUW�2\Em.h���x��,$�LL,�֌mg�R9g`��-��Q��������Y�K��� X%)�M���mY�zwF����z� c�|Kёv��s鐻��	ABP�zi0�޺��PY$���=^FNS¥Ɂ���.�l��eDɇ��*�[��S�E�hn)l@��JGi�Z�+C4�[^y¢���su�HKVO7�#Yv��[�S*��#G����J��>�X��7a'�|Z��o��SL/4�L36���s�u����
�e( !�G�d��e��ڪ����_W}��9�56.�!"'뜧h�RQ���i��J�t�i��N^ص�q���E��tJ�J��J[���#���B���I���[�d�\s].��*��*E�rR�򹴸9d�iۀW���[����_����f(�s��݀�p�T�����b�Jo(`��u�EUtPup3\}�Ԝ�Eo���jk? ��LY�
~P�2Xܚ�D�qv�Q m�VК�.����\��LA!o)�!�m(���r?M_�U|�I#[d���q��ߦ?\�0d%p[����6���2!�>{�~:�h�9�E7zZ~��Tw�U]h'�\�l��|�uG��y�?͚'��r\9C[�Ф%��DM�~ddK��d\T~�o{ZK��3����Q�A��P����ţ�vr���+'ۼ#�����ʆx%g�����q�А��~���ڈ�jؑ��������9c�Q�E������Q���3��n�����b�d����K�k����݇9�A�o:���
��J����^+�mn��'��hN��B4	 �(�aq��ӢTM>���Wݑ��p�,B��y��\�"?�ϸ��(��#˯��;w��"s�����55D å��S\q��iq���4]9n��%��+�ob|>E̍��ulݸlnA<�dRIy@�ak��Y��uye(���% �*�IF�r�������ɓ�������jzf�C����B?�,j@H�턾�*a��Xm�㙻����Z����`�8���ɫ�*�q�����ϴ�2Z�:�4i��a!hV�_�E��w$/ɟC7T�*�,x��ju����86��\��uW�C� L�]�cNo�[����7�A~�'��*�vX�H�ȵ'��;�B>��Td�D���3ǹv_oC&D��V�6�����^�~����� �<���J��Y���/���h9��-��X���܌E�:�_Z���rJ+����&%�y��C�C���R����,:��Z�Cވz��7/��d�5���[����1si��f�j�%x4�v��%CXe���Z�v3�w�����Xxz�nb���i�M�л��4��ң���K����()�����G>Ozj<	������h�y-;�-?1M�0�=&���.%Mv�����%��8�:m�$�bټ�E�֘0@���r��[���Q�9�<3|�.���{�B4�q��y�����T֤�K��0\�� |���Ǿ
�kG9���O?[�rUe�lv�����X=99W2�%c���%LP0��m�)tL��?��|�x�� uQ���V��H���Z��b��6�	h�Dl��k���i`e+w�t�7��*H�_@
��&퐴F��ٰ��[x�eo�V%d����9��g�8֚�v����#�*(rlwַy��T\�H�sǎ�ޚp��L��Y��*[����gs���82;�]�iǖy�М��h$�j�����y��� �bс�iE�-@� �*�P���Iī��X��A�rO'6�0�I�"�&� Ѥ[�_,�8��=�+˪��F�Д.!�N��1�Z�$�������0��K�p��"2���rMԗf��<	�d)SX��
����L��p#Nc:�Tw]��S�y���D���dahe�'	<j��wn�T�p	~�JA��W�~��V�#�Ρ��U��i9�K�"�����GF���q����~�+F �3�ĝRVF�C��Mv�H��[��z���c��@�1�Wp`MY:�q[N�M�G݄l��4�SeG��"���6��2����\�y�%��uu�����x����-�-���ю���J��՛�)@�28@Td�X-���,w+��s��r*8�D�؞�����1��K�c����[l:8XQ8�����	*?��3��;s�C�PBS6��:Q&8�]�rr��87��rS�{�K�v)� �a���|��2e�k�8�VE��pe����e֋�tK*q�/���W�y����G�U�X�?8Cf��9���Q����Lu�&����KKv�H�NƆo �b���hh��!q�!��#�����rg?BA�3o�қ�W�~�m�U�cC�g�ύ<6�sKi��q;�]O;z�2��c�B1�TG��Hm�p�����0k\X�و���Oֳ��>�6.;�� ��z�ԃ_��$G��\؋!D� 8_r�}�5���k��UUY9�Ô��8�mXp��α}��鮽�n�:!�%y>��Ɨ�Z�rw-yBt����2{N�}��n�G�.8eCj|��Ǣc��\E��_�V��o�?'�=ںw�����٫��Ҳl��g���6^����/ш�-�hY�uR����!G��i�"��-
QvL
��Bu����D��p,�`o4<��s#Ǻ5��!�(6ѷG2�?[d�Ѩ\��$�����|�O	Ay�˕+�B������Ed�*�2�-�o�,8YG-D��	���&�a7�W�E�l]�iDE��Q���!�:�e��$ߖ�1�����c#gf7��.���L��c׹�|�/�*>27�Y��+@��;|��'nt쀍�+A��2�����o�Ks@)G���V �����q¯4��V��,�ւ���$���t-qz��`��,��
=$�����q}�U
���~�Ń�/up�z�n��T`\n5#?M���NJ����&��#.qѿ߲y��-��8@�V�)�����ƛ���F�;es#�>����gl�IG��9���k�^���7xc��l�C'�iH�p�EUi�l�ӑ�u�>O��h��?�Z5$�i���9^}��4�T��fÏ���;�  �8��:躵��<�S��@�~K���d�R|@x���7�J@���Zuܢ}�I֒��ʒ�*�C��p�o3���f��6](np�(��Tz��Ȇg���0�m��j�J��e�ld.T	8TO��ׇ��L#�A<��� ���'�&-\��e��k�kS�akh���@\�k�|�+i�a��z��9�]B�I���(r4�Tx��d�:��m��͆�-���v����\%o�DA� ��������5�;� �M&������71��4��=^p�B.�?��P� ���`�L�Gڰ�d`����4S��ӓ��|��������-sڨ����Qc"*D����bZz�2e EY�~�A�%�DL}��*i�d6�!�h1{t�U��E�0R�M�X���h��2�k�h%45BcSjNo�˿��G������$�E\���i�r>ݔ���_����9����Z���g�g��YM�D��x�'�B5�Ȼu�҈��~;��vQ����]L@X�<F���z�ºy|�#�^̴h�]'�1梁�����4p^�X����¼�d��p�}dݳ���F�Ȩ�B�8���y�߉5�JHu4��b6���57ՏH�A��:��[�}j�����ji�Wo�5����:�op��*Ɍ�@�0�+�J���!9��01�{��w������LWT'�ÝZ�¬�:V Wp��x���� NL4��j*�O�u��K��L���|������>�{�&������'��ɛ>��g�J};m�c<�����61�M���g��'�>\�br����*����?�+��n���)>�^�`wO���j�I$\�W[V�ݫ��wǸ��i�=����f@6K�����5#��n_q��f��)�T֤� }.������|�$CƂ>n?V����$���(��n��i�/m�T��c��MT�;�+Dpji�X05ǜ_{	���#�$����ˍ���=�Ғ_|�>9X|��2�p\�dPMˊ�������|�	�xe ���<P�n��aC�S,TJ���S�?��D�w�7ye�P��4��8���e`۰X�Ժ�Z��.�׵ �eON��TxW�W�[�WAנ1�?*K�͙�������P&��;�2r�n��wZ?��*j��!� `�׳�g������HR�P?\@�yPP�<�9K�FSe{!���t����86R�I��1q�+QE1m�Aim�xێ�̼ذ��
�[ȰQh�Ь�f���&���U���J:WR_0_ .��~��ۏB���XJf�h���]�ł���T;���6��m�G�AO�����4��XNM'�G��e���~Z�Ix ~	��n����>���cD���肉�*
loW�J��u(i1���9b�x���(X����.�����^
ܫ%�T�=�	a�ԚK�(D�e&�j����ޖ�3k�o��#qn�X�ʧ������. �r��Ba9<F�;�f(��ږY��yMQ��0��Ԛ!v���g�_�普r9a��&�d-��;�h��%���DCI���]k! 1Ot6�GQ:�5��c�Ы�)����9�Z�}�
	��=A?f�sV��&��"A�17��	��M��N
��*�V*��M3��a�C��k���Nq�(�A��ď����z��\�i�eW`��tס��J���f|�*��縷3=�S��м��5�у��m��zV5Һf�g�����ֽ�o��J����Rq��"��v�cz�AX�N2g�\��bE�y�j�se��	�g��x�e'�G�)��?��_��o�/W� m����>��\W{���� ��z�Z?�J)G�?�Z�-�2As�������u	ŧy��h�U&r��T1f�^p���:Y�i�� UH���s��T��>h�b&��y��~-h� z�ٖ��1�����������}�V%��c�*_<��pK������l�"�,��2�7���I䵲nG�'�b��RY 1.>.8�/���8rX| l%����*���HB����?2^��j�� �7*G��8��B&`� 1x�BM��wlK�G,\��-�z�Y3Z�	/�%0��Ui���y��0�n��(gxWb����j'r�J�{�V�=��ܯO�O�^HSue|���j�s$]��T�G��
�d�w�φ����a��c��+����lQ/}��`Qy����ל��塞�"�/�/NG�Rb���nJ>��I��kL1��3����õ��:K��l`:vY�Y����2�jF��E�j���2�ɧ@sق�z��*�>죨��!nQ{�̺h� %���-&���))�����
=��0nie(WAl�2���Բ;��?��l���+q_~L3����!#V�Y@���u��`'p6m�^um�7�mƮsp�1����;~18-�j�B��9�!�`͞��E����j��c.?��NW(�
lDr��p��G�OA�fF&ɉ��ִ�;� �|}3�+34vY�y�s���7T�K$'�b/��7.!tN��4ݾע��/�xL|��p������#Y��(�?���k�[$�ƀ��Lܸ��EQ���ypR��OR�Ӫ�VE<�F�C�"���\�v��K�e���hS�����Vh� ���'c�٭S��Kh?0_�bJ���FNq�ezxu٠��.�!*�Tv��?m[�&�p_�i$�KEe't�f�~����`nD��ێ�zo��xe��R��"\�H#(gpF�5�|��ר�h�X�����4�=��s�r��c�ȼ����0c�=��=����,Yy&��;�WF4�|[ ������Z-8\���l_���4J�=�#l���5�.�Dz�X�G߫�O����]eHq����,ID �zA�0Ӭ��4ً3���Sc�v��[C����fD��'f��L���j[���E�2����u�VJ��ǐ�2����%���/-T��A.o�%�蟵�\�>�������[�:����!��0�����s���,,.۪]�c�x�M@�*�ܵD��%���k��y�4��Za��Hn��\V�~9j�7a��mH���N��k�\8Ʈ۴���C߳�QR7����u4�]�C#ٶ�:H�/~����@:�qj2�	�*��9�v��4��O��E��oX}�����{D�]�ǿ}^��e�rH����[�cXk-�ckl�ǿH!���mI�r�!���pe���K������ցv��D�/���$#�~��7П�C�H������a�<�<r�d�� ��Ӻa:pw�^��Xa~����z)���=�yt���n�8��Ɠ��m�?	�acz�Ƣ �z�.��5$�#~Pd�
�U�5��ݢ��.v�ǒ�V�!
��D�Z�u� ��� ����t�eB!7���{���3���T�Bs��7��p#eO��6>�>�������՚[;�R�^�V��&�Cd��ntζ���ҮQ}jБ9?-�7��zS:��W���]Ghʦ��݌� ������F�V�6�&��!���R}�X�|.P\�>:HlEJ�I0��b*��Q�su����R!�/���_f����#y����$w:m�k���s������ˊ7�|�i	�c'L阚��h��db���X�OK*Gv1]��z�0�A�̡k ��	��6��1�Y�!!n���H�(��!���y���߇U/��� �,s{o�;�[�<���M1��:��f#`K��� ����&�����Z�!� d�[v����J� j�G�@UA�x\��/l��R��|Tj�C�C;��q^oǴL桒���6���*��fՉg�-�\�i߭�rleY�Ć�tg!8����A*s�d���ep�I,�ŝ&�]�:k�c���6�^I9�Xk�T|vW�!^[m�g�z���fפ|�0�#�)���Ҡ��%�%m�Ģ~��0�wa���6�"a,[]�"�O�Tf3?����F��c�5�:���1��$�h��[�h���w���F3�\W��`���@���a�q� �S�z���쿍fg� ���q�NYH���Л|�R�#��O+����� _4��c��5,ch�co�ݛ�{`r�q���3�
��p����&^�T���qYD�@�l����_�f��Z���'�Bk��hEm8 S��jP���f$�j��l(ɩi��W�X�m�}��ӵ���-��WBeS�"9阨/=y�`x���|ﵪ�{���m�Yw]TY�?ۼ ��w�m�6���Ƨ���=�oJhǬ��Mc��P�q� *��Zݔ��� L�Y�LX۫R��=g{��״*�O�'�Y*|�.��-X�ɂഌ�� ���J.)c�^��9�{��y xd�3�~��f�?����!��Җ��e/�t,�/,G�|����=MSn�+�a:8�>�G�_	��t;�Q	 6YQo��d!���kJp�{�
J�V���(��nq?Mny��NE�7RD?V,�ar�m��ʑ�*73��zxV����S!|N����5��}u�s�� � t10��zx�=b_��DeW��^�s���nF�^��v�g-�DBI�jZhY[��UO�74��Ԕ5�_�E�\�5=$�'����� �/���̤��]�p���b{�#$�������^0W�E闇� %��9���k)^��ϣ?)��3h���[͙�~�Z�Ȑzc���Lx�F�����B;���kD�C���?�Yku$�[ u���d���5JRtn-|tX���D��TEcK���!oW$�p�p�/�]��
~R8����U���(�ccH�"�hϫfK��g
�bk��T�<z,��.d�Q��s�t�dg��0�tt8S�4Va�C\��)x����:� W3B8�L�N͛J�'�s�GpJ����Z��uY�Y�#��ho���R���A$U	�,a��Rީ���f_I�W8!=^Aq�`x��&�ϥ�0|<���^���>Ê��rm6a�i۵���ˉ^�	�QRn�Zn���M�Ya9��m;=0�|0�'��ؐ��lɬ=�ɄΟXD���]Xn�w���U~�}�E~�����J��ϰ�a5jY�u�-��"�{ ����^���nZ�.���Y]m�!h�AX�ͥm������Q �^6,1�y�G����y��'�Iu�6���1*���7TM��0&P���ޫ�k|CO�n�><�n���B@�pEe>z�҆� �]#�s�a����oZ����ؒ]j�=M�������ܧO��gl�?N��t���\x��>:����E�d��<���	�cް����fS�c9�)��d�����N���	��?�T���"=��"��ܖf�z��]OM+��#C���u.�`R91�0c�
I���������M�U�� ����A�f������}����;r.(s�t�o)
����e���Z�]�d�MX�?vR���*ԧmq2D̝��%�i9��(k�~/_�x���xX����3Sgv5��[��2o� @�>>�=Waʲ�v�����
���H���;�[i��5�_+�5"=��\48�M5M%$ϛ#���;�ݭB�}i;��uJ��KGd�YXz|5�9܆�}
J?�N�0]L@F�^V�:�{S�=�PU�.O�����5�(�TgVA³x�cc8���@��U����f��7���"_0Ya�PpS_KM�+���T���*֧�
#~��Gw/�P�'z��v6b���>�֘H�U�+��f
�L��԰�rC��A�X�)Z-8�B��(8aay�<��-�b��,��
r�B�}�%,Q1�e!I$�/{��~贛�߻ц��c�pǥ��>c����U�nƥDnf�݄I�))6�+��U�
���H�7��F�A�Yz�$Rz����-��F �=s��f*�"��S�舮���V�n�E�0�,�e��)�x����0�X�,<�JX���ĞN������m��ՔN���t
ؗ3k�߯򹓥�B��ғ��-,�z摁F���Z�[�BGpƙ4��d��N��{�ͦ)�36� sf���	��%|���d��+�T��o�^0�M��N�@�T�����˃u�8J��O����M(h���dh���MU:�m����.y�^�.�+B+w�j�j�;%�.N�:����.�����|7���#��%������Z��>X�=�I@�]�}ѻ	��~��ǋZ��ˉ�z�N�j�5���NT��Y�x�󤔇�W��������F�:C��ȿ!�,�ؑNb`�� $�ޙ/y\���;ϰ�TMv��u��{��ȣ��w ŝ��6����k��?W�t!=y*� �*߉z�k.�`�H��F3��x�Qu�C�*�q��D%��Ӓ�����d�Mi�e�.;�+����L���Iï���R��#�mWe5@D냑��]uԣ��z�&S.�值�w5���pc�̏�;S׮ٝ�I��NL���[)?�C����L���08@�%�� ���k�����0�T;��.(m*�,����`��K=7��fZ�nw�ޕ����q�C6���.<�m���~��IZs�H6�A�$�3Ž�-x�5���ĖO���H�#����c'�N��a/���=Ws����p?,��ʏ馰�K։���g�5���z��%=�0��������~	�B�<�(gP?6�2� ���ސ����u[�໯����x�M�ӷ�\�m8L(��-.�3��]_h+��H]��
���]�������@��A�僄�'��ݩ��*���^�~w���l��˧� ��q̆�<�LD���Z\6�乱o/Ԛ���5�B%/�Y��g)�MԒl(+ӭ��w~(����)� ]����f�����?0hwj�a�OHU5��'����-:+���2��n��k���J_6�6Y�G��OC~UY�G(Є��;�W,,�������[�W�hj���&�'����&��S}Z^��������Dͮ,�]KS1��~�˪�׻��~�@�(�1�Q�Ȧ��*hڭ�߾�j��з��}u�̔ac�3���>?��eR��w
�ή1���0>�t�� L{����K�r.�_p���4)>EN�����J
֡$&u��(�$l�\�.�óg۾q�h.��纈Sٯ�~��ϊ�$��[O�	ȡ!�D�/������fM�z�7(`V?��\͌;]O+�HƘ�-���Gt+���)?}k��C^��:Ƽ�%�M�X+����E�X��md�?�6�o�;�?�J�m�!�@��g�P0oB��-�h#�V��	�h?��n�ԭ.���c�кt����1�>�|��5)��������/�:��ͨ��4pm4��ζ�N�dV�甕/0����h�T:��3?�(6nTd�9M�e/,1�^�{l�\�*���\&�$(�z�XB�癝�1����.�R�,�d)���䲋O &ϼ]kyo`�kE�d�m�7�`�a�r������f��g1'�<����[�c8�)���:�BY�n�`*]++F�������o@N���-�6w�]_�Dk��>F<^���Ag�8���p�~*��9_�{ñ�䞷P��>�2��n8L�a`��jj|׳S���H@� 
��<���O��N��qPqn����1��Ϩ�$��l�c�^��+�fh}���.�m����g�U
��}&|��h���mե{	��P���HV�oaH�Kyw�B�6�6B��m�t�Y�|�i�_'�!�]��0a/f�\�
�2��l�&���IR�&�����r=�Hz����u�:��R����j�� ѯ��	���}R+c6���x)�'s�d��#�����\$���-��EdD�cʋ���}���;��h�{�� a���Q}q�\�vBwģ�Y�O&,����KF�=�1H�p�fځOG[���y�����'�-�V���\
���j�Ž�jͿ��I.<Mz��l�/'�K�p(zV�p�̅����a�'��~v�E��{w��y.;�N虭y���S���N"?R��z�� 5Zm��1rr���
�a��H�Ȳ	�k����3�|3E��7�n��hBَ�A�t�r�)�E�~��!/`�9��r&Mr��{��a1���	��BH�w����?�������x�o��h�I#�t4Cѹ��>�7��3��m�[PF��)@p"{��Y�+���P�=�)=y���povK;ŝVU2��D�ZF�BL�^���p�
�+�q#P�gHAY��nb�yYB<�w.��"�ڌ�b��9Xq��2=�U�nLz{*���䅃��UO�òJ=�����5��(�[)�[ð^,����S�(�G��@=�pth|�ڟ�D�Іq�݈I���i��P���y�8/b<��!n��\���C�M]�xl�|���f��隵�Q��DJLZQ��d��j��?�EH(Ԭ}|7i��d:5��1�k��?6D��E�'qy�����[��*?1�(�C� N��c>� Ce&��B�%H�P�%p�����'t��Q�g� ����nEH�ɵY˶a=JR`�f�V���qϦ���4�Z�ru����K'�J��"�rȂp��s>/��b�aѳ���
|`p�?؎|������#1{�S$d)Np/(��,�zŰ�Ԙ#����8����ǒ��:�؝��c��	}1�w����;�*bB|�l4c�Z���S��M�.a州+�G1����ׂ���q�B�q݇~<|N^�ydP�26�\:0!P,�};]���%a����E ��������+\���x/�,��钑����2��R������u���o�4��C_��(K<�� y�|�,��-����G�X��$�SspqGq��Z)􂿅tt�=�<���U@..q�őcm�~,;N^<�n�����G��4��&ξc1���_oMAJ��J�n7�_�@��W��DL��р{�c����l�a�?c�9/(�t�l�S��"=
^r�p!ŕ�׊㜙V!�\�ɞ'���}=ǂ��i�Ҩ׹"��zX���� �{%2���i�>&}͏��}�7"2�noT^��V��?����ݽd���eĚ��4��
�3�����k�2_dR	ڞX�@ c����h|b��dV�պv7.@�k�|���Emogg۳������ &�P�;]O�dx#��Ң �~��W������NtI��C����:�P�Y�u�G���JXuK�%1q�T������([�^Y">f�L^��8ρ6}"CZT������K������.��?�>���&I,k7�U�l�&,��<��͑�꒷r��^3"�(���[;���RG��� l�а�B�bHv�k�<����!�f��ښ�;�J�Mx����9f<�1!Tn��'K�%,�6E��@jk9xD}>�rq$ �{�!���,��3�����9��ӽ���������&4�vOR�����U��o=}^[��9%�|�[��B,ڄqGEm4��I��3\-;���P��wf~��E��Q�{&l.�"�;�G5�1c�g%��g0cNc[���r�l�a�Hol=t�M
���]%d��ds4�Z]N�݈ꔌs�l���`=K���@�ro&�L��}�
f6�!v�3�ؿF4p�DO蕛E��F�e�F��%Ŝ�����Q���g�ǚ�������
k"�;�?J��]��TW�K�&�/��$#jQ?,(���j*c�ެY�{�po8'� ���1�b�������(z�|�-s18�N�˓j-�UE+4r�o�Qqv���3��H�=��t5{�\g��>�BÆa�>|�Y]�=�����H�5�P����q�2��O%��mzrT�?�o4��Մ*w/��^��u��H��)8C!�/yY6�yȲ!J7�(݋�ov94S�.����h�:a�I{a����Nǌڶ�*ݥ����F+���s�7�eh�9)�e��\O����Q��>x̾�cV�T�P�m�֚�1�d�m��28�sK$�Җ�OȄ�z�I2��b��Ib�NVGo�nf���9I�'6O��J�sDE��^'|��n}r�ʰ�p�v��^�\�����_�a>�?�[1& m�]H][��T�x 5,�w˹E(F�o�W^l��8?hޤP۠3r�� Fw�L��z`��,_u��3����l��亚�I)&�'S|��o#�D�]#�P��*��Kyq��Ȅ��c�}*��`Y�i�Y���lH��g��)�T���`�тY\�t������{�'}Zz[��`��>��p���E�)�i"�`����Y�2v��d/7�ϬK�9��GU�fYuj�S|T}.��E������'�&х%n�[5��>���� ��?`m�6��$�|9�:���^�`i�����)
2|D};�'�v�z,�;Mg��+��/�i�N��o��y�˼��+p�N��A?��Ǵ8#|o��!�zӉ{릵�7;�,`t��dKs��B���ac?W6��`2܍���`�J��6{j4��g��A�(Z�C���.$DL�x�'<F�07�6��}2�)XJX{��,�x��\��ę�b\��ڟ���eV�c<�S�_f���|�ha�������̒�>���}ˋj�� �~�>�sΙY���Ad������k�/��+I����`�2������A�Ǒ�ڄ�P����6a#��Y<m
� @|	�"�n
^-�\f.Cm��`�u@L�A(���ZlG����0�d\�{�a���u����X���a{T~�����P��L��L?P�T���P#�
��Ηo�16bOb�?�����֗o���H:ß�  ���qosR0��� �1�2?�t�X���&"/�YN&����B�MMOc�
��؍{GRL���r%�E�� �;�U�S��Z��ڣC�*����\%�!��(���V��Y2�x������|��KJ��<��x}��#����r/�5�Ka�q�܀�0.vZ�s:�&��T��e.�P���d84*�����h�ዌ�؋�a~W�M[��T/6Vh��τ�[2�0�2�Y�Q_:��|u�%87,vx�wO�񄁏�,��hd	���k�t�2��4y8
i0�9^~0J^��Q�a�����T��7oM�C
<�y� ��u0I������8yO	��@u�E�@��G�~����`�F�(b�Mn�q	a��s.x�R{flqre�G�[%�y�� 嘌:��i��_fqں��O�F>z�[$ݴ��B��1&���o��m#� 2\|����5����?�V��tS��6�s�'60F.-$C�|�=�����6�c���޷��/ơ`��D����+�T(^0�s|�����0�,����6����:�E@��V�dpK"B�}A�ͣ�1�.��mj�����������"� �N򵜠g��kx���"ak�*:-0e�op;�r�TJMx�5t��a���7=׶�U�(L�_�An;R���ir�'�/6u�K":*gփ0�Xd�����Ԙd�;&�*�,�=/�"�w�l/��WR�sک*2@9U(L|���G�59�����\�e�E;��������~/l6�檪���}e-��עNe���{�v��'v���aD��^�TuTkDCy�=������u��_�h�4�.U	������Ur�V�*�F��T�3����lb�U���3 9�i	�.B[�7M�R"�m|��r!(/R8�e7h%���Þ�5y/�j����>���P;Ľms�U����]�2nD���cj�]�����S�n�[�;jߵ|b��M�98D�j��Lc�*$��U�.��_e��z;H�=�օ�{`݌�q`n����&cC����֓��4�!_{��|1&Q��[�<���08���=n�jj?!� \�,� Z�-	�h[=����tlV%<(V�-[���A�V��qM*D�#xɗ(�V
�G�Ƶ������*����>7���:�ORMll�	�����E�Pn+�q�Ĝ��3�TT)�G�U���
�τ�x(�W�6~\Qf�(��)�@�@5�KAl��%���`�B.��,4
�"T�-�n���8�p+��>R��ز1�<�F*��D�آ�7�6��t���Q@aKo�-�ղ��X;��J*t*�Ba��j���;��}1Yvʩ�pBh�%��eݴƑ���s��pj����8!�-��k���S'����(a.8��� ���a�Z]�dDv<�m�c����O�� ��k霤��Dc4L2�J�� b�\�u6~���:�-x�M>���Y!����� G9�81A��Џ:
�r��w�5C��fñ%h�{��@�!a�gŇ1�^G��&�A�dq�N{*H�������:�ǙT|Ts�@NO\4jm֧W���J~k�u�>�}�qr	˜���,��������.B� /����(e�d����K��A��V��9������~�h���.��;X��PX���]yM��=ph�?&����['�O-6����Y�(L�{B���7���/F�B3Z���pՄ��W���_�2���vS�Yr���uY ���O|w�
��*R\����hέ6��ً�\�a�<,�~�F��+'u���>9���e�~+�g���o^��a� �k��Pc/�xBʯf$`b�H�âf[m�C^�v#|�+��q����ۜ�@Tq�,���+Z{l=svvk	}r�Eo2���eRl~U�E��V���o�dn*.�4�n�L	�t��H�z/�{��R���+xfa���F3E��Ҝ:��r.�<���p]%ɬ��m�>��5˨�P�X�b�l�\������c��Wʊz������k{����v�7��4�S(��:H3���C�U�9���ΐ�x��8�$�ZUI���g����������Pl4T	ܦǁ���s6H�T��p]T�x��9i�~pZ�0��U�9sM	�f��
��0ڿ]����ޔ�|�p;Tܔ#o?8���?/�aQҊ�5T��Bp !�F���$�:��L<�`'���P|�?�����B��4���q����<sy�V159�H;]0$��C��5z��t8���.�%%��O��ucZ��xct0���#�H-2x�u5P@��4�Q1Gv'2�+esBM����r�a*O�E=W�k���$�r��
��_�4���Zg��ҍ�����ǋQ�N�Axx#,I��L}��gt�H��J��u �(�;E�Oc",��gj�Ы3�j5\�}��w� BĨȁF�f���r�����P���*XY�	�D���%p��Y<�}e��kH��{^�~��Z,@vL� �\�񰌶�N-7c*�1�RQK�|��Цٟ�柡z>�R�VC��q���z��	 <fٱG"�x��/�W*L�;t�8��q@�<���y������3'�/�$�FE֠L>:�@�%���&����ވY	�_�W-v̹Z�Β`*.쉇�v�6��S�k�/�#aa3g�}8����ҙ����B<Κ��N��I�G�#l<��.���C�h����^r��"£e�[�qWQ�K�<qOy*"�:��Q@��r��T��	/�{.S�ԑK��ݗ��E>MJJ�)�ɷ̘��D�o[Ȱ,K�0���m�f��a�H�	w�Ȋda�?R�t��_H�!�7���٪2��x1�G�`Po�$�+���_5]P�r�Df����B�rj�����s�iyw�Y�Fn��"���=�7'S�w����:9�$���a�l��LMs�-��}9982�q���Ѱ?�T�J�;e�!����?0l���&�1:z��[������N�͢���̺�Դ,K��T6+�fީ�r�$52�-Y�O�Tp��2���T��f,*"�\�TM����7Do�oYu��J�=RX�P��S��!eq����K���\v�<X������Z	�2��M�Ǩl�'�W��1^EC��7٨[,�ɖ�y����ʂ���MFFL��r�A���.Jn����ɜ�W{�&e��b� ����
���E	ذ�#����(&$7&;��-����,F�WF�W?k�-/���j&ؗ�L5�l��=��ƚ?Go�q�Q�$���v�u�MbX���$L+������?��5l��L��@�[�C6N�4��`�]h��H�H�`/!!�	'L���Xʑ��v�������n�4��U���}��O F+e`! !'�� �.�t%�{��7g*�G�TX�e`g��.�����y0W�� bs;�Bć\�q��������(�J�;ӵu����2�ד�b����$��g��YuY�5��"���*����+jOL�q)�o9�з�gf2�J4�)I���fƎ`�m�ą*tP��i����]4�������)�A:fԇN�mb���DM���,���"��@M�l";fr!���#�����^*v-�n���p/�σ�V�T�o�n�����l���e�5Ytr5ڬh�~����4s�O�}�v>6!C�hg��EC�)�&
>\��}7y�bӬ��6�{��Me#��J�ug�D	~�aǭ�Xl��13�cF,����ges� H�>�>��������pH��q��F���4�ٛ�H���$����I���d�\9̢$�2�������p���P�H�i�< ��k��a�m��� Ao�C��|�9����e�T�Cs��LZ1O?�6�/�����n���U�S��U�
� �!TE��9��9E_�ؼ�ߌk�$�m[�_;ׯ���+�^N�0�-�Mȳ�A��Y�{� �r���}s�ͯ�7SH�y]�����ƽ��ʣϱw]��1ҟB'����<a�������z�{?.�$V��{������E��;� [�]E����(V8{4�0��6_Q�;&{v��G�$S�.���;G3Y^���P�4C�y.�@*-M�C3 2�ߔ�����rGϫ�O �Y
݈�r���|q3[���B-�b\]��0�
 �qSu�k?8�UJ�ؽ*���RI�k��2@���&��2`|Y��13����Њ��~"a�� Q~B�mSGD�Y�q`�޻�|bU���k��dhI"�9��ԓ^P@�|�1�3�TB*{l^۰|�E��+��hA�3�M��	�O�+�?Qԛ�~� `a��`�4���� d���kg�Q�oz�t�9��[���#x�G$��9t�Kf���F������8#^�eh��*�� ����o?��˭&ܢ4g�DO���CM%1�0��0����A�Ƶ`�H�)���|J�f�w1�l��İ#�⢨��a!��8/��>��0g��2��Ш�N�aR]���)���3n:+�_RB~�;V>��k��G$��Q���������h���K���`Z蘆���"s��E�B����:���ף9�E�gE�a�
�̲JÛ��£-�A�:�O&p��������P��� ����;<�g�&��ۍ�i\���{a��h�F���I(Iߖ���X� $�m9toSC���{�rҰ�s��E"K~X�z�%������'M$�f.FG���c��|�7�=a`��������xF�IOc��g�ׇ:�jA��w�i��m>�EvK�d�^��J�i3�S�Qx�|����1H����Ӆ�G� ���Ǎ��������T�IIQ4G=���#r���K�� ����r�bbF�ExꦝQ��N�i�[|���"؄�F 2��/�(���,���LPGt��G�wAY��&�vO��>{�'r�!�Vj�BƱ��q��f��k�T\� ��эS�.'+\�.�&܊�4%4u��ǅV����`3[��vF���3*�w:I�����)wԄ�׳�>����\�|\����|8���.gb���3s�"56{�*��V�5�,X�jB
�v�#8|�3`/Rc��)D�n��R
�n�}��r��m�	��������_���dGȸ�-���zS����}>���t1=�y����N�â��ɸxP���+�HGM�Ƥ#��o���ٵ�{��g*	�B%�Y�Y֚���6�&��s'�=��˿N?�ɑ>rhv��O�Q��RF�>��+[�L��΁��-��s�\@Y��I@f˭�~xŭ�vM�5'���c�Bh4ڳ�Ūn�j�N�n��<�J#�[e�Cz6��TO�ZJ��d��]�\�F��s��d�咺���XW���s�،s�oT�)LC_C�$�eV��P]���g�|��Hv��(�ʅLD�[������HĊ�f��u��mF�}WIL�{>̤�x`:���)��
�h%����3����Yב�E@+�D���>���sY�!�i4���h�?�m�*A�l+�4#S/�C�ׇ`��#��=����v�&�הD'Ü�.�b�r�o�l�Ґ7U�=/�;���	�)�x�>����@i oW
J�wXC̖8�����/n W�1��$�P2���~���L�+��0���1�����'�M!:gDy2��>�ڃlO%�ݮ��Б�j�u���B���]�F�(�Y\��p��i(�V!55��f��_�R��*���"Eܨ��s�c�LRv}y�:��������m
�� r��ԞV�IFLN���0F�5,�pbepO#��4�4I��˽�Òt���z��L��3Y�1��v|�]�gj��@T Y;�;��/}���� ����XR�3��
ޢjj�H�`{җː3��ShYԼxlSL��R���>Z_~����������Go��N5�a$�u��o�jQ%���6�����9�d��.ԕ�K
fS\4�*��w�����܀�"r~o�tQr������
5�Z
���O Y� �C$���h�d����Gyĥ�g���S�5	�)vH���'4��T�&&����4_��W|�n�͗�~��cG��%���'�WI�7�fe�@"w.(J�,�/qx��
�f��E;k$!q��C��-�nC�<�[��A�����i�=�:~��r�E��3x����� 	($XC��q��ť�˶��xR�7`LH��x�P&�2����˻e��*��ӝ����1�����I9���G=���|[���Hso-��<Ȳt��ǚC[N����H���ZX����MV':'��}^:��s4����{\��U���(��|��9)��'E0����H���)�/�r$]��b⵽ht�F0noI !�ȸ��%�^��XT5#�h��q��A��'��
$K��DP���Ay��^�C�ٍm��i���S�������^��B^��]6�c#��_�e㖅WZr�r�CL8� �/2�c��օ�^��̒
ؾ�O$N�wc�2�
���%��p���|~~K+�r����xz��U�W8�OG��Q�
ח?�Ӕ�-j�G��v�
e}���4?��n`�f!h)iIxY�����[��}\o�r�B����b$��Ͽ���q�R�������J�\��o:�w��)}DL���	AC�}O�x��<�_���1��w��*Fr>�?�8�6�#��!�)���%3��uXyo�T�16,��5WyT"�$�8)E�����6��sl�+�r�oĵam�%&�}IDH�E��v�bZ��W�18[@�7?ƚ�|#PW�6�+i�xe�/$G	�b��/�A���Qj�����	���]��R�jE�#��?�B��$��uQXXʐ-	a]5��9�[Oܳ�	]H˕�3:���f���.k�����U9�ߏ-��7ə�y�W9s�Sݬes�O�eE�`��� [@��:=�^�6��Xg>�p�� u�</���:�x�Ģ!�@��
����-�8w6xv$��+�GL*tĿ�T��)�XmH^�r�ѽ��=H�U*�%��VM!�S?�%S>1:���[��-dƥ^5A���ڟw�+@ASM�)4�&'�6:�L�zT	�?�Zj����]�y����CY۱���ze��Z��_�N����Z����$z�t�C�A��I��/���.��
E��^呰ȇ[�����<���8��ڝ'ӳc��:t$z�o��}�<�IѾ1"�8�~���`5��,Q0� ������]�ɩ�IQ�� ���D�S���PI�̄r.[�&��PU�X��McqZ�8I1��W�)��c�&��H����X}���s�z6�qZ���i��e��&�j=�=�|.eN����d�s2&���)94�|gy-^Z�Պ����r��b��r��5�:L�[�;�- ��Y��h�v��7�wџ:�ߛC;�)����3�����K���F�e%�Y�1�AO�����~�>�5�?�G�V�5b{=i�[�vvdK�k��}��2�1�fi����ߢ[����-VL�C�m��9]i�7� ��q�0�ۏI����O|V��h����J|�,��
�!��9T�J������]���
�j^�8�WL�:!f����pP��|ء1T�U0�����h;�����n�z�=<M�j����Cq�� ��hZ�<�ԧp�9<�.tҜ~�t$�-X�q�ăuv/.��35�?�"Cb�"���.ֺV�e1٦����ǃ�f�y��H��I��@�d��k�G�?��k�P;~�24� 6lqũZ�*v+ōI�h�%��|nm~��L���B kcR[���Z����_H-Kl
�����`���:�5q�l�'��q�E,c�正]J6��I`�` �Iy��e��j(�NЊ-���Wa�?u�|���f�j�{
�R2����P�I��+V�G���6��!<�W�a�$�i�L?�:1ހ��PED�Ý�K�~˗(I�����j1�oP>����R6Q�J�Z��&+�>���T��B��ȫ�U)��,�)�Z,$��o�s��P���@>EܤH�U���CO��4{�������ll@ն��5C�F֡,c|��"YEL�,��Hɫ��Wܟ�v���)����������!?��HR���+=!]��/��
�i��ǝ Ob7��S�5D�,y�J��Hy 34s�:�o�b)��-r��3ݷ�Z�l�V��ڌ���Ф��++ߵ-8?��R��~��i��f�9�t猚-U?�;[.iv~ZBZC��h�|1��@��A�B�������#"�ð�ywt��sL�a{�K��:��I)T��Կfd��.�d������=�K$*m�3�,�$�M����]���qrq���<���?�ҫ�ZE�g��D��Q� a��=�9�1�X��^6�k�%��z:�1âC4��E�N��I|G>/*�*�_��i�n���br�73����&���zz���c�N"��]wI6�Ѐ-��|���T~����5�l�������y�˫N�A����B~jv9��e�5�tw>`rs���m�"�D��x�o�ٹ4n!�^:���I��ln���(5R���V������۳���n �ߞ$�q=f��b?�l`�DM�s/�=� ����dԖ9�_���~�|1_��M ����u��yx�8��IT]:���ܴ32��f>��`���}E���:���1n����@'��t���]�t�"M�Re�5��gL�y��t�$�y�� gO�0����I +!^nZ��=���H4�3�~Bj�5;{\u>�r�C'v_�:zzZ�8��D�wz��c���0�HP���������#>�H$T���/,��U���M6��gP� 0cG �}���	�]����Yxq�Y� ��,_�+�:�a�;����/�$Y�5�X��Q��G������ ��{�P����0�L2Ws�a�x:�q��~k��ĉ��� ���P��f�)��1-�E�:`&���(v���&m�$S�u5,���ԯ<�h��n�i�.�p�նY����Bb/N�\���V��B\Ӯ�$�_���j�u����֭s7�lj��6=fJ��1Q ���>�����<�(��~�H����J��GHq��a��&�����A���#\FH{tq��'��Ykz�/V�q��CQ��$.���țԁ�m��ͯe�=�t�PH:rR���ƚ�'I�Ɠ��I��qdJ���f�}��P���w�+�d8�cqwԝ��pMJ �w��/��QgȲ�`��kE%ȊW��v�o,��$�nm�OG@'��;�t��C�)��LE���n ���5)���qA�+�˞qz��e�~,͈�;�����mz���Cu����WY�����O��֪Rk,Z�k�\�zV �F*1�{'�pu9��:���EdB�J0zې�>ϟ�F?���� �i'���+|K���*�I�>������w�͍>I��(�t2~����RE�x�v��)J�f�
����g?=��<��y��$j����7���b� ���M"`��۩+�D��@����q=��M�ŵq��է��+�=.d��TƷ����c263nh�����eYQ�{ݠ�W+B��.�/*a5̨S�oF��%���!!)�㕈^�]ZL��lXԌZ����/���PX��A���
��J$L��-G�Qj7��⑺|tϷ��)�}D��D@�Ӧ>#b��yъ�>�P�¿��H��̰��J��&t
�EZjSFğ0��D�F���w�06͢w��N����\ڈ쨩�*�5���k_�ԒG_�=�Ѥ<=���p.*����Z��M���~�����?�m�Iɰ�5q@Ҍ���bt������Q}�H�X'�&A��nQ��,��X��>���)Zi8E��8��WB�?>�Ґ�y��1�7���y�܁Cc ��0ڪv<��Ft�g�����aR�핁�.G:[��g�A�sҩ��:뿌����T���R^�c��٩]$��@����b�;�ٛ����t��sG�� >M��ac��������G	�.W�aM��u�.���+HU]s�A����6�P�w��C]�VkΝ�WA���B��u���'��k�,��xQ*^���|
h�G�r=��Um4	++/�K�� ����65��8�~��PȤ�M��Y�C��0	3�m�x�׊��M*h��͍�F��n*�)_�#���V����a�Y��A/��ߍSu}L_�.�#��3�(a�
2�+��d�O�n�  7����+5�oj!�������1��aɧ8=sP�W�	�� )���۩�i�:���§o��A�6���I>� �wS�V{�m�GUt��	z��gk�*>��i�[�Tp	���B�y�%��;-[r�x�wQ��+��5�x��$�gG��,q�mXm.�L�
��%�db
հ
�;�I�1B���[��.�����>���ܼV#�����h|J�$����q
B,F��B^�߿b�WˀT,�ϫ�xUE:����K�HL�Hw��/�?G�*�y#�4�!��H��Y7g�Q�`&mj��@���&M��3��g����*܅�W�g"��'�|c��$�7soȳ5�R��\��'$�o+��/���v���׿|�����[���[Mnd��J��O��!��Y�-�د�E�����0�_�s�

�񒦢����w̢0w�r�S^�VҾy���7`��xځI�!&�C�|�y���Mb#y���� ��b\�;r뫒O��=��/��*_�Y�au���RlYb�\uX8�T\��sr����]0~��Y-��>��W'KM��5*o���=��<��l�r�bTh�}&���v-BB�ݫ���T�[��N�hT�Z"x]C��LI�ap[��4�{J�]�G�/ ����؂s��87�����6���z�%Ae�|n�̳�+�����tqG��{��Cufr�P�W�O��O� `�w�l�6��CS�u��� �ZVy�}6�k�'4:Q�F���Ԡ�/�O�~�Q|�;�mB�+D�F��43���أ	.���+e�c#�.�.,�X��ʡo�����
�zq[��"�C�f��Ky���u��,D���ڔ#�a�
ϙ,*��Sv�WG�@�5� ��w�N�Y���O9oʿ׭-��%lDe9RD1([�F ʚNV뇥���!����Ӗ�' �*k�T��)�}�̯p��7<�ϘǮ�j���"ĝ�T���R� M:�/c�plZ��a������g�ƷǱ0�9���/�)|�PKY"]��@�rY�@��H�:Ĉ�
3LWëK�Ȁ���7��D��aI
"�������\W��hύ-�xSA���ƃi����}�h_����x��h�.+�sOҸ�;��r1�sI��߀��41�V�d��|렅�(t�Ph��s�q�R�R�M�� sC1��(޶���3=��GD�ٵ��ZG#��L[0I$eB:g�ȒҩC/X�3��5�qV���!�m���~m
�)�us��'��
'���a����m��Z�v�R�����
}�5�n��T���ڭ�7h��H͚8Zj��l�v�.�`��:��<Tl��N�qHOTw:jN�ZF�kqh�XowW��[-���cam/i"�U�/�5/���&�J;�S�����s�cU\/��n����#\{5L����:5���,S�O�$����K�?Q�d��L��"?�n���%ru�eO��魌	�#*���;�k�ށ���7�I��;��7ߺl��dm��;�� �P�_�#��S+����۝<�<DGXЎ�6Jo���9���}�_,��1S�@�6G9c�adAa�v�J�ɩXJ���Wp'�����LD^y���9��,��pm�s|W�JI�`RjDQ���b�?0URX�
�Qs!���������%.B06��Zh�w��Mɠ����*o�X�+�WZ�M¿N��c��{9@�2oj���c�����EV���8 �)R��|6Ʌ�m�L��],[��rW6�mj.�އ����p@������g�]�Q��(��� �[�.���)gK� C$���-@��+�A7ES�J�ħ�Ӯ
ޤ'�_��P�U�+�cd,��ZU�sy!ך�٪����~�����scxU��84MƓ��rP���i�Z�rg�i�,0��,	=�t��� R�ԵQ�{��$u��s���1��$�\ya�O�����kSV�=�����g�nUڟ����=@��m��<~�~�� ��~&/A�8
q���X�O���9GΪA���XXx��w���<h��Q�Clw�0�k۾v ��i'�>���Mr���4	�����C�E�NRl"
�!�}�E�8jic�on�L�à%���l����%	��� xפT�1�:"���z�� ,H�av���\�1�w*+:�������4'�ƥ�1���	�r�RHz�G)f���J�;�+EV;��TJW�ДX�@2tǻf��'���k�o���D.��T��9ި\?́���]�Pf��p��1>^l�i����]P{"��q�b,��[�K��'6�s���A�@����E�>��a(aZ��:T ��bD�<]b¼�뀕�� T�	��%���XA3�D�O�՜�����[��q��5�i{(�q�B9���:���YaYP^3��w�۹B�j3�+l��(O�'��Fu}�s�&Dy��~B]t�����ؒ��+8H����"��5��G+�Ҫ�O��-�c��}F�.�U�e�O�6{�`��,�%��o�X/\A�O柱ju��V�ȿ-.��ݾ�������cI�O�}�����[n���>A�Rn8��t��b�S`�Jʷܶ�L����G.ډ ���	�������Ƿ�v2ߛ<�JS�S��N���Dr� E�N�똸e��\�I~|x����K���;�ş�H-w���kg$�N�;�4��ްa�6�I�zE����mHUHe�M��W'�<q7�2�ht���uށ kun&�ge(՗E*��j�)Oָ�1 �}(_�|ũ($�.��D����q�����b:��jT���<�;
r��U<���̖Q�xK<�5p@�(�\\}6�%GT5�����C��x�}֟����k��R|"(X@{��m�>�4Ǳ�#5���E�tn\�La����a���9ô$������!|��Ԧ?��˙;t1����C�b��	i	C[6FxȢUxr���M�� Z%�D��?I�;�/)~i���Ed9�ri�`�I���3�Q|��T�,m��>�^k��3i��?!�ϵ�����%#�l����Ǝ���0N�_k�"г��f��
�F&N�z�B��p_:h��!Q���m�D1A�x�e��/��꫘*\b��l$l�5�[m�$T��
z��&q���9I"�d��>�7*5�&��G(���A��bt��1���*��u}�*Ҋ��P�ZQʹ�����R��f��:j8:Q�Ѡ�;��5�+%����d09���c�F�Z2~�������j-�ly5,##�f�(U�+�,��Q��QP��z����g@�� h�hm���"�e�"���7�Kq�d��'E���\�г���ﯚ�Zfq��Ѩ	�(����R�T�*��/��x�3)����8���۾}�ֺu�_&��~�88iyd��� $��6ިCLQ�����"4�R�9�F-�[�R�}���m��f�/od��R!N4C�hIi�pT����6G1�-��s��<>D��c�Vs��G����V��mՙ�Y\�`���]�D�h�2��D>*jpٜ�GѶ�m,�ᖚ	�\H,y��j��gM>��|FJM���!���P5T8�Z��[k�K<@ߚj�8��!f+S�����Zk��|/�l&t�rW�\?�� �O�a�֡���vI.�n��'#	�4
�3�a�k�+$2���p�О�(���}��=U?�P��G�e��������<`g}��nw�+"�$� �낻�n�+e=��q���y
;{���9��C۸�1��Q�V��rŀy�s��9/���KB����j�~���uì"�C��řD��8����ܪ�� ?�T�y�ߞ(�F�=\��eUu ���l�����O��/����ݬ1���Q�r���b��f��ts��A6����M�"j�oi}2`�F5���I�p���D����T�7U�T��)�pq�V��4NS�1p�.�R`�cy�GIm��G8"Յ6Z�ʚE�'oE��	����%����r���*0�l!�W�����)8����Ư�=�_??������3�ٷw��Dd��k,��S����/�!�ڎ�%:�*BUr��ܴz�RօD�Z�u[�_��BIiA���ٖ�|߇G9j��7+�� ����9��E�i��Lk��("8i��Gݐw �99	���5!�H&���kj@�iEM�.\�X��ٍ�q�����Ⱦ�
d����
��u�����V��#6y�d�i��LR��~������qJA�B;�!՗EB�@X������p������5�m�οH8�i�'�=g�ǔ�%n���i�%�t��:Y�E�/�pa.�[*U����E�?�:���D�������d�1I$�L��Dţt1 ���T�F�c�]����U�T���%��-2��hs�7��Q��O:+��~�a�P���O� .����r�*�?������������+�9���.���+^.z;<y�x�c�s��Ó�v&o�/��6�8�UO�2��=9vJ��.G�]�>�kGn�����>�l�ǈ)EO��(bl����-4�B��<[�a؁�+�IK���El�n4�_�ȇ�w�7���4ۯ�	�θ*qM�ǍD�d1+S�Z�/52��]�'�_�;��G��/v�K�H�e���9P��S��l��z�h;��3��z��)��KY_�Ѵ�{��_�ƅp�9A�Ct�����Ų�"��Ry����E�0�f`�~{��b���
r��
����1�|�;�����zkn*x��h���Q�$տ���5�`���L��T�,��$I;""MB�L�����{�ct׎�xM�Ck�ݰ��;8�拓��0��x�1M��0�u�����T�}g.D~k�}��Q���Q�<�^���A�c[��-S�I��=?h���Ҫ�Z��m�F�|P��GP$y@.%_�/
.T ��hvʤr>FSdF�m��$-�����2N`�[r��l��Ǩ�B�,`��Aw������@E�p�A�s����9L��Q����IGQ�@v�C�&���!u���Y.��S�A��_�ֶ� ;�<(T��`:�l��� �d ����,�w�4��+��u�������bc��yVF�CJ�:�0��LE$�aD�+Ѧ��
��om~��!:�5M�v�4�嗍N��h��ʋ1H�.<�Q�,�� ڐ��"�1��K��|���N<"Z0n�-�h��a@��F�� �5�XA+@F��2�jrt���يѬ�	�����<��O��ف������vB��􃽜�~"��-�`WO�5�CR_��f��x�����!�l�ݑ�9�2��>�f�jB���?\~�!<��9޹5�� ~Vl⡞�X�d�+Y�U�"O#�V!��<1q�N��!��!�����	� y���+��䨗9�LY&���9��WӉV�J+�O��"l˲�ȶ?5U��;f.�t���
�%`�����l��iX������9SW��7���w�+p�]��<0��t"5|�맷�}�=��M�oo�����] \��jqj��<����,1J���G�v����]����CoA���Y��prRO�r��.k+0�,�tz3=��ئ!7��ztK*����&Ǌ��ZԊ�K��{@�����\�|c��pf����b	��ߌ��Ug�q�S�7�!-�R��H�E��8��Њ��FtD]��=V�k�DN�d�(ϓ�N�-4J=���@g?�_�.�UC��.��`�sB`��)x��z����>� [�,9~o=�z�d�K����m�gv绗�a^���S�԰ulD�.�(�XsOvJ� �`�k�8 �F���9R�y��@����.�z~�ҵ)P����n�@LC�~ !�EF`{0kY��g�~�X%af�8����d�0 �-D�NR)��؞I����Φb���0Fl�}*88uu���vY��n���pD�M�"�g$V��O��0����&���(����D<��ӒV���%V$9�q�b?a���u�Kς���K���F�=0Pj�f�k�[=����}Z��w��(S��^P�gW���rY���z�.-Z	�r�Ӥ�����c �|L}{��O�v=vn��c��6-j��������q���qkȦ@�����yy��6��Y� 9�֢u�G��-��ả�?QL�޸�!��@Hl�F	�#��zKFc_�;��ڛ}ɦV5��o�?�W�4W8���V�d�l�P}�-��Y-*}��L6]ɹ.~Q!r�W�P8_L��]ʁ�g�!s<ܥ����(H���h1�ϩw��(P���>�=۬(j.��Bv�5p#� � /~�6%��T����Z
;柘>�e/�H���G,����<WQ��-����C���ޘMv@ZU@��
C��ޡ�S0͇�\V��Er,y��{`��)����>������B�	(M.��
*V݋R�4������m�~��i7�u���Q����N�r�ozKdI�{O=Z�����~jyo��ź�
>��d~?�����k�lC.��@�XS��'��Yz�I$��&��F��	B�m,Q�n�!��]�����I���I��٩
]�󪫧��i���:S��c����k��D�����+�N�_wd���	�#ً�4p�5�`��⮾�t&O����7ae![��c��|��7��:Np��V�o7�
	5��(>���V�qU<�i}axf��H�}W�l� G�U���o����������4�RR��B��;h�; F�=c�.]=�S�X�fe!��E�=��`�ah����bUD�@<�-IPqZ�C[���&�A�U	riʀ������$%�ogu�E7lf�w*%��rte�NZO�'�6��Te���fG�r�__+��%���ab�b�!�>
o�E>k�i]Je�Lj�%V�x��Ɯ��48���y.���5BSoJ!�*+P���n.7��pp=�#p��mW��=�;}>tcR�.��;v*�g*��z�2���,����;�_e�nl#W��2PR�tx��-,C�%�O�*>��\�+W�1��`��C��&G���6�IK�;\��3���{:�>�
��:�NZ�0�����B�O�I���<��JM��M����"��j�}4�E��5k(�ٵj�ɔX�5c�d�k~�_s+U��	t��ז���C��]/��Z ��[<G��tr��+�!��~��lZ�uF
dq��\ '>	�T[g��E�sM!���G%(X1��.]�d��ഇ�9���(8^�I��X��eA%7�: /����
H~��K�pS��F�5|�o�y���f2}��h/C7V9�j&@��5�~{V�l��XP�p��[^������E�@\S�B�F�����
4Z����!v����`r0H}�2V��5���	���`�oW-[�Q>ꕨ�a�ho���ZNu��.��H���{�3����3�]#�g}��)<2$�~��۩Y��p����x��E)���|/~2|8��ʢ㍁p�B���E+�>�� zjJ�,�G�4��1M���m���T�c���'	u"�6� �?^����o��$�d�ñ���51��-,ө�6���a��]w�$�`���ڒ���g"�7#I�͌˸��>]E�N�����R��H�q�u�����7
�p����Qc�Fѿ��D91�A*8L���e�o�+e���c�l"������.n�ŝK�}q�Ɓ�=i`�U*j�
us� ?��)ZIs\1�x�c���}����e���ɬ/%�b��`��`9Dk?W����,���v�@��m�ts,F'��u
Fz��Ɲܩ.{�=���A2(���6�����y;�"TZi��=������o˧ۥ���&Y��x$/��>�P�P��헵>��lڞ6�䌆�g8���'��7b�Z�ӓsǽ����삆��S��������I�y��x�Y�����F9�g��Y |�������.��<_|~��R��������ފ��q�8�$V�+��^6|�l��J�z���@J�
���iU�}�VDM��aOuz��v-����51ؾpm�<~)���3(\:��
JPS>��z�E0��6�b�]aIλ�0!�#J�L�([�h�^$[����O|�R��A���{�-�v��!�V�������?j�/�ӡ��m���ۓ���A+����������b�~ %��1.�nEL���K����S}�"�7yDY+t{Lʮʾ�}+���Q��Q���{&f=W�xJ�R�"���cv� f�����D�2\xԙyX��	�%�pJ�+n�[O����"hwZ�ߵ�dH���^��Aǝ�`��Zm;,dig1�����K+V�7�d�o΀��v.�?�A�5ryM��j�#�9I	{��/�_J�b�o����Sv�k�i |� �)�SrT��/^�"�����*�>��B���O��40�������X��8��"�{rrBm�����v�$gQ�K%�S���ά�gޔ��4b�+�I�Q"�o�45�{�U�âo� ��)שf��fFZ��ޯY�V�}n`����)��>%���uC(8�u�wX��ĭD�ړ@y���WErMA��P��F��U�,����3�\����a�������lNo�� �䪆����y�<&Xy��dVN8.5`��P�!�=��r����'�[�[t+_(�+�	j�s��TD�:f�ʏ��S�)Yze�G5�>�\�y;}�
v؛�d���T�����[��ȡ,�����0�7E"��39/>j	���H�s�C�q�.Y�?GFt��8�2�u9Hx�H6,$\זO�ü�:�����PE��TPm�:���X�*�o}P�ԜW����s����k�т�y�x疫C�O/�h��t�H��y�ڴg��Z�-�N������uvl�/|��� ��9V�Z��$��5�a����X��ʀ�,��CօŢx�q�,��|�'�6����7�X\�+nO�A�y7>g�dHqlh��h��B��-���U9�h/L!P���Y�kW�����~ �h��V�l�#�W�X�4`��g�ۣ{2}�����\	�[�Vs�xμĦ�B���s����8e��Ϥ��v��{>zz�L�ţ��Fk�اu����g~S���=����8߿L_�J�6�0um):���W)�we\�%��B��*O����DU�R�ۆ�E����ԃ(ˣ�vC�ePnU�w�R���u���l����f�ƘP�	��2��]*�,��=|�������7X�ʷ�M� *݁���	.	iұw+d��83?���S���s}�]@���=�Xi� ,���d��#"d�������G����ɂ1[���>7�-�s�N��|��f��]I�XQ����4�+e0�<CB|z�'ؤ$��[����^�ɰ ����-�T�F���H���q�FK�:[Q��v�wP2e4��0.�^$k���v�t=��Eq&7$Z�R��u��T�'���덡�Ky3����2�Һ -`&#�:�w��@�o�u@��Y��`���	I��/�"�EX�� '�=�� B���'�\)F�m�V��}�S-��oF�a��$��[-���&m8�	�~���q)�>r��8ipB|�_��1��B���h�Ƶ�����Qvs�&o�ƺ�6�Se%�.�2Lq�J�b³�b%�w���H˞<4�MȔi��2�-�
ۄ�G[t�6��Ѷ)��j ~��;";v]M�sM�10d���jOR�������ǥ���>6h��v]}���Ky�����V�2`�+�d�$k]/���Λ��;"��t��`^�q�����C8���v�bm�*~(���Y7k-�Z�S#k�Qr��[,P�z`h5��s�n\ތs�p�n|����V�Vo��r�%3�W��ؠ#(W��?���Z�K���A�.���j/�Ƕ�wPL�S���B�U}�f=�Ln}�f�bu�������]�#5�	��H:��� �i�{�co����˼qOot��Y�ߔ�:
�,z�Y��2�. ?R�6ͦ����u�a�~�z�)��ɿ&��}jY�x�Hg�ؚCȆW0\~E>w���ʓ4�*t6��ד�TF�TKٰ/���^������������b��4�������/��V.�j��f�QK��^`Dj����L�5�|�\,�&�?�?�q:�(,�����B�y�fI-�;kW'R��5 �^l� e��%�{G�x�Em!O���+�W0ǀ6h�GA���6�Z]F�"ƅF�-���E�R	���u��5�^�jۭ���.�& ��� �x|�(x]t�]ԪG�w��6�\=��r��Y�}0���ڵRC7����-� @x��#������^����grҼHh� 0_�l^����7~r���9{a�7x1��ϕe�!�KC?C������i�E�>�0��C�����	�I�E��AwC����z��pu9&(����K���a�E�Hĭ���oUtWF2�=��=nF�+���n4��q�l�-��{�BO�*�6����u����\���UqRFlT�Yٲ��eᄦBһ\`Q/TĪ(O�QI�!�͆�S�;�����g���p��풉r7���Y�*���PO����[xe�w��5	&c���DՐ�b�S*�7 ���lw�؉����c,(B�p�`B�!�����ʺɹ��J������Plm6{���2JB;�#L�V.!��y~m
��w�^��#b��-���x���>M�5'[��m}^��s�VR�r�:���d$�x�s�Kz�>�g�%�,�\�l%�)y	�T��f�Xg}A���p�ք�J1E����*�I�B�C��H4�'1��AZO7vg6�|����݂�1h�ޑ��{Z˴��BUnV�9��Tc�a��"� I�lY֨�`�/�����u=���p�T0��J��`�^���ؓ�2�큛=�����{i��|��G�AG�Tp<|l�͊5�.J�����dP�@��$k�8��9��>�p�>�IM���}lyP�)���2t��Hc��6�#+�U�@�5�i}��I�B����!#�H�
�"$ט ��Ơmƶ9���L����$��9�����`��9�k�z~�^o�n�G��߿bU�q�]X�삿RC-�84�v����I� ��Zn�`��4�EƏ�3�7&,��9k9ߢr)s�:�J'č�JT!�e�ÕV�tJz0lz/�R�(X�SH��JQ���k�8K'�d��
��rHe~(�g�h����gJE'oN�2��W,#% �n�w���a�Saa+�D�iE����2�肮KV���Mv"�|jl��s�J��ڌ�m޿� G�/j��=��+��c{\���SSsY�m��� �i�����e�ؘ<��]D��#]ң@92)��Ǡ��~<@��+Y}��7�[i�A��ں_�D��4�%#��J ��:�o��y��+CyĂXڶ0`��U�����(Z6�e��9����lB`b'�\jYcO�*󙓮R���B@����3��&�%�^���r~D��֞�&i�����&gY�����l(��)ۖ�"jj���z�)�F�N�Z��IYQ������WPcr@F�.�O&�#c��3����u�t�#��9^��v�,8Ok�:"@����s�ɱ������'g��;.�ߚ�X0�Q\���K~�;[�A`�ճBDU6*n��\�gdK��1Kbxij]��Q�@&Y����nx�ī� ���a�v���ZN�>����9����KC��x��+{�e�I����X�����B�<��#2<�)��b�����ԕdC�I�3b�����K�M>�ME�-}, '1;�\v��D�~L2�FYF��H'��8y��P��R�O�o�yx�kh�Š�h)�<����
�h��9u���*���~��D��ȸ��������W'A~o9�ä�|�,���29.�5�)�WA��R��Ͼ�ߢs͕1j'Oլ�����N�Q �	��B�6��2���X68i�tո}]���B����j�h:+!r�:,h�6�Qo��8��@ ��Z�un+����3�`"43�+&��Mp��v�Y�g`s��Id!����g],<^�t���yA�C04�}�dx�U��Y0��DPv|�҇�LF�ܵ}n�3�Ӱɶs�@d!�F�'�h���[��wM�nɉ�3zIV�4nBX�Y�x\��]�+�I��A)�A�SMby�h�M�<��R�'u�(W��d��������7�#���Zw���J-�<�	��}��<��� �7?�����ݟq��Lxz�|�y��~����)1qa��A�6C�v��6�����z9n�W�_�U�.̢��OZ!���ڻ^#a��S�=�1�E��r����nP�	 ��͟3��������o�#<&Ƌ��â�2�q!�Y���k�,4/���eO�%��Q��p�R]����Tu��:
���m��N�io�?�FN�S+�U�W�{�*��R�����n&o�mwq~�j
� ���UeN�4�>C��%�L�:�Cm�v�V��{���<��Q���U g[-� ��� R�����Y����t�<}��pqE�|��R�9�T��hNdж���ѽd��������� �l��	�#�$�Nҥ��&�w6��"��<x����n������u�<��׫Uݭ�r��i�@�}(Ԗta�ѣ�V2�Y��j�_�I��I��G��H�"�7�{ Te���&���N/IZh����%(��3�9��]�F"c�Z��ezP�ǥu��@��wpZc`i���Vտ������'l���n�������%��N�l���q��*�~Y�ʄB�c9��R���oŴ��}�.�����b�W}0���K�p���J���W����=ъ�"R�І&g}��o���������L^ ~ ]� �7c�G����a8�rVr���n�)9ө�}����!B�G�*�m���i�+�4�s�حP!M�J���w�Ao�Vq/�k>>q�1����_V��Ƚ���6
���q���8ɡ���g�x� �X�U� s�/��:�N�"?6�~��Bs�U�f_�q�+�S��E���(�&H�AܛCm���^�Q�s�N�Q#_	�"��y;)/�ݴh�ve�5�R�0;i�s�~og	"܈\y6^���Z��J���2b8��N���N��Y6۾��$"^�K��5I8h�E��D_c�$#W�^���z�`#=L�#7WF*�Y�I����7)�J�b�S��=(U�W�s��9�:�r�?�A�p8Z�A>�=G���ElWng:�l����!S��!�\�?�A�������ڐr�Y�"y��&^rW��$�QƳ�=-�(��gS
�$��5uA֙����j����޼�d_Wk7q �=K8q�R����>��a9���pV�����Pz���ZR���wV)AN�l�V�D_غV.�낏j"���ƄP����V��l��5���NXz^#(~!W=g���g$N��>f��ہ؏D-�e.�<�I{�5m�W�r��r$D�[s8r#���t���p�℺��!(�m�s�����͖�L��[��RE����9�RE�<���Ɖ�$�y��T��y�ǝ����tw4.sebᑤ�%�S+[v�$$�vJ���*הe���o���aT`=Y(��1�㲦�wpS�;�|��Xg�V�#�}W��׸��],��Q�/{�x�r�҅_�l#�Q{�(�V�2�f��S&,��)�d<�����ʔ�eO�w���8�ܡ|����6�$$�s�B���̧�9����go+	gW��w���C���F��.�_�A��f��`�jw�O�,�@�(Ĉ���囦Y�X�(]Y Z֙�Fy��KJg��E�U˒Ek�������wc!�b����ݜO�ՉF�yE��'c��I���$C�JՑ+���V��C��E[�Na(y����v���f<���C4��lB[�ǐ�S���3a�If\�� ��P��JcLb�(�q���e�xRI�3�&Vr�����
C��D���W8����v:4���~����!�\΁&�W!���<�5�sv�Q!�+��>ֳ�f��'�g��ZyD@�xb�D0ZgQ_�������7�L�iie��c,�f2i�-����������S)S����9s�{<F�j��}�r+�����~�X�e��������	gF���ʊ�-�!T&��1���iw��z�o=6�֕�3ɕ;H�u��`ܶ�]���}�o\�CⰧ�&�� ,�)*g�B�&
�m�es{�V2Y�R!_6����6y0Q�R4ޤ�y��r��h;�U��L(�UÒ"���S��uo�Q�P���L���/ %�}��ђ8+��Vk������L�k)�?������$�&��� cF�$�R�m�
���=�=.~�io�sL�vUw�����&	�m(�O��J�UhL�n�Z�Z^��W�"�^-�Ը*BtR����x~k�V�b+�@}GJ�h�"ωh��f�%���#���8��"eq���!c�
e( !�P��W�De��J�J�p����j�]Up�2g�+~&׌� _+���ʽTQ�79Q	Ek�UK����0��¸u}ƙ�)�̰�3��+�"�aq�&Ĵ����Oh��#��n�9�2.�O�,�^��:(sn�#�}#]�4J���"�z�9����H$X�aASBR��3��0 ����S�;�ۈړ�kwI�I�S�}���WT���оPo^�"��N�y(x���ًA
�x&����ע�r� [=4��g�:TABWp��.|�	���l��Li�	�;ɵ�����T�a�F`��`qi��*P�ԃP�����ْ���ݶu뙹�OB�b�A��܏$`U!M��ȁ��p7�Sȡl�÷Q��7���,�޹�"�� D��E���}���V�s܇�d^6�&����*�{}٧;����[�&!�Ӛ��~]�s�P
��Wv���N�o��+`�]�#*W2�d�E�j�ɮ,��K% ype�&�2���]M���KRS���H��<��2y��y��fC!Fk$�UrS'G-hL�^���������]������_��1��~�K��� @�R������:7���s������S��wqe6?��>:��V�f}�s�']��wa���
Z��.�Rw"���a��T�S�F���?��K�) ��� F"UtҏГ�_�(G�LՉ�	8����4�+�G*�/�|����~%=ꏮ©��in�/<�N[K+:V?#���S-2,kM��:
]����OC��fX͙� 361M��ݘ�::�%��q����J@�!>�SV8�J%�(�&>��ڪ-���RM�o��cA��q1-��o�ir���Ws�D��8P��$'D`x#&w��ɖ��~�Qv0�	ec@v}��8��I��W������^�!Vd0�3�>��ZS�%N�6����%��|��.H�p3V����w���9����Q���伮�w��
3�����n��Ƌ������iؖ��ǐ���9��=�8h�}X��p��r��n��,w仞%�pf*~��Q�8�IXXP�W��u�+8���>���2d��I�~r�(��P�6+�i�� �ܿllv����H�4@J3_ݫUi@9���v5�dA����5h�nG�jeu�pb�P�dl\���h��P�װ�.�_E�e� ;�R@?��V�P�_.�������Im����}H��$Z�u]��A028~�	}9��S7hm=q�0r�(��������COأE�o%�N��1y�����)� ܿ�K���.?��(�?;9�!6<)�!��bQ���Z���p��.@

����J��ڑ�,:әQZ�p�T�h��U�>E�����y�{.1lK�zi6��	^�2w�0[�&�S#����m`�:l 2}9(�V��2�>���F�Sp�QS*�V�z�7��|���˚ -�2�	�<g�66ag��E�ݜV�/Hg;�P�eAȬ�<��{�6#��?�Da�gQ��}�Fe�b3o^�)�1R(9	ϓ�Qx�y� �_�LIG]�
n�u�zaZ��Hx����2{xG�� T��k��c��@>��O�� �$�/���f�K�����Y��H�\._0�No�2 ��@�TZS�Ѫf��u���v��.�TS�����F�R#H^E�����(U�a��<{ި-\�n�Y.]Ȱ���A�/+k�5�:ɰ�ַ9�J�}�v�ō���[|��g�E�D�x6؝��[���c�`1ѩ�L�,�$��4�L�4m��]�����K�G ���� ����w�+g��Nr�T닣�b���O�������3���Qd����-�_4�ӯV�V"[/ 9X�zP�����9�wM:�:��_;��f�@�������s\���*��|���C�'�Nx����_���'����rw�UH]"y�c���.4�iz��B!�ȷ<���%x�*�|a���[��`�>k�j�]!������>���Q�1�Ba�ɷ�&y
��i/׭������-�A$#�,;kP�L{f��d�'mc�,�c�|�RD�/�c�N�$vDe�H�rm��k��dJ�'�I%�	3�����-�w~j�B����x�j� �V��X�c�孌�l��c�Ӟ�LM�̅o������۹��K�Q�`�,��]h��&�A�/�:ĪUo)�B|�=aa��ܙH��e����h�f��%�k�>(tX���W��p(�'-IS:�������z��e���@�̑ߪ՞
̅�w��8]+ǵ;�crEY�R:c�!�"J3R�7��z��#X�=;%���y�m �hD���V*Z���Ԅ̀�͈�Z�>�yb�����	�-�<�F(F����~�H�i�����v|WEq�@��;N]��05cH�s62fQ~��d�����-���R�n��mfA!T�;g"}�2?4�_��z�?������*����-�ӑ��U�������ٵ�ö�d�#�	VAà�T�/���x�p�V����.o_9I�ƌ��,%�@�@%Epx��r��ڧ(wv�4+��ꪞ"��ׁ�<����ׇ����W�����Ѣ�c���c�Rh¤�q����`|A��ʛ�����]�P�^XT����E�B�̝���F�9\Ķ��.�E!�w�;���̑*]�����6T��~����r��C{ũ���e\��i�C�>�|�''�y���z�2�FM�T0�dq8�nx9yFdϝR	q��x�,q+�9c��TYS$��}�(�h�ߧ�iܼiiQ+"g�B��[��S�@v"�����=AP�� �w�Ys�^G'�� Ǜ�/!�8͊ͮ�'Y�Bpm�|���~���(�Mw��%�[�ө6��0�T5���	D)a��Ai05��a��3��a��;L�P���heW��&�����-�-d}�N(>~3��,�#^�Wtal�<���5�w��@��1(S51��Ӣ�@9?��DѶ�a��M]�V��o,�vA��w��Fz�2��:�����WʕnJ��Ag��Vy�cR������֌d�/w?)y��}�]w�C'N�{��so���4m-o�ӭ?-x�(�kB�NB���(�H��|5���^��xG�R�*�V�ɭ�����m�gH@�l�~�U},����>��W����;��#gPj���u�����r��@�e�	�8�WXj�b}�V,��EEU�������[���#?-�Xƶv����Yӭ{e��F��j�|��ԁ�@�"(���W,�'����k7m3.4~i�LIZ1+�x� �[�5 �h,�X��h�9�@ԫ*lGr�\�LR*B?��߻��g���
�e���Y��hy���/���\�)(zJ�*�|��si�`��;�E?B`�Ҳ@���	���7rJ��O1�<sҸ��7�� .W`$�V>~���d��~��;^���VV�K�s���j���Wbń��W߸�����:��{L��gL�z��WN���"J&��֮�pyBQ��f>�hb�)��<��O�d��� 峞@���G�?"����:�;����������c9Kr5�OȲ��Kr��g�t[r�Z���tgfڪ�ء�B�9Ϡm�XS�OJ>�%4�^�'���V2��B3B��~�Lv�E�}!���-y~��R}�I!��w�u,6ݱg�+}zY7<5�&�,��\��!��k����ʰ!QX�3���d3CY�h	�َ,A3�X�d.?t���ɰ`���% ���:<K��L���Lg�SQJ�(I:�_�Ud����.�u��v��]��\�b�-�@be28��86�P���ԚE�7SrN�Y�`Qc:(}�?�����,��]���&���^��	[�∫�r)ʆX��-u��(��;�b��\l���5�X��?�m�Tw�D<�x"KTc6��`GS��0�Ե!�K�_�^�rT.Ci+�%V�X�[c�v�|�6^ˁ�O���`��ɲH����I����-���[����@��EM|q�x�փv`�8	)��<�(�	UG�!<��/)�F���CG�a>[c=���\jS��(�Tm��CR'2b8/��!N�"ֿ������IW�Ͷ�jT��۫b����_��Z/�_"�N۪��K�g��ڻ���=�
�fާ�OpH�g��b�)� KE�r���l1dȮ��b	v����0�u�(^Wvrb��K�,%��t�g�)\�]l��dtO�����d��]42g�_ĶƷ#[��;�]��|*�\,$IsqyF�$B/�t�P�M���|�~_�����+=5GY��%���JXA�?F�[�e6:�\\�V{��à��*��xd����J��(��EW *M�&c;Av㴁�	>d�M��������8r�����<�/���m_9�ʩ�$���/��Z� ���`0×q<�r�א M�[>����R �6h,���&�^S��>�y���X�{��߇�%p=�T��Wʕ{*� ��ȸt��33Bɯ�+� �ws߲�cN��ђ  /�=/��u3 : ��0�=�����ߤ
���=�1���F�B��~���A��~�3��
 �=�4.�[ ��z�35���I]'�2W]Dc��
����Gd�%?�<�� �̿��������^ˁ	j�/��$�|=��m�'O7[%�Z��E�IH�J�0/���0^��3� ���"���w�	��8y��'[�[�5�Ytޢ���D5!?�8�j�K���8{���+��$���]w���Ƭ|���vӒ�u�*�q�q�u�.o<SIH�b��>Lbئ�}�˴$M��s傳RǞ�(@\�x	��tI�t$��*�%��f�=�� O态��G���0� |1�/��!�a+ʩ�E��G�;Tr���27a�@=/���Eo֗i���|30wx��\�-��|���!��� F���0˴�x�7�x���@!z��$0J�s���T�8;w�Z/�I-��&6 �����jPgid�!�hu���;�N切&�C�H�2�5b	�^��w�C�I��	���W�E�L�M�֧�F}�k9�%<�Z�w	�Yi �׼.�8�І�7��s��3d�CF��\Ӂl���m��*�~BaT��؄����.8L�*!R�o���K�9],����6Ԃ՚���z�y�ma�1i\(���+>�38�>�f�v˥iltІUf��`(�9�W\��6|C5����Lľ@;�s$�
��� o
'�Y�X��s&,�ș��6
���p}U�1�A���b��W�s+�:�#BŪ������O��)Q[����H1{�i�03N�.c.�eDx7R0Fxv�?qzo4Z�
Ѵ�N�T
�t����H��~W�!n�R�
B*؁�C=Z��:���P^�gS݈�$��K�c�s��"җ��d���O�:��_���I�ݬ�R�.�-�������G٩�I-�؃�it6�x"�9��]�j�;���4��,"dmT��3Ga��r�$��t~S����&8��Į�<Ԉ��x?�8�,��lN�K2AN��}=7�r%�?L�u�v9�;>n9�^�8�Q��N�z��g-����e�n�e��������`�����4��>�*Zs��
#Hh�ק�J^���oTX�툏.�*�k��9�.��v'F �LO�.:S��jħ�'4�]k��\}���L$X=�����x�P��(�R!���M)��|�v+!�>���ۂ��Ц
)dQ���U_%�:H��V[Yə#|D �U���H����.O�XYǨ���3����W59���|b�J�1��*¢s`Q��E1�@�!f�K�/���L��M�8.�9��j{� ũbR��b�Lgm��r��6Q��+���U����������g�ڈw�4�v�z AF����n�ڢ����]���Nu�WI�\��m��d��"]���}|?��׽F\� ��c֠>��)E�m����OR�������,���o�Rtae{x �]_x�r��� |�h�.��z/?n��$R���C/��b=;�[@J�¼�kу�ׄ^v�I����Aj�X��uV���O"1v�|js��09M�w�gC[�d������ߐ�~ ���_�'��_+K�2�7j#�3(���IA3��(êux��V����6Z`��'�$�<��?�u��J�xfp����3$��~��ПLN�<Ï{ ��+JMM����i��*�94X{q�EL���g1W�2g'Y*���}��=
�׆K8�~��+T����ѹ��Rim<�=  �N@��l~��]�U�UL�����zC�v���/�|3i���1a�qu���� ��,3��J���fenn�춠�����9��ƍ�]p���7 ��	�f�+v����y8=�K vN'@	t��:D���H>Ȝ���0ƲRY^Tʣ�
�0�]��-�_�xc�2�����}�=K��O� !(��U���Lu%�w������Wh�0 ���rBE�X�S
��z�i���7b�۰q/}���$�
}D��L�K����8�L�{�h��a_f킣���~Q\�
�v���^��J(��J�{xm������1���燡B�ן:mE�����L�b
���e��@�י ���E8v�~���U�_ݴ��^Q����%:Հ����g���qPY���HZ"˝�_�����!�)�Db���WJ�'�Og�`���x9�p���:7�~�������#��e|�ų�#&DAx��~'"%�;#��560})����ͱ��a't��\9c��Ix�����VH��Tq.GT��}/W��7���|iOl嵎���9�WSR%��*Jt�:waU�E��泥Wl�%Z"e���*�L�S���0�@Z:�]L�4��i %\娾���R�*M&+�6Ďv����Y���3ra�nF�{"�)չ�]h<����a��N�9���9���3���$^����?>כ8�:�a��Ku��
&�a�b�!���� q���s2��k�0�a@�>�Ge9P��ZC=B��n�q�y
�x=D�� ��%��q�R���-xp U�G��mN��0R�\Y�:gyYu3��N훜g��-�ɑ�T�QZ\j&7n�����H{8���!>���г����t�%�5���w����TҞ{�n�KJz	7߹z�������6y��a���pPy����I]����������"?�v	H��̬�kse歵�&TWcB��]��86T���N��k�F&f��)X������
2;�%����F[���)7�ΰݍJ2���3�����3p�5����׏Oh��B����;�EK��j�0[l)�ٕ��f���
�����Nf%��t)Ҋ����R\c0��=  P����m���U��ʝ20�Q�t�t@� ����Drޤ���z�Oh��Ւ���V$�h�U,�=�D�x���y��w�d�U�"@!�p��˫I���
��ńZM�L|)�þ��P�DDN���&����ps�*���� �|���M��=� X�[���i�����9芦�M�P��2�3�VLv����M!N�G�u�9���I�&\q�sgl�m?_#�]�C�\+9�/�֐J�X��{��'>�h��F������*EL(�҈��`<���ו�9�]~܄��Q�q^n�|��׼�W�~O^</<��tm�X���񳨈%N*s��I�/|��Lp	��Gه:�'Ӝ^,��(���\s�!��J�*c��3��`_ ��;����k~���+��ӵe~��2�\��, IFwBL���.��K'IM'���fe�D�ID��@o��FbOEg��-�Ў�Gc�P,�
�IY�uj$2�k=�exZf��i�Ɓb���hЯ�b��*��"hX�~����-ZA��5?ybU��W�k�!d�%��,#�$ �������*w��\q]��,��m��X�0n}wF�C�C��XP� ʃڊN�
��Ъ��u;�:�^�IN����x�E���3.�2� 8#_ɔ�#�`�rf��lI嘂� _S�e<נ����;�o�1f��m��|oX���F�����B[�T6q4���8�Ŝas�#byw�����btƭ�H�lR��z�q�EJ�.ˉ:�W��M�����ɵ��=�zLґNU���̻M��g��"�G`o�)�K�A]��.�����N?�sG���	Y�_�K��&�c"��ƙ�!�?I0��`���EY�����L�rX��>Hmp�X��#X�4nr](���ac�w32�DM�b��Yd��(qh��e ��z4G���D�Z�4;$_ʘiJY7m%�-�M��tb�@���_?n"�d�iF����+�<�Җ�0�y&�5[��d�&��(2}���aT̟u�ao�lYg����ѐ\Lnd �K4\9lw{����7A�;��ƙ��+����R�d^r*����Bk W?fk�!c�1t*��@��I�GG!�PDpB�UDB��vp���2{�Z��K?-��f\��Hq�\1�ٴ\�U��c�+Z�v�Խ����X)��-���ջ�o���"���I�oJfcC�f�=�[V<�	=����bkF��0
w:�Q�z��>m��}�|������|o�\�YFD�`��J�wF�r�~�X��ޭdX�p��?�$�����E����`9պ{�985Q,�~n�j�쾶@a!�q4�	�.���Đ�5`�0����8��y���0�׊0A��Wݠ�r]�!���h��þp���I�X����Mf#QK%sp�2<$���*��s�U���E�EC��ZT��'ɱY�a�z�'��~v'Ƭ6�f!�[�!׈�o��x�5Dݘ�8v��ܻ�7�6�w%��9�j&�l(����=���D��&΃��[��Wv�����V���8v���'�u�\�%m[b���YŎM"�>
jR�٭�%>�Ӻ?O:����l�� ����@�dÍ������`�~ �pr�bH����q������e'�a~��S��Fe���m�Er�v\��ε�.R(��ɶ%9����k}Dߴ�!�]�Y�0��S%�5���j`xz����$@}v��m����.b�X�IA���:7���߾'���佥m92JX���,pbw�8�p�l�V�%��"����ÜKBz����<Ro�����AR���N�2 ��-|W�kU.�
v����z�X�\�؞@Ŷ�	~o����_S�z����y����i����`Qs��S,�`� 0�t���Te�J�Ŏ_�2��� �x��R}�=�Ƿ'9'��|���=iԋ緮ksk-FJ͵�m~	�($���ޓt6Ih.�Z�o�}�~h?���j������و�,�u�T؟�Xc`�؅�Ԓ�ҩ�U T���`��m�y�OX�=��Q�ئ��ud���\�5�1��"�y�7-��[�LG����L���?�O۫kg7�n��A1]a��/W�VD�[t�'��%V�@o�� ��&J��m�~��:$�Sv�%��%�r�d�y��8�;$��'%4mf`K~N{ב��.�K5tS^!��M���3�+C��4����;5�`��Ӏt���/lέx���6��w#�D��߇P4��SL�U��𿰃�t[�K�[�7w��O�?��$gl�.^P�2{���eZ���W�#�҇rs����4B�v�L{Mk���;�&�S��ο�[�с���@�����r�S����&.
�ڀ���7�\6ک-�
-�^����_��9����ŏ�i���?o���GY�w�z�u(��(S�f�@��Vq�^\gA�/�(e߈pR>����� �R�	VO|�HU�s�x5�
��}6��ewYy��˻N(���n)�B��}�?�\@c{�J	*��\q��̆hf9�j+�5�}�-�^�5���bN:�8��G*���<}��%�_��[#��[��pqzi��s�(���:��$�a��31��&-C���(��t�ؿ���L��]M�yCP�i����zސ��suQܥض���]�<�ہ31�- v��6)-��ߨ���L��η��x�Q[��3��(��Q\yɣ6s�"�[�u2�����]�M��R����K���1�{CAxB	��#�+�h!�ETJ��X�g(=�ŉM����
�I�\c�u�>LLz��$�&��|��m�0��#�>J�������vN/"nb�i�ol�Ռe��%"0�ߣӸJ����V�wӛ"�l�9�D���<O����� ������=�5�oV%���&5xs�+��	�
�p�ɚ,��O"#/s��V_�D��$7�}���`Nҋh��>����{�
�l8�!�����aߓ"�j�l�XS�PY�=��AC�{��/sE��ܽT����a��{?��'br�b�_�� l[��!�������Z��ץC�_l�*7�c9=P�c���p{y�	��e(�k��b,��t��A}��rFpF�v#��ow_�Ni/Al	+age!]�P�٤R���%Փ��2
r��-s���#��9�
I'���݊?LLU³Vh����nm12�S� r�й[�.�*ѪSO��P-\�N�X�<�8��W.����[N��1�8�Y��`2ʺgW�.��@v��I�>�bL�h������bفI�8�I"��9?�;wŸ�i:vT�ï�qx�=	]K[�*G���R�@}i68��x����z��;|�ygϢ�Y����eȓ*�)Y\<������>�)N/����E�Pb������m�f'|�^���-.���r,)(�͘@H�`�t��W(���F��q+��W�E�5(����TcD� ݬ%��݀���S���y��YY���H{��)2�PWU����O�U���^�o�������m��Sa��r����40�ƾ\Lm���Ϟ��X�&�5+�p�˞:�n�l6�ׂf	3�֧��b"��n)�����Ķ��IHU=J�-�����%0Q�S�f}JE�`-�l_�CՊM�`Atj����0������`�%�Z񥀠X!;��Q��,R�zܘ�dZ��q��Bq6veb������)����eX#֬�����u*�"XU�����0�Z�1�hb*,��H�{]���I�,��p�<�:�έӤ���Ģ/k���A�ъ8���6�H�#�1`]6>�y��-O�a��Q�nI5�%�1���*�X��d����۝Z�0j&���Уs����ʆr_�ipax�q���Nݯ��a)^�Z�x��!Tx;AUmv�(0ٔ��Cv- W�z�M��zF��)�X���α*�W��Ɉia-�ٮ�w��5������8�Oچ�$�#P�Ɠ^]B�����s��h5�`	:�i��Ħ,@�1}���Hjs�����X����a�x]��j=d�-:�]ʾ��B��|4�Uz�P`a�eiKq5u<���09��^V���7��dxE�=�/i��o�q�}\��X��cC%"�h�Ѭ��Ғ����:��<m��q~È���]$Ѕ��S%v�=�|t�6�[�V�իR�8�o�ԭ_~*��O� B� �q.����Էw��v�nd�"�̪�쥩�Һi!�Rg��ަM��c�N����k���A����Vo��	�.,�WR?ǉ��Asy��Жl�g������և�E5�_o`��Jq��z=��7G&�+5�������|�*{i �C�S6NƆ�u�tH�t^�f�Ao%sIX[�����a�1R�ez��(�����C4�ҝ��Nܭ���z��(J���>���*�?��7/D����]3bP�Eʻ�7�n1վ~��E�����
���Rl��>C��w�S� ��;�eKR6���3��ʩ���Ι,P}�z6�n�7eS�o,��m�C��~FЫ��fX�-��E���#r�$��u�粦?䢤�nP�4�R#�:��4`�., ��
�C�q�:�I""4J�����v\/B��O����.�@��,�&hL/\M�l��[Pg~��]�����Q/���ë������"�  [n>הd ���/{>#vyl��-)S���-G�o���{0:~�c�����V�9���
���T^���_���13,�4��$d�����(�1�[r=��J�W��x��p����,6�������2`:}�N�\�L���Zʆ�q�q?矧d�RI<?���sk��/������O�C�T�X=(��Ű��3-�ǣ(g�8��O0�Z�-�\ C���_�=��)��"+{-j�H�va(�M��_n��=$T���J[�U��@�x�6�3Iq��s�Ƌ��̈́��'�r�7F��$k�J����^��,�Q��C)�|��7:��E��Z=F�C��k��7�\e~2Z�+�-��0L��e�.c�?�U�~ܒSLG���P�|݅2��2�'ר=T��ms��q(�J1Y�
��c�D�S�Q�7�@���gVr���T��ː�t%��������H�Y��nm��E2�z4I�:PY9�į7ڵ!Qv�E>����_8�7)���p
	`�ف��%)�=��qz���^�gķ[��_��B}��|N�8ۉ�un����F�8ʽl�0�KJ��AU��<��PT�'/�+��ڧ[HCf����L<���G.�1���
�J<LO�m-�lđ,.l�w�J�|;$��~�h������]N�7�y2����eݯ��v�<!M��i<�kL
�}I�no=�I�2{a���;L���S/!�h�r����M��z<���qg�a�>(�M��){�n΍WӍ:g(�z%wC2�F�Q�jf(-ӈ��Rp�@\y�{ף����Y���]��%8��߷��N6u�	��((�L�ǌ ���Labe(��y��波�% �^�@�"l ��D<\,�|��O,���Ƽ�2�κ��΃�|^>�0��Q�E�ȸ?	r@�`���������z �RV��ds��$�{<�z�0y#����k(@�A_'N�gŹ�Tѝ�� ��f��MԺf�RVTw=�J,B�A��8�$�i�	;��O�9��0d|&���rg�5�d�cez�Ą�;��ג	�OD�S@"�ZZ�s[{:�h��p�G��P�e�,�Ա,#s�K��fP���jhKΟS$.�X�EX$.K����
@�`v����C�:���OG)�U[�'1�H9C2��ͱ�4kT�86�ҽԆ(
�s���3�;�d����4r���+��]�~��)=��T��z��Xx7;�#~/��F�7�{큭���K���\s����y�������� �rhQ/�Ӻ��AZU|�I��Yܳ�d�?��u7iٜʢ�'5���ܠ8pBT�jϿ�l�%�Z��gz_$6����[���hW��L+aM�K�P^F�Y�}Г��)�W�����$'1��к�����+H�G�´����m�i�t��,Y�����Atn�\�i	$4Gw4����a�t�wx� �^���`A>�ק���g�Aw�l���|S<�~�3h�'U Û��8vF������{���p艙��*��E�:�n��w�~kP��:�Ȇ���S�v9w�6`�n�)N�� ^$c�X�����gy���9lÐ;���z猏��e<�?p�T=q,��'HEtL��o��ھs§���1�K �-��)�@'�EC]�H��[V҉6�7��z%�2G>���� 3Z�e�c,�b�d �reG�#�3z�+�8��'���Ņ���9��X�U�e;���K<�eҳM���z����nA|�,T�{	�V�]�Y�X@�&!n:dy�l�s���F�?!t-�����Wr����C���z��g�N�բ�SQ���Լ�?��-�\#��`U�rx�3G��e�d��'t�����|�����C�l�R&22f9V���MDp�(]ي*j�+L��'�����]]e/l�o����'����\�?�c��،1|��T[[���A�ɹz�8蚲[�@ԟ[��BA�#�Y���n/�AG�^���u����/.80�Ow�cL�N��D6wzk�,�׊
'��}-|t�Y��[����s�^5(�}���w\�p�%�L�?`��\i�%i�@}�GK��> k��1HW,f�dӱ>����js��i��`1�d���ƐNzJJ�Bv��A4F(&OS�'}ُ!�{���ê^�}`�����v�ƀϙd!c�#$�h�ч����
]�'�[�4�^~�X�*i��E��n7Y����zq��1*Cx��^�Þ߈���4s[c75FvL�Uċ���������ƾ[E�ǹ���1�(b������D�7�>`�]Jv���Et?��݈;�Ɣ�c��^v���iC.����Cd���<�LʂZ�K��'g^TdO���1��~��j�<� O��_G��zd%k�;d���9��y/ɘ>�T�.>s{-����z0�D�i�P�C*�Hb~k�Ix�%����.u����C@pd��=�O�.m*�U{~z.G�
�jΐ�C9P ��ebt��~��d'��M/)����< <ET����Y��0��s�$2�(K�9�?�Ci®�g��!�2�nżx�Q�����[㵃�
q΁�N���EgA|�,�2����R���5Bt����G���ǼV<ͅQ�9ay'����K_R����p���rY�O��|`FLp�V���-�&�k|�;�.��yX9k��p����G=q�w$��a��yɷ���������רg��an�g�f_{����T���_�(*b	#ψX�dt{|������mELiE$�+��y��c���osT�oJ�B(� b���2eA�ْBo�^<뚧4�t���P[}Q�B74�I�����l��I�F�У��$0(T
ÃAΠ��4�K��6�M�_��ɕ��}*����/tj����!t��{����x�gB��l�b�R;�0�au%�����r�k&_.gɚk�n��x�:<��$|�i��y��CYd�,^�1��>"�7u�8�.�ϓ��gl��0��2����F#f^D\��~��VO�)�8�-�Q�^��Ժ	�<�頹'�����;�汱E�ą|�Y۝XP��n)(�8`&�[S᯼��p��%&k��U> Q�L����$�ayq���5�qx����'��`4�y�K_�}�>�2��'sQ�UO��I�k�Z<ek���p��|9�S	�^@	�E�8�7���Q��E�
_j��e�G��;D�=d1~��n*_,�>k\;�����PƬW�_��Y=�x��n�bv:��;O�}0�&�����(�F�bF��~����S2p���?=�lu����sϐT`��t��y��gl���:N�
�T�`1���h�P�g��M�yz�����t��T�c�A���,Wc�<I�L��}�i����tA�V0*^���Iю�g�u�9k� ��!Z/v��Ft��>�ʱ���Ӄ�j�6��|�ʯW%P�����'��mE�w�%115i��=E03�F�������4��nP�^��% -Y���9���4�J2:�ڙ.1=R�� OC��*ŅBܨܷȚη�M�w���9��(����_C5�(���:��	�m1����
czt��D��[����>uT�?Ca��{O��D�+x��i22�q;D*�K��p�ik���vs2�Kj�V��4%����+�Be�\�6�Q�-��eȤ9'���������]��^��"���a��٘H��~�B�S�2�&�e1anڔ��%f���ȇ�z��#�g`*	��pp������g;[%Q@P�����bc�}��F���mi�*�^�4��N�-�s�FI@M1[�zq�W<`��M7$:Rl�������O�C��?ʃl�/\�˽��F���n6@�T�����Z��ir�&�v.Qn�3� ��Z���3`���
<k̐��˗q��(��� ��͇c u^)�y|��S�oC�YVE��<���^�E�+��@+�1��G�x���J_�ZȰ~!-W�=f��(�?����2fGғ�<Y��uΈ}�P\,QC���kWm���|�ҧX`W�,�U
��{1=T]�]��Vl���ˇ�o-
�W���οc�K��R+c��M�>���*�����@ʨ��_�K�Z�X ���[�7|�o���n����n%���y��S��B���ф�O��E�Z�a��4�#��
�i�HR��
���[�)7��9�ܮ�*&�Z`��1fH��0�`A�_���h6	?�M����M���s�>���M��'�_�N� *� h	a �������i��ȡ�w�u��g),-�g�F�h(��}N�Qv��ٰ:F�W^�?#�s�I�aEN'I�<ME��_��� ����a]��#��@���#xc 熾ړ�T��K����T�Z����F����`:���qy�5�8��iN0{HfC�jIz�tH�6F,u�ӡ~)�{ѐ�ض;�)�0�Wh�h��̽���Ӝ�'i�@��3���4�e��
ϛ��D_;�Na�N	�2��	k��&���XW�P�DSIxo��a�ͨ�(�L��yK}����l�U�g�n�����e}��k��	׺��Ctq H�������j����C��J��h^N���9Z���0����8l��h[��UP�-� J�e���7�L�ܷ�2c�y��ӏ�(�-g����R�������7$�Jq�``���,�����r�N��׻ -�+X�9����5�'���j�,8�S��SSr�U�-�ڇzwp�L�R��jI�!��aڪ��J�Ԙ	�h��~ѣ0R����r� ��Y�����K�,�/ޠ���ܐ��Ur��v�R��2���Մ�oVu��>��`���߅+u�#�̛	�c�K�l{�'�g
�	���?�*62G�j�Ag���#�/��D�"�qZX˓R�&�s��3&&�ZD����� yh�a�Qϡ#4Ԓ��7�f4����y�y���d�?>ޚX�Z����m��2�8��D�!G&*������	�%��Ʈ�"�����&��>X�ٿ�,"d�ђٸ�9�=B �%ϩ!LA)Ib�Wa��]O��J��^�|#8�E���Ѷ)S�K�v荿X�[K ���Ux��W�4;h�ΟZL�~tM5vH���@�vo3��nQ4j�`ӕ�/SH��Y�eW����x䢫ץ���b�n��խ}�c�����1�Ջ���C�N}I�s��+B�ߵl�Tc�� 6�O� <hw�9�A�^!�~��s}�������<w��F���'��*E�Hʮ��gNK4�a�!K��x��x��>ֽ�T�a��R��u�ET0�����ڠwv��E-(�ǰL��x����\��T�����z�N�2֛M�3�Va��g������9�]!6h�,e���
���n�_�H�<661m��t�l�E����b�6�c3�yoЖ�<����9"���	��Ņ�Pw+��3y(2X3�]���y��Aۡr%�B�z)7�fF�e֮�0�=�:�.�#4�yL�Z7V�G����Ҍ��عݒ��B�<�-����L?���mj����[Mr�X�y~N�w_�F���F��丘�+�HP�9t���9}R�#B�K�=�7F���Z.	f�W����K%^�����4�u�x
yI����J&Ws���+9�aH�J�tbİ+��v@�REDS��"���z�s�\啣b~w�G�3qu"� "�OZi�[L�t=���Ľ��M��Ha��mT#m���HY���	8���bI�ӯAZ&��;>��a��@?�F�ׁ���g5s���V��u�+��>�g9��=��[���[���[��!�\.W��CE�01��a����[`{j��L�h^(��b��04}�T��=Nt���k� u�T1�n������G
c�r�C?����4�,�U4�u�٧(�Jr���S�lO�~;bm�y9���g(<�F[�̼h>4��( ��1��O��O�2vi`�_8钗�n�n��D��F��̓qPu��(�B<|B��ȫ��"2p�]��e2��M�mKJ�C,���G���B�_�+��
��nЭ�똨�k���L^�n���sa��<Z|�UH���?�*(yu��ﵬ�lQ?f�WW�Yޡ,��x:Kf��e;m/���l��etV��g���h�@�^q'
:���4�W�l�	�Z`�t�GH���̈njq��l�iT��w6�G�H����8�VT��}��]���!_�:�#uF)A���.[��T�u���_*�ͮ). Tm�t\����a���1T&tϞ5�]�Z)�����!XX�1Ə7�}�Ffq�jx��PD��@�y�f��T�=��t�v���	KZ:n%�h]�6�+�J�@�Z':�d��E�����]p�ɋ�����)ԭ�ө _�٫7ޝ�����7��0mI�8X��?��ʛ\�7X߲��'�b�{I����L���7�G�ո�c��ߏv��77�-*����
���k��B-C��9��<�����I	J�5�an&���t]R�jT%���\�`���K_��rw[
��#;��q8C�G�!4gD�um��e!;1���{������m{@����X���Q4,oºRP?~��m6����ّ����v�f�����B��cs���'ظY#�G.d�7��P�5�0�.��&��M�L��������'�`��Jn��P�)L�������xM]���z}��_A2/�B�<�[2|�O��SO12�>:Bi�q���o��Nt�B�fN��,k>��=���3���}�f��T�u!���^I�F,2|�=�*�pĜ��iaI�$��6��g���K�ұ�Qh��?�(��l�����G\��t���1j�! ���C.ބr$Lj<��0��R=ou���~N���O�T��j����)�M�f����vA�tZuLx�� Y�H�} 8�����м��qr����
#���ق�/W�~�_d�����
��e��*¸!��Y�od����v��r[.�B-�jt��\ �<�RJJH�Y��p�X6ZT���ګ(�����c�C��ۼ�Q|�p!!T��iR������P�2[Xm6Z��_��/�3�"���r�u�4���86����a��D�{&��*��M4��J��eS� �?�if=XC4Hh(VK\]nR��EFxdNA�Ϋf�K�h�T�	2�-��Ѐ����_�-yc\�:��:?!�&�)Z����b?��<R+��<���]�߲I���@m�=g��Ka5}�W3V{%�A�k��	RMJQ�)�����5�D9ӵD�b����1�?�?��̖3D�f�L�! y���Ȍ�����S����V���Nw�<����xٳ���o���90��dS'Ӆ�H��h>p�y.�=%�%~��X��L�T�����1CJ�V�R�����~��0�9� �do�>��JL|�y����La�ųz�z{l֦��Q�DM�%X=K/=,��OB�f��Է"�N��E���;��q50���(��"�FҲ�)�$!��m���N'���d1�U�4����^����8��R�<	8a��o���j̋�~ɳ݌nXE��%�93p�b�؋g��m�p�}<מ����~��V�ЎYVDCٿ��l�H�~X����_��3��f]�>���o���yW�ݓ8*M�&���d�Op�hz&�ݠ�Ǳ�<m@d.�哸��'d���a��ܔ/vń5��z��$�M��C"�!(z��x�s������s	�GV��N���%��g���O��G0<����c�-ۣ�`������I����G�DVܐM)�ˢ����KPI�:����nt�߁5��b��!���7)k)Ns���p��D(��ұ��`�(̻E��Q��Ҕ��z`zP�K�2�5vlY٨�}|���/���7V�S��j����CRMW~K��f�KC�w>�k9�%c�2	i��*�m�'m��"�*�zI��ek۪nTQ�b(��TJzj
��6)ک��P��7{u�5�`M2�n&�����4��#i� ;�9��ťcO��j@�c3�]5v�m	�mv�t fߋ�㞬��C��>^�<)�_m~�y78��@ռg����xaY��r��ܟ�<���4�A�	~�=��8���1����V�҂2�1��M>��դ����ze����>��fΪy����� ��f��*���o��z��ކ�?�v�=����;7ZCZ1aH�n�,��3P�u�Hpj�Y{i�q�m:}k�1��.{��:��ӏ���2�h�÷y�&�z�,#��wΖ"p��n��n��<s�8�'�-҃�v˚�p�iY���7�Lyy�y=h3P�J,��2��0��z��@���Z	��j2\���9z�:�
�F5lؠ.��Dn�\�R�j��o3qd�@I2���8����l�U��% f�6�����bh�l��n#�k2EX}�Y�H�[�z@`*�w���\�&iʤ�BZ��۲���sc0#Sg�O3�{�g��b�F�į�kb��wc-K �d C@ɧ3l'LBU�5��Q��!8K���m�+�uPx��W�F�*w��㖐���dJ'���?ǦՔ��q_���x��h��?N/'�q�\�6�v"u ����)�Q�Y��`W�is����U�NoA�8��:m����m���\G��_�!�=t��*�(��KZ�cٷՆ6r.�	;=Ȯ�2ͳZ��2Z����t�U4C�_��R����[�׍)���]��)hMá[���� �1��ul�f�����lSWd{^�3Ur�U�w�C�r��(w��p�F�=ˋn����۷���/>��I�^�X�F=?�r5w6����ye�a
���3��3���7�����`��A{��&%�)�_u����a?�Y�y���0�?��C,D}/kj�"D�������V�r��}C0����� ��c�4+�%JPf�A{ȳ������	��擱?���~�*CA��/��ڐ%
Ջ�AM��g��r, ���A�1TE��g$l��L;�,ɛY��y�I�B@P������Z=�-f���)q��@3o<����ƌLȣ�4��<���!L�k�->�	��U��[��x��̲Kl5 O���Kz�&�}�<ܴ]�2��Cj�9�X[�v��K	�_���|�Za^Ī�q<1Re75��q�z+i���D�t�����̣XI�sƔmϠqo�93���q�ʰ�o�(4�����'���~�������u�k�]�<82'�2�%�i��:�fD��~g0h�M�{��$��}^�j����H�I�x�NQ=��_>�E���%U�\`�7�0(�+��SN刱L2�)�0X��u�vŨ�djG{��%�}nW�>��O�Qa5ePr���u�����d���n��:PW;�����"!p��="޽v�+7����E~#^�a�4�Z��[˼"�Ӻ.�o�xᇽ��1����loA}^���<.pJ�{�h$�{u���u��W�=Q�v;�R�qY������E  ^pWb@gx#l�R�挵�#4mS��"C���2m]��~M6��a=w�>�*�S���]�*���v���������4�쵷�Rv�e��S�%���U���@��3C�4�t oe�y�q�83���qq
o��F.C�u���l�1��R��Dު����X6#�nf^����R��n8�� ��BK�(ȢD[��B�������j�@

��7���Ǧܞ�(SQT?����I�o��Y�k���5N@�f_'69"^��]�#@��P$�Ɩ�(�p!�+fK��������	6W8��Q)D{4��j�Ew�E�q���X��:��@�N�2���~>/D�v����zl>�M��`}"[B^�q"�(m� �L�������4��l�\�3���ym���-��NUR�:)\4Q��M���>�[�zdg��%�ɍ��A�,a���ya���i�P�Ҏax9�z�/]x>~��gM�u�3ؕf3s����)y@[��yf�FH�w�."�=ސ�?���vu�4P��r,%����Twv�����4X�����_���i����i�Ϩ=86=^�B�-ai�5���d��}���W����V���� �U�%�D����\�ꚇ�����;�9��M�7��cd�{5���f�ЦC�\o��v���zƿP4c���6Fʨu��m�Aj�����%g9\���]��5����Y�\�q0�d�E>� 9>8Xk�~�����ec�i����܂b����
��N��E�#Ƥ{�r�"e�I�ﳵ ��˺c��cdx��<:b��$����&IU��b_H��%\f�D��[����p�A�+w0������?�Q��T�Ǡ�}�;�6��I�=�	gQ/���M�?=��P��\�&yR�>�9ǥ��\2�v,�04L�#['��܋��ۓd�h�(�vȆ��$��ޱy�Ȱ��Ϡ�[�O���ϐ���]F��޻[t��To�y��|xx��޸cz���Z�PS�KJڑ�1��b?��e�c�Zo[ �8B��=�G�S�����]�כ�]�D��bC��Y>���[�TAoCБ�O5gJ�|����`� ����QBnSph>1�{�)�gp��o�,@�~Z���`����3K}'4,�	Ut�_Ѭ�u��:Nߓ�n�����$6�(v�:0[�c�l��(�^�wq��>a�%�������~�8�t���/vFufN�gLhaS�=N8��^((� +��R�	����ʯ���I����-��O�7�
�=ȟ�Z��^��x�R]� f
�ZǤcm�Lx�����J�b��P�ķ��wq)(��el�ڐW�.]{K�$����#Z�
���i_&Ĺ]t�O��f֋~u����)�x#�Yj�8QϦw�$��wUD`�]��N�!ʚ �8�HÐN�;�GkB�mwZy�kr�-���]��b��7K�h5��@y0y���ᶶpi����3�QH&������7Fq��h1�]�N�+ߗ¸��\�"ݔ���9��p@oJa�V��n5��Js��LD��?�VBpѬK�Uj٫�[��8L�O^|����Ӥ\i����v���l7P^��s�C�~���Z���d1�Fd�J�w�/�w�C�,�c�rƷ�y�7	J(��3�Ss��cS,�ݪ��5�=���AjC-"S�E��e�bt�%�FN���6[9���>����A�a����!:���qX]�Q�#4�>+�p���̒yq���B�I
����{h�k��!��D��l.7�7�BH�-���.�KqY���g����eY�����Ap�C��҆N����/_m�Rۓ����Fn���?@P^������<�jc$�'�^XKN���Ӫ_�t|��&���.:�偿i�������b|
�ei�+T�!ޚ�m���昕;�6	P�R;�T����`@�+�Z����0#y�Wt��b��:*����6��d��Ɵ$��m�[j�\їgGnd%y�@�-���ʥ���zI���7o�h�B���Sa�k3d��(䅩�& ?��r؋�9	6�����A����#@.t��>N�W�n�:�i�i�KćN*��2���^�^-��Ť=������:W��:\��/_�>3R��k�~E�R~�ݜ����:z�	�ԜU�L��.� u��z��-s��/����G���&f!�%^����D�	�Ơ�$n���#T���;>@�a�����ZY�����C��q!�J���ϋp�k�{b*M{��=���]�V�;� M�XTm���O�ބe݃@7���ur���lto������c�Y7ORp��20	8,>v��]z���vM��؋X7�'A��$��P��4���n�\:3i�x{=_rg��	���8��($g�)#UI�"�|X�C^�<>���\'kdy��	�
��vw��1��J�T�˟LT�J6�C����s�}�$4b�SG.l�~��f~�k�;��b���o�}C�8ʒ�eૼɼ�:?��6�T�W�1��#�<<aQY9�u9��/O�P��p����	���b�,�J�*bemhу�qLS�K�z�^��&%������Dc�w��#�*����:O�@�Oq#���!܍��xV)I�8����5e�R3d��π�"m�ejþ�v�b�j!*���!T���Ժ��ڕ�����9�Q��"�=rn�m���A�rv����d�MĲ��eb7��&BpP�4Z��tv%�J��f����{n�Nu���߼������_5�[*5V���<��>ڪ�	MS�`ь�?�J�ޮ�y���9���K��.IN��+��̹ӑӮO��k%Z&���b�U�A�޼;���ݢ%�1�����P�E-&	�����!�a�����P�p�ش���Yu>$�|�=yQh�+�#��qb���3�1�6E�
�� ��q�����,)�,>�xFB���1`���J���2��0Θ�����&�z��{���t�:$������J�?�)%�s��0N���.N=����|�t�]'#��C^���-��q �h5�2ӿ��;�c��]���x4�y3�Ƴ0�hࣅ��4����htam�14l���!Y�(���%��*��E�A����M�~�j�xh����%# ���%���/��;Y�5'5����{{��v�����Q��E��Ib�~�1���!��ڑ@�7:K�a � ��3�!�O8���@�9�2V���<M�qE1im�W+ҏX���ҸPc]x��):eI5x�r�po�>�����$@1� �v��َS'
Ö���p[ou"��gt
�h����k��k(���?�Y-�!,���H�ɾ�Ve1������5m��杲a+U��zڿy���tm���� >FH�~z������c�4�jy�#��@�Sz���^�f.Wn.�^�z����w��B���\cN��g���U�}(��������gf_��%��٘~h�6C�.m���%�Da��� �r�2���\�`(�fL�>fVћ��;��U��O�K%���W�]�'M���I5�?�R+N��1�0$�*^�ۗK9F���.!S�KWo�=]������"��̷���������+ZH�X��Y���^������H�l~-�k�H�<+k�U4��w^,��5��b�]��B���nȿ����-��x={�Hc�&r;h�
��c/0ٍ��.g���E� w�S{^�^6�	2���Ś����<e/QL@��ﮦ��TwA��fL�����uu���5J�����h���v ���m��%u��V�ƃtB���uE0��˔ŊG��.ͩ� 㮢 i�i|�S#����$����GF�߽L] �		�k����a����_�cys��6;�̈́c��~��Y�y�&�-	��HZ�O�M7T�N�� |��v`B�ɗ��7����t������#���tH7W�F��ߠY�B=�|�]<�K�p�9��k�3� ʈ9�L�Ӛ� ��w
�j��9��+v�!�CS����O�'U�x��U��R�����VR;x��BI�`��bQ��,�3y�Y����X���W��}���n��e��2d�H兎��AzP�����ڀ�!��q�$��+�Jó�pf���-��� 2d7G��kf��I�t-��xT&���;y!9�n��,B�`礎�h�7~*?�H*4�0F�߮c��ݼ1����~�+q���-&�f[�v�M�X�	"�3/�SW*��@n�5�$��Ta5��Ig=(�%{�\�bd,ё�s=&���u�
2����T���Fͧ��)���f:�͘3(!l����#����08����=S(��i����:��T��$�
o��h2�U��RC�"~3�L-��aJ�;����e^5"1���6�%��yf�d���3�횮�a%�R�
/�����l46D���|�|�q�'.@A�}
m�Kd�/��#��'M�q���
!gjx��5/��u�9�k�����������S'�z�bpP�Op���o�\`r�&,�b�[�)��Rem��ҵ7(ɶ���b�8U��نJ�E��O�$Em�A^�5�w��Qn�+�Ut�NEoY��zxIY�d�vH流�R�%��8`<*��7����9�����B��|�:�wUx)
��T��ގ�ȨdNH�2^\��Jn���4g���3��)��$䞞����}?4%JM������d�M��IVr^sc��S�2$��(�W���Ԥ���V���A�ZĚZp�}��N>�w�#�=bz:	��H�+;^<��}��>M}.����P�nM!K�f�`������ň�40G:˗��U�����i��'��	��l����R�}��ú��2 �?����a7��-���?3j���U���ekRu1��:y����k���1I)���I�3���{ę�K�JR	?�_*��g-I�o�y͍aBV�������k��A� X|c; ����l�7�u\W��!&�8���̨�Qb)��%o=������NMp%���Mi�"��0��=ƩU��G�ʳ*Қ�d��:�K�e.�u�Wk�Ư>Y����A�9�gvV��5�Kk$N�p5�\��d�\d�I�?j����	�9YFY�e�[A�F$GL�	�8^�1&�ߕ�����˴jK��l�$���H�����q����V~Z�J���r^��8��H��IU����9��B.�bqeXU�:䮝�)؍�>��c�Eя�-ݍ���Kwh4�[�Z������_�
 �5F���Q9�+����f�b)*0��n�A��4�箂����;��g~��v�Ӓ{78sQe�]�&��!��m�+�ȵJ��ʓX6��䚬T1���/�e��PIҧ�M/��䬴e��<#�m�]��睾u8�w=�YQ+e�ױ�F|�NMI��{6��m��OK併dQts~v���G����8{�~��3���$��v�궂Q�3�~>���x�8̘9c��8e CԦU2y�0�D"�l����]�?�����Y���$���t}��$*N��}��"��Q��C�$�F���H��H��k[��U�9V��p����~�4�qj�W���o�e���'7
��F(z��U�o�|ݣI|�
B}����C��U*EQZ��nQ���a.'4��l7�b��'�!-7�8�YP�AM`tsm���t�<���i���K�ks03��;n���0`�ݓ�>Xk��S7��J����
�CѼMkS~�Ϯ�8s�S�|�h�ޜKt���/���t��38��0��C��>�#�c�I���S�O��0�;��a6�O>�������>Z��C� 8�'��:�}p�A�R5�<L)�k5UmmoǍ��0M%���E�s�Z�E����Uؐug���[���>�+X���� Y�H6�����%���č*��c��s�:��xa'j�� �Y��n�Z������\�
sy9s���B��-]ǡ:�������db��f�,�(4���>4`�R��>d)��ai�3���g;�ީ6���!A��ǡYaU%Y���0! �8Z9:^S�$��Aն�5�By��"��ۅ�I&�ue�4u�������c���1�F߁�N�
��9uX�%��Ǹj.����#�}����Dl1�d3�hX�;|��	�(+(��7<νI�7���W��L��1=�|e�1t��!�?^+G����Q%����jM\�Չ��0>��nyIx���	)�.O�jjL;��s�d2���.{��_�Lh:�PY���&(9b:���N��G2��dj��$y��G�<�֐���ܱ��	�}��xؠ�L��Tx ���++�A`��C�ѭ���v�oi �44_��	
M]Wʍd�Į���N;��-N��'󠄒��L��ˀ]E&x�0�MSǻ������f�`� y]�@�{[f[�$��-
�~D(�H�E��)�uJ꣦3���C�ti�#1"�g�i$�^H��=Ϣ���9A���A��*>N�T�fy<�K���FP}'r\Ήo?ߛ������,��ܦ�ӌ��:.�\�`z[��&�%y>��&����d��(j!�3�{�5/��T�?m�$��1�z6F*2?�Ѣ[�ͰI]��&$8�a���ꅎ�k�;`��A�lg��&h�D���E]���P+�x4$��{$��k�#�<uҖv�޺{T�\7�.�1 �&,&m�2;�9n�!�z�T�[��-�B�F��/���UhN��2�����ݭL�ڿ�h���5ۊY�� ��f�}g6�. X��S䧂x��bP2��Xjx�L~��ɉ��I-�
X��mY�M~kv�!֫B1�\��N���d| ~�i=tH4�-̠�� ������/b/m$�a �B����Lر_zC<�S5��0��{j����N}��=�ce"|؜��F�'���s%l|��3���ܓ$#��>��њΦ���w:�ޤ������Qa���tR���V��`0�%࡭�6
<��Gs$�%kѥ�+`S��A�`��څz������MO���@�R����|�CL���'pu5 ��Ȭĥ�N@�0l�2}_��n��X-�q�X5��|h�G���}���)-�8�z)�_s���E�5c����?Z�)`���Cr@4�f��bz���wj�6���I�n�<*ʸ��"�_Uf}���P�,�=URL8L�yWܢ/}2^TH�����a�U�����ʹYa��m�f�D
�2����_2H��?KW� K����_s�co��o[|�d;X�3�(��Wle$�~W�+��ADiw��ya��$������Ʀm��>�]��=71n|�K��PJr����]ƥ�	<�J�G�Q��8l]��9e1y�y&i�<���\�P(�����r:ڧ7�e6��tPV���H�!�"FI�����'�s�>j	��A�R���P*�a^3��;�p�^������4�X�B��.�"tiSP�<y�CU��W��J���AA=[_��|U��~b4j��Q���*����A�]���N�[��~X:H�����{}���9�4;�ז^v+��ÇN�7�9�o�UY�cx#5k�Q3EC�	�?�J����}D���l�&����h��#��b%:�̜�K��/|������
pa�9��m�2ͼ���|����{�ݓRÕ��4 �����PGe�*F����!�Ey\S�96����.�D]�OIV9��O���s���e���nZ���}��qS(���o�L�{��{v��]ؑ���(�Og��p��j�p�����)�((K?� ���)O�?�T؝A�V���z��H�����Rʈ���8F1��8'�N��k�ʬ�*���I@�J��8N�^`Β9��\��^��k��MyR�Z?����HVc8�W�K�}Љ��ƃ��b|���]t��K�i	C����Ww��e�6�TW������Xo�,����_U�ڋ���On`$ÿߦ��?�� ��sAB�p�)���D0\T�N;���Pًb�T��3Ag���	s'��"u��&V6.J���.e7�O�ǻ̧'H���P�|k�m������[|���͌U�B>8�Q�hi�HM��tt����s2y;��&�������Fn?r#�W��o3̓�}�:�;��]�Pu�	ʂ	��>'�͔!�G1l]s	�]Lѿ{��و���;��־�1�'2R�wG��p@��w��G������Ȱ��~K�b���
����CK�[�F@ھ�l�k�n��Hk���zB�5C�_�4�5�>�Li�E�W�t1�=K���nSqH���S������mm��T^'��>��q�7���~�$������BGpY�J��Fp��2��+;�[K�*]e%�Ӕ����@Zfs�Jns[ӍB�+	��^��/�7��'B#��w��*O
!�X=ҙ�<tA}6�9CslC���>8��Q"	���b�<��[t~���&�M�A<nÌsy�*A��ɫ3,>��f�< �g�}FXȪs�t!�$G4���o��o�"K�W�����tVǌX�걑�X*� ���v��<E~����>�gv�<qv�_��O��S���q����6��$�P1�#�j�;�t��|�;>Rӹi���W�����#TRSݝ�v}�6�!�V`P&;�s����9@��DB�"�����(�/��&H�|�홐9�#7�i{�B�ϝ쫤-u���j]�+쉛�����=G[s20c>��=R'P:A�&��b',*-�<�w�E"�ܟ��T��~����w&��bQ�I�
Z8��N�;�<8���o��G8��XJ�Y�`z�� n�K���QyN���}N����E���CV꾊����_�����K�A�"�IoU��/��}Eѻ:Ѿ��t</ۭ�i ��*����>����ø-�r�~h�֨F��κ�^6LK�n��e��c9���I�b�I�y�Bo���eQ�����;o3�v����M�� Zﳃـr�`��[Jj3���1=qlgzz{��]�(�9q�c�64G��4�<!�m|+ X���Nr���2�D�}����G��[��
���ߠ9�Ѧ��F<I1GrJf�Q�E�%wʬp/���� �'��j��Y	Qm��%�/�meQ�զw&��RM���L��+���$y�\�X�H���q19q�s�m��L�z7���� �ZYBv��i	���W���s�w
��q�<?�-b�U���D�
�L�:�z�� ��B�rr���!����q� �_��~'Yj��K�G�l���n�?�~���!4s,)8� C���M[��9IR�h����\����G�ݸ�X�u��&^�e�څ�x�=���I�V��^�o�w��Z������,���8o�^|,�A;�|�c���o��ɪv<o��<�̣1��f�L��Im���̡�
#Oʌu>Ӝ�!Zr�p ����`�Q���R���t6�d}9��J��������(��\�zU�S�$��0�w�	f-�� sw�%ɜ#e��D���cGV�>�7ug<�/�xKx\9�=+���ɶ�Ƭ�ݫ��uTta�D��	z�~���2/�N@�:y`��[ ���O���0�xS;�ݚ>����4��+�ԪM��h�X�Y=������c������|�k��lz�c���bUX��;�BŲ6[|79f;)P�Ҏf��Cׅ�)����j?��1�m ���D��-�8?�����}�� ��?��=����bT�Х������������7�°��z�EWi����u0�F���k�VX�����Ʒ�z%^cJ{��_�ϸ0�	��X�db����k��s�S���@�WƢ�L�W������\���!��ᓢ�C�$ǯ��	K�O[�<�UB�W��D�4Ba���"芐%?;q���5�[KmӊQ������Xf���/�U �.����2fӯ�RR��Ea��а��'�^�P1�����q6��������We�DC�㉹D�/?�K��Ii�`��7KQ��|�s�vv�ċ��_V�Z(WV�90h+�񅤀�o���q�y'�~^��O��ژ�ƌ�]l|����v��(7�S��9m�G%�aǘV��?f�;���b�4{�p9�bN|j��վD$�\�%O�NdM���2fJ@�N�'p��B� ��L��Ї^A�d R���4BGfߣ*�|��3�=c�+�d��&n�n�|�)y6��<��c;�Q{+\���i��9�9C�ի�:��:��v��7��jyQ�9Y���!�����V2�x����%D��9�|�^t��M��2B~`���ռh��-�c}u���v4>�.eOa?���tNo�����u��Ml�x�B!���g�(�P��z�?Li,L���O�i��g�PT�
A�x��*��7��D�(��yez����	~�2HI��vrI����̇�?#�l8Ts�
�aa�!Q޶���NB�U��`�������d����U�oTݯHa�H�ܛ��K��Z����)`U���a�b��=R��w�\��iQOy����/\>NW\���G������	��ԋ�x{m��%���U��BD�Ң���=@J�X�5�R�D���\,9�&���&��Z�����<���Z:X�%z0�4�%�1-�%���ٓh�!��Ѣ� ƾ;= Z�lT79ͩ!�}��v�X�^�WOv�V���աg�G)-��j؃}��S��\�$�^�j��8�	�w�
�n�+C�x�A�NRA�{Hv�n2�����P~�0 -C�'�=���t�n�w�x�^���k?K\iB�<�W�
Sv[��8 ���A����i��n)g3D���6gBL�P��%Mĕ\�W��`��|�{�[�ln��$��g&>
�W�1{�˪�T��H|%�H6��
���s��Q��Q9�d�� �rl�{��٨���8����9�_ڭrf����Y�P�/{�,����c��]��l;z%����YK�K�phJ�.�lc:cL����Q윹�A�k���&���۔�{[q�Qp)F!��8�2��s������{��|��v=�_��;�9��s�Q���#��腒��h�	�H�yӣ_�A�m4�O{����0Z�3F�z��	��y���
�`�ҙ��&֡ E�W�r��-&��9C35-��z|��Mզ6��(���Mj��HQ3�\((����j�鞋z�i��6�ko[��SB��|�%qh���ì��@�t�
�5=��C�����,���QZ�3n��7�T�9����SP���h~%�����޹o��1PB�G]�U�?Y�~k��g�}Y�*̼�+�Px=H^������*�Q��`��Cw 	7g����(m��@y.m�ns��Zԟ��pcQ��ݳ.-<������ �?UW����*���z���D����T�(�T	��1��N��b)y��1Ee@%��=�h`�	���P��.�3�#�Б+�tY邿�R�[ǁ�I��ǂ�mZ�Ν[g1�-�����k�3I|��i}��\m{�a��7iHe���CT���oP4@����7Bѓԋh|�DK����gl�u���	��������ޗ�V}UЅ�Z6,8:�Jo� �e]���d���z;Р���}Ć),��)ql=����e�'s~C�;'�7�VU}$����ЂѦ�ZW�����R���i���v���:��v�XV��'ya�=`���ǜ�ڵ�s���ắា��n�H��Ôs���Y�/�m{!����V�����S�wPOE��Ek���,��d-�xY��PT���B���!�@H�� H��Z e�z��p�'~���!�ʛZ�VP0��ްA/�q0r�����7߷L+��c�Kw�ֻ�:�O��p�B�������5\R��M���m��f�
�&��d�D
��S����F��'����bX������|Ł�cU��q�"�K�0���|�[孄{�����/H��¸O�pXi�dх�
z�Ժ|6eg��-䝑��4�kŚC�kpg
��hH~����ZQϭ�(O�n-5�Q+�P�Y�>c�q��e�s��j9����g���9��X��+L#�H� hKL)����^�¤E�B���m}4�mpƾ��3�2�z��t����r���n�`s�,�BX5��a�CY!�Q�G����(31�Y�k[Vo�#��U�iRq��P̧(/�>1�)�����R[�2��Dt����6Z 7��N�����L�.@:�&�˷ε�>����"a��Rv~�B���)�G��e��uqs=��$�k!�e��:���W<� ZW�����s;-}z�T�7��LF46�Fr�B�y�m��-��{�~�_>�MR�rZ���H��Ʈ,��9�x���wg���Z-`�W��?� ��]|���;1R�q8JGZB
�!��H �����a�fx��!ܱeӀ1V��a�	,f��,m�/�����.��x"[e����@�����v�)�7�Z�	bU���1R�#�D���7������q�#y��v��&6ʜ@1���#-��]�@5�w<ڡ�eE��vE��3tK���jt�Y�t� x��>��)�O��\���hI���U`�\��P�t�Ø��L�u�_�:
�]��I�3y�����2kVk�޾�P6� �_]���a��9�%��T�0��������C�a�N��Z�Đ���k�Xm�te�4[�LC�_>[��3��ݦ/cf�S.�"�Fm`�����X�?N44�����Ý�y�N������!X+��K�03I����j�>�V���I$��M����Ni��S��M�D���_�3�n��Ϝ��.�ώ�b���Rb6"��ND��զ���s&�T�&��v�{���6*3�5p�@S��P��p�62L�7���)�f�a��A�,�}�4V��DeR�fx�b�T:/�����ҥ��RVi��*��a̶����'(�����"����BJl�y��,	��y�;����}�Ϣ~x�|�c0��w^��-Ub� �>y�8�����^&��O��B��b>�x�ѐ�a@��Hyd�m����u���,j�G-?�}�R/�}�K����kz�BB��C�ޚ�J6��QϿ�VD��n��V�/ة��E �s�ܻ@� fu�eH�6B���g�V�����=�s89�]-������4, S�s	��T�����4��?H��=N����%@HD�c������A8���PAv�X��hZ�չ���L�Jn���~�R~W8�6����:���g��PszFN���Y� %�(;T�6�����7:SO�������q$�|%��(�m�kɾ?O�݇x������n��i��Q}A�$ߩQ�_�_�`9�o�@1#�Y u)č��;3������u���cf"�>v��r���Ψr�rr�ۃ:M�����SZyǇj}x,�,c��A�����4#|�-��z�J��L>В�l���6;_�ۧ��ѡ��*A��G�8�QN��S[��_�`v�\%�̔�I�U�����Y�T)X(��$r��<P�{L�'>_3���d�_i��r.�Rv�/q��ť�d?jK�ˈ@��r�^��Ns%j�FAo�и�R��{�����H��M�4��h�����d
C�3�z�--n"e�:�?V	uɖ`��w�uS�//��2�Ȼ�D��Ү
����]!��<!�N��~r*t &%�k*��;v�'�l���ޔ!�8�!�<
�g��M��TYP�L�p0��*и	�U��n.�K���"^y�����^�l��j�p� ��G`|�v��:[]*q݌{<�ec� G��y��J��{JMN:���9<Ìϖ��h2Er2�+�șRڄ~�䳤U	���~�i�F�m�Z�T�W����M���;�&�Ŋ��lwq踍ۍO+{NB#zx���U��Dz��-�1Q�ޙռ�eA�)]Ph���.ʑ�F�T��W��Rg
��iЯ����kKj��I�_60���FF	�y�px-�oJ��42qą�\G���8m�n��
'cu�1�D����mD5��;W���6[Ш����C|��*+G�z�
^3oˏ��Qwg���!�;���M ���P�f�v��v/6g�	P�щ���g��+Nb.�i8�ߗ;ݙ[[���sd]~�-�9mK�5�������b��V�P�ÿ3��9�H���B�ת,$�	��5
�s��m�cxOwK�q�g�k�M�s�jS&<"�wؙJ�5a]��ͮ�������>.�t�)��L2�J�����2-Q}y/1vr�����|qY�$�Ғ�(�1�TP�+��vc��k�r�#1���㱃���9)�88S1���$u6���<E�FWW.Н�'wۗHS��q���Ԭ��ف���O!�O['B�E�n�}�j����s��`Ġ�ċ�����=CGZ�Z� ���[ce;���n���>G9���w���P˚����<�p�����mn�*�}j��8;C6�I��\�i�U����Q� �px�U0�C�HEar�%4r빦&��G���a�/R�����(z�X�у��ۛ����!�E�,߉���J'P�!#�&G�,�F��K�h	v]��V�Vkmd���&�tILo��8�}���j����A�˫$��FX�x�+��Ǒ�u:X\�MOKt�S�)T�B�{�o�TI����of��~�.�R�Z4~TЅ��w�zO7_'�A|l�B��-� ̀�cɎ4ʶE�kK#���bRyv�M�qu��K�]���QC�=����O��k2������ �{�)������*��
J�V�).�U��dQ@�(�}3E�fմ,�ͤ����h1,�gEKPF}���6?{]��W��X�hK���;�~����P(� �.�N�P��A�}?Y�*.�R#���;j �Ԃ�>�
:
��{G��aP�}�[����)�ˈ���/,��y�G�Rѡ��~*��A�"7�HW����_Bm$Hdo�B�����d,R.v�򩇵*su�Zi�8������5��_E�ȏ1Ȳ��`���j��c&�O���;��NIM������I�Y<:�t����2-rS{�(�$d�8ա��q٣{������=�Wf8JFk��υ��L�:��+�)��_�35Aby��z�OB��k�� %���*�Z�:Ybfh�#�b���'�GK���酛��}�6 ��[{��^���2<�(��
F�%�t�	z���ѿ�Y����!y�3"<���H��j��.�� ��(>Ο���t����*eʈC���i��~��
l�noeC`���A!JR;���a$M����-H%јja����D�)�˫�=K'�*�=8�F5��stճ��Y�̮L�|X^$�Q�ʐ��;����.b����l�G����m���
�n�22��V����Aܲ�R*a
	tw���|�to����3�����]��D1rP��2ղ�S�2�wԌ���'KT� ��}{/Uj憸K�"<�p��G������ԙN����e.v���Fb���OS	���:��^
�>8�`iGhrY&N�o_C��d�ؓ�n���>W��H�
�yp��vhX>Jl6���1��]�z��(_���H�Ȝ�j`��� 5<���'/�焿�#�*e$u=��2c��J��[��j��N&�Ĕ�A��C
�Y�!��-/R*<eG3�9���`���-������0D��*
U}M?�MQC��!�fw'j��t�*�z,K0SpW�
m�k�KD�a)(c?@.��8e[?�M ��c�#�2�fQ]>�MB=�����ټ�(�[�<�n����I.d�ܟ�r�v\���(8�9c�}��'�-Ϧ��a^�&������]���>�i���M����D�%�hcsR�9��z�I�'��p��~��~��֦Zg����O�u<���I+�*�y��Z,�z�A�=9W���e6](	����I�#��jO�5{c���������$O�$=����N��� `��й\��w����y�7E*e�6�$�&��|ۿ��p;�  �xXSw�i�?�m`�P&{���]��7_�7�:[�P
��CB�;��%Q��$x�٢zP
�ν�]VύVsŢ#&-}����p��h�$�Ğ����j$lˈ�0��qa~�f}�������ӵ��g�)b޺��bfq��
���%��8i��lf�A, �_���Lpդ���ҧ\���e3:C����)s���]���~��Y����Ϙ��^ }	o|p>��/ܗb����&;�F��O	���_���5c��Kt�؜��F��B�Jp _�獣>oB3���By�}E�q��p��Q.�Ӌ�~�\Cxw+^'꾗�7E?�PtA�Iv���D��n�L4��˝!�6w3�+G����jC��9�:�V�GW��6��જ�A�|FbY�����m���@[L�oa�h0iBĤC%y-�(ԇ E����#�^M�g$e�舑^5p�ܹ����T��P�)t5MҲ�3Ty�!V��Z�Z��%^����T>��0b�G^L����hJ���?���r�|G�b��A���GA5�G[��L�߮��u��#!(MSl/��o��|��f�0��+�-�}hrp4^L+�-R4��Ͱ����d�a�N^�r��4�WTR$�	���_���J�s�P�����#&�?*�8l�$���d{�z�	:����ϓ�r �Q�06H�����mYGF�J�uզ�$WL�H~;���"����l {g/B]�J��GJ)Q�Î���>�l�rzP"�(��LTڭ>�'k��U�c*���$�s�=�˹)И�Nj#���-�
�k�C�7Ws��M�S������i���M�ݽr�<y�^(G�ǃ��k���au1:-$�܀@#���V��}���_�K�Ws�+����ת��hg��Mw9�5�}:��g�GM)OwT��P��f��/��$Xy�v�ވ.�E�&���>�ԥj�%�O{b����y�G<�/~Rx�[y���#9�p�BU7)bH�M�0� �*���Яpy�i=�����E�����VU� �J\ղ�����X�]���"�b5i�W�nL���m7�T.P��ϏK9�\�<Vw� �����4�¯��U�O�tnך�����P�53���3�1k����g[�y� a�o�|f����n����
A4 �ͧ�`�::uYl��X���:�U�4�����P+��7�#K����ԣ$�,��?@uԁ^�r���o�� ,÷8�R�)	�Ƹ0�x 2u�6'[7�`>_u���\�Rg
�5�����]X���w���'�:������*hxLs'�ޜ���#݀Y�܆�"P��֋vV��)>��̊�`9q跕����2sn!n��K�u`)Уe8�W&Z�Ƭ�hk�G�E�����uWqYӳ�y��O�׌'�a�ɕL���wzͣh��8�(F���a�8bB���\���31K;8Q�|�	�����p)c����֒�4�_5T�е2Q���_g��&RO�@8��V��`��FtH��S�j���_XYM�^Ͼ�b�Kg���=j����h�i�>��~�L��_���i2}v/�wF������Wj�(�e"�ݠ8�F���Ÿ@�r1x|�2eH�Fj��t}SgC|5 F v��޳���.��4�{��ىs��o*�Cfu_1p��@�!d\��iήV��dP=v��,��ӷ6���[�|��Ѥ�3��LƽO��E�
c�w��2�l�|�X�0��U�Q=p8F:/D�:��F�fa||Ȗx^[1n ��$��n�f���u�%єUY�ױnkr�F����Ese�9N�ui;h�Q�N�/J�eL���E��a�[�"�ub�!�T��L�
��)��ZCZt��}����H�)Y����Q&��GP��IPw�Q��}�x�6��%_�r0�3�c�����;��w�N��<��ϙf�=�TY��ݢ��h���� @ń�
��@�@j؏�w(�k !=]����&F}�8���܃��(f��Zj����f	��K
N&�\�S���I\��{ߠ�:��/�(�\,���˯&�O��Č��fK���:�UY�Bk�rt�֖��!�0��T�=4�;�i�I&���onBnTixA���x�N*E�<��_��@#��%�f�Ϭ.ɔݖg�+���(ȟʡL`(��I�Bj�	�p/�t���vrr.ƞ�tA���rG*������)5��!�,k7K~�N'�A��q��/��2{=��"l:U��z$����)���/�=y^��,�K��̐k�@XK�^�מ�f��|����"4|(��D�y9'u7V��_��a�an��i��X�X��N�8j��ɿ���Wac�ꪾ]��gx�5���h[Np;�����S8�c)�C>@r��X�^J��F+��e��҅�*0u��K^o��.��5�(q`�v��B�a�'$��.�퇣c
����B4�k9],-���i(�5ݚ�(����U��K�|��i@
��/9
�=��os�s\B2�{�<l��aHD���_^�@�찋����#���G�aY,�T?`"��%�i�U�K�A��$����%�SH0�\��d�ic�k:@�}�����~{����3�N�}�%ʌ����Quӣ��r�y��mHM֡���y�Yu�x���p�\�q�D��r2�=��T�ƾ���,3v�1dW�JQ}/�h��+��p|`ׂ0��G���2���B*�8�W��
����K�w���d<��!�p���2�zs�!/*�F!�)�G�'�Yf$a��{V��o���$�ـ����9t�j]U���σ���H��Ծ�ȸ�GU��JiL=Jh��IdU�|yp��ٷ\��b��g���-��+����m�{/j_ߥ��m]>�<�LQ:q	
ijM>v��mn�R�bx�ɑ:#�SI�LԼyx�_���3ŀ7L��d!#K_����j6f��i�;�^�২a��������Vc�����������幑�p��R<���9�����,^�V�\y.��^���x�O��1�0��v��xb����T�t!����q��;5z3�,��!�&���q�%D����#���s��8��B�%��gY)�����=�̱��{�A�/8�>B�_�C�7ΫP��hKF���Q������I�	��Ǐa'B�j�z�p�D��8[F�|���v7�vR��Ȋ|\z��k;��u��v(��6���q�1b9���у�V�0��MF�6�;@�}M���~9��P�����MK�Y?6M�,�ͬ�؎�`�-Y�_ru�q+Oj�&7a<�1b��=�Ԩ����q�\�X�����d�qiq�[S�7LU�Bl���aJy��q�#�����>�>6&�t���qW{��&u�P�>�JЖ��`튌�U��rՙ&�x�*�5�67M_�p��\���4�8����9�{:�1���E� ��7�#H�z��Y�;n��@R���/���$}w�h�){�^�P�
��I���*is������!V ���&7�Ù����C�d�k��pZ�߲�r<�h�RK�ctby1 0pX�Ֆ-X�T5,������] $��žY�Ϧk�V�%??������̔�ns	�P��41�fը�����u�I"����X�/W�a5���V!�!�߫L��Ғ��IU�lm��]&�A��Q���L��W��d�lN��=�I��K*�cAL�Q�#U�=u�d�d��*�f#����yZhY=�\";^�Md���.]hzr�E�5�#*k�y��>���RTq
b���U�(�\��q�o��`8Oq>fiZc��{e���;�^�_ؘV:��,M )<���8�'�1�H����	�'�I'��'�I9�ӿ�!ޕ�d~!��,_H����-L��F�.�3,������u��}Q���3u1�����aw��(���۳�L'������G�mT*�
8ˢ���
ke�t4��ѲdC,x]9�N��<��U���ӫ�^sݛ�*��M�9v(���9CJ��EUj�,b��d}�O%^ky���:�qi��a���+���F��#�\���"(G�����Mڀtw�������f�x�i���Þ(��r䎑��L�F���k	9&*w��C��ݣ�]���zXs��p@IՉ��>�Yy�	�o�sƑc�5��k�0�+.�4�=�Ֆ�E���-�ȊO��z��[s��F>��#�{�5�<�֕g�b �ap�dnſ�f�?�b�;���/�MS��Eud�(ƻ�K��TI�	�HsV�%�u��0��ь�A�ѐGb���Q�@�-<�X����?VՇ� w"c.V��ݫa��W\�z\�6���_���d�r�n�d0�`=�>�r�y�����}���f��}i�?��=��첚=v����2��$�1��WawK U��A���&��NW��P.�����y_�/��K�W������D�o��4��Q�r�{Z��0s��PwӷQ&����2�I��!�}���"HT��35g%d��ز�қ:��)���x����/� ÅK#���.U�'�=�����f���w~�:�������c�Z�%���s��f�o?Ho�<a�|��I�;Lu=w��-=�6�g�F\����71�Q�A��(ႆ;n����qJ�8��M����Έ󠅤�<睛2�`�� ��vA)��@e�Q�r�[����	��"��l�.��[!S��t61�P=��!u�Ҭ66j#��kX��\]���,$c@�f٬�Q�3}��7u����bLӗ}z��>�N�߉�/�$L��7�E��_=U*��C�l��$�D��?R��ڷx��6A��eQ�P]���<� �,h��'9$��p�^v��H�CHƎ�� �Nݰ)�9�T��c���U��q�zAV��H���B?� {��i)��ڄ'&����n�=�6͋XT���qg���4�x`��|7?���F#�(cM����X�-.�Т�-w]d�����#��P�I�.,�R���d�[5?�%��q�V?X��4Cz���'�.$g����\�h��:�2�UY�&�A|��4.#� �Sr��0���Bd0�;;ꗢ�ѫ|È~�h;�P��.G*<�6�6駬��ݷV�[�zZWmKvvV:9�B-pR��s
�� ?�v��Wn� G�i�g�O�Ϛ���=��N�|&/��1P��t�]�T���9P�',,`��3%$(͟�J`ꮻ�$'�Rp�>���1��6U�I�]ф^��԰�oIׅV���L�cD����?Ƕ�3a2��ã�\/��u}ۂ	������>u���br�v��0I�&Z�	W!�@bF���I�%>���E< ���y���A�ZC^v۹�CǕb(mѮ>�qg��3A�`1�=���0s�r��ƺ�?,��t���);�_H�|�eoY���W7���.PGJ�Zj!�b�*<�	Bk��P��ƣ~*P��v�ӱ���u�Ɨ�*1-�?;��G��wc�t%�8��H�p�l �x3 "���{�j��&��t��+{w�*�j䩢�9Ō�)~[k�~���?�`�	�I�hx9e��7=�l����	!�I����������NW���ڏWHO��Je�-f�<��E�` �83�=$���ۢ{qu�i���t�.��_�Ew���t�d*��c��QI����_�;|i�_F��\)$כ'B�9b�ۉ->u�A�}�3.�ѓɥ�OcXM=e8��K>"Y��g.����ȱ[pwz8����JE��w��1�!y��LJ�Q(X�6TZo���P��L�Ko���,��LD��$
~�E���L�|���ѯ�yKl��!������1� ����<��I3J5��#�l(�.*|]��2V�q (��SuAI�D�k�m��+�)6�0��7N�5��䩨Em��&��f^ԴLG4w���_��g��|9�չ��ls�#���?Eׂͱ'îRh����6*o7�[I۲d�jgU0Fz��D�pڂX��'�Vd�B�8��"�4� �����-���.l�da���&�@*����=���Y�rC��M�L'(�����%�����ǯ�cq�p�H]��Oa�n!J�J��3S-������o��YG ���UX�d��*��s���@�<�g��:f�f�<%��`O������`�$1�B�N[��=<͜cǱ_��k�%�OY6��#z�e�H�p{�j�����J�w�?z�
���Ax�;M%2iɔ���}��v��d9^��%:�_ջV��k��O�:m`-�N��z S:��{���KF!%��)I�6���L�!s}���^�(�b�T[,ae����=fzn��+`�:*d�⣩�I�t8.=���������<����mIi(<�i*��쯥h,%��F�@��6d��#<�vA[]�x[����&���0'3M���-U���c�řF�H���lq���� THc>�^���,20_��[�m*��D���������/����t�Tn��8h��Bca�:��T��[�Gg~@#	�PQ{�����������j�v6�,����rIX?��N8����Ĭ�|-�ý�a�6F��t�	��8e�ǅ{�re|�A��2V�b�̂}��BE,�x�˖�f/���Y*n�tb�"�'nT�[�ŀ-m����lK7������z��Ҝ	��J��,�����B��QUM76A�����)���o�� �9c4�u��:��ݧ� ��VQ�f�k��'|���Ãj6��36؟-?2^+WT�GF����Wtr#>ڐ���!Fd�[ؘ�"^�|�%�*c�Wv_�,#��rh�\۬#��윯�>5PXj!�{������ֈ�>#'󬙙� u$R�$?�a�]"d����x�s��I���}ks����5z�b޳�g��L�2z8���=���
�Ge�n�ތf=*�kOʭ�hn�Qh��c>�ޤY�x:*Iv��g������ގ��&��;�����~_?��y1t�q�6] o{粶d恦^�+YZ_J�H6-BBT%���h7̢�QNhS�c���N�����_G�beڣ$M R��Bں�I"uح1]��LɥP��JS�0�⣞�8�:�U�5e5E>5Z�v�kI��a�WV/���<�R�޾��n}io���w��<a���%g��u�˕�#����X��b����� ����"�_�"�~���ٶ_�G#imlW�A�_w^]�K�;V �S}�}>̎~EQO[ݛB~�-\�����c�u{DB@T��w ��//^�J����j��eB�DU���ү��O�3N�mv���(/-e ��K���c�w!������0.�oj8Na��Ef��������J��$2������e�J+1d��S��oW�
�<�F���rE�F��"���K��iXR���r`@�+��Y?/#��u�=BЙ�a.`�U}�q���#�S�[b}@�?%��^/�W�C�O�����d|��W�P���T,�Ԫ}[s�t���b�*�ʚI�<��d��&g�x���J:�\0v3q(�yO3��S ��J1M:�fL��е�#߇5�^Pթ*��A���0�˯����3\Q����;"'+e��+���͡8���G����
�6�3����8�����Hz������x�r*����1�&�'5p�����qx=����`��b�@3ҿ-ˈ���
��M����W�r����+!�)8n����G��D&[��{!U���<�ES�<��}��s�{{��c	7���$�u�1�G�=|TWbr"�s��å����T�=Q�OvX����N�t�%쁍�,5�ǂŶME��>)22#�p�ݒ�]���Kk��|��ɋ��{�r£���o�`�QE���~��V\Ɍv��Wdx��V�4�\=:�T����#��Ш���4@+&Y�#t"�7�?@���C�u2�j�ۨڏ c��EPx�A��]�#�9�/��6�.GTmC킧�a��~�e�Dh�e���(MQ��w�u�(]3��1��j�4`˫���+E�QO�|�h���5�>�.n��n��M�S��9��t��^�~J��+Ȟ�$��E���LB��#"q� ���kS�
��)VPJ����fs
��=��kW�L�8���h�n̪*�#ҵ��!|o	"�=��ߕ�)��s=GӉ)�33�={��S�?�^���$JWG��a��n���Y+��ԝ�9�FD����CY�+`��f�;2{_Ri?�VG=ag�ו
^��T�{j�K�D��鴹L�+�n��3�XT48��*���6y2^j'�4���"Ǡ��G\|t�7����K��@R�4�K<�U��Ce��4~��xfJr׏�+�m��\G��f1��aH���;a�AD��o�*~��(:�Gl�x��SJ�q��O�<OW�D������48�y46��?!�YN"�{�R
�\q�q���%8V�@Z{$���\=T�3��r �v���`{/U�����#���v#���o�풓�H3��$�BH8f��� v�.��� ��u}	���0�9����~������@]Ԓ#:��%H�x�D7���!�x��5���O��F�ܥh?�vJsY�>�P�,h� +�?	��N�i1]ҷk)�o��<~���m��Mƺ�O��ffz%+�o�Q���~���3A�'����YAF؇I�R��/)����d���%�!xzWCDɽNiy�"��'��}6� (wt��������׎N�T�X��2D�����B�Eh���R��)iV?�F�fy�i⅝�R�.b/Hp�l=p������H5z��3�z �u�+z�Ť�&/<�p*|x
�q~H'�r���)���!�^DNF�6P+/6�`�v�Y�0=�
V�s�"�/?�����,#�:��'|�4��w3�,��óLfv.3�+���j_&��# �AfoH�r�v}O���sq��`/not�ڑ{��0�L��HܤXcW��l��Yo�X�_P�&I��[�{\��;mY~G�v���#�%�Z��Աe i��T|$��sNZT<�7�6����e�_����W���@���1r�g��!�����pw�~X���]M>3)&HW��t[ߞ^�Qo�[!tJ�P��+�&H�����<�����>�h8���qz4�L�93��QF�*��i�v�򕖤�t�>���En��"֦a��>���Xrh"_ub�$�>�`1�c�d5������H/���o��H�b9f����6���*�6�&?s<F��1eLi/8y��8Ǖ˻m0�;���\Z#�dI/�N}p����jd˱m�&�P�Sa
^���������Ī<+�u�X}��d�r�k��'�S����O�r�sٻ�S�z�c։'�@�H�b��N�)��O��ܱ��N:�zw�~,mSS��
'/'�d�?��Q����gҭ��$����� �c̿4q8��]%k~,��)0��Tm ��S� cќ�O�/O��� M!,P�p�E,D�):⎢l%�3��s��`]ѿ���[n&I'�)��d�7�l���C�˕�����Bץ�`�K��ک�W��'��M5sfh�bҭ�_!�6X�s_�}q�T��:�|����*��O��<�R����s�d�����xztF�Ѿ��&o�jF%*���T*;;ǲ����@���=��Q�Y͋�GU��Y��<��JR
�@�ϻ�Eݳw��j�5/�3�2�T:N$3޽�}Q"�ȱV��[�8H��ͽ�,���7|;�[�o٢8a�>i�A&/3�[�-3��h:~ePu��"P�7�"I�*n�ޯ�>�"H��(��||G	��E��xct�]!������]c7��T몊� �yw=��E#�*K�����¥�ڠ�m0��!l��U-�to��U"��
g����pgQ=?d]Y�cxz:�l�؜���[�* �NT̆��y�^�Zx�7/��I�L��2�(��p��W��6_���Y1HHNF��c�&�z��F
Ts՛�}��.�f��8�ݬ�'��A@��R��D`��@�\�>�1Y?Y������G�)�D�*#;�f�o�������T�����
��$�!l�"��?�n �r�2��Ӌ�Ẏ1rԬ�r��ȋI�y��/� ���]ALz��/�~��(,�5�Lp!h���¿.R)b�RT�G����rMY?�D}�����Ń�L$�.���-�p������A�i�L������AT�h��<�>��Ӽa������쭾�Z^͵�3d꼫L�!U`N���� m�S�V��sٵ� e=Ro�ҏ���C-m����-.�a����`NW�R!b����H52��"'�j"���1ػ�v\�^�<�X��Jl�ܶF������ba����@imڭW�䇺{�h���_�cZYB�yh�'�)Q�I��u`ko�����W���.��T������9���\]	j�����'��Rr�ҙk��^�OJ`��o����g�\R��v5iл�K~�кS��0���ME9[<�7�Ey|�.2h�3�j�#0�]��I��${�Σypı��m�2�N�3p����-�X�'Q�/L��9��<�k՝��zOlwg���I��~g�Ʉ�n�Җěx����~�����J�{��C�}��}[�B�����7=S��p%j�Ʒ�A0�T�&�q^i}dw��%ꧏ��rL��z���p�%:}h3�E�M��'��&ݯM��V�D.�;�,]g�	/Oq���3z�(~����W��"=�4O�0�Ҋ��|�2.���ɹ�톩�:y�p�f���ԉ�� ��Ĳ��-:D����̢a>���P_�)s�����&�?nh����
N��}v]m|O$���@�R�Hob}�� �N�:��L�!w�օ���+
�xQ՛��ÂY^y���J���^�5J�'��,� �}a���&֔�d|%*�E�;+�b��?��	��vN�������=�7`
������Æȕ�	"��&e��s�y�^@)yJ��?������-1�5�S�����[-u��Җpy�n���f����g�6�j_�����6-�ʨ�9�J��ꇧ���R�w���Y�2�qp���HJ�ƪ��	Ao��l�>�I����R���/�Z{���C��g�(���9�;n��&'�K�
��
@��s�5p�Z�#�S�$<o��R�� �[|傔e�x�Q0��FT�ѠEP6q��o#��-���Sjk�� G5*��؆�X
�Y1�-��4�<O�^���Q�[��GE���\�t�x��
Η%����(��F�3q��i��Q�р���_E�l�C2���!.�4m����qTΰ{l�w��|o��>y�^%YeÏ/��F̚�B����f�w�&z�>�&F�p�ſ�I$&OA5 Ǘ�:�R��w�h��+$4�A��S�-6�j�a9ۋ�1"d�K����'^�j��8e�ʧ�ܣ<�����$�h42��]q�J��gJeZ�����U�{��~Ua/��N�d<y�h:�;&���_,���I��l���?C��l�_��gq�Z)�TԌ�r�]0^*d� 9F�yŸ�f�&<|A7�9��"�0m�)�Nj��� ���t�{.ޓ�
�6��GqN^v,�@���m���{p)z�*w�*Ѓ�)�;���4-R`�����H��$��WTa��	rDvo;���Xhq���גh1��_剠���<(�������E��E�s�Gh$d#-ݫY ����Ԃ�!�!�7a)\�|7�AH�T�p�s|��0���b�$��y��rdUrۢ �0=�� �FK ���2=��'��ul	M_�!�$rTT�hр��vs��e���lQ��Gl'8�Oƞ��o��MU3C�C�ߐ�B���X2�u<�3eЭ�tH��}���)M�d@@\b:ć�)���d*�+��`���U��.p�z�^�E�����\����,�`�J���l>��w�]�$�,���brY|͢�2%�Q|4�X5�tیh�����8�<�;{�PF�<����K�?jGO"{h��bq��8�7�I��4eW�`>~>w��#�2 {��l�)8Z^����c
y�f�%=] I�~��b�{b����S�Ԥ�v:�jW��)��j{�G�z��}���.��يٍ]�*0WY�t:#[Z6_V0
��� ��`A,�� /)�q�͟{�E`.uI��,���bJ紞�4�%��f��l�K7��7<���=���% ��!��O2�jV/.۟�0�I�
hu���R�sS���؅[�<�&��ljl4�Fs���M�i�������x�P��<�ȴ��� 0�qMYk@�+����2`^�՞G��Y#�;�󪽖��v���������a�n��h�V�˧4��3��!�~���?}ηɎ�[��_	$A�+�t�Ȱ��7�)�����74��<�c�Ŭإ|b����������^S��d�dᩭ��%X~�j��G�/��M�sP�����~�er�6�VN��lx>�%'h���<Q�*.T%��T�Wæ����d�L�'�B�nЅ;i��פ�s�q66�:��[?�k��˦�%�&�t�D��%S�d6�F�&/6z��,刅gx���&���*���*V{��e�ˆ=�̠�a)� a�E��d�Rmi��L��z�s0�������FP�A��� ��rt�Qq|�#9��XRO�/�a�������	/��0�$�4�{h�mL�
=0�]|����+:�Ӛ�����4�R'�e�q��U���|�`�>0�v�k�5o$�yv����&�>�킥m���<��%��I��Y��]�Px!��|�7��'�1��[^HY*�+�ӝ����d��)|�p�Z��"�E�p-��
�#
#�ꂣ*���O��>�>��:fً�Wi��͌仸e�-���O��p�5jY�c���ϛgo�MB�+5҃0���w���ϱ$c�3=t�l�c�QF�C���LX'�x��2q���v��v�
F�r/{|v��J�P��j�qجpٍ��SX6�t�� ff�F,�������ʑ��胸����@?ƙ�`��i�k{�9�2��)-��p_b��X�+.��X�� NS�qn�$��#�d�*�	��c���q<jW�hKb�2u�8���;��SD�B��c�j��ܘ��fl��)[��[a	�}�����c�W��a��^���g�%�F���՜�E%���:��`r���3�u�*g�4�{��:��U��"�����B
���nY7�(�*2�J��.���f�	�bn�$䢖t�y6�Oc+Ӄ��Y^7Q�<���j�ޮg5�����fR�m��(Ʀ�V]g��
���l�b��&Ri�n�%6��oc�Eד���X,x���K�qO��W�%�7S�"�6����|���s�g�{xg�6
�=��32zS�)�9�����yי�s6�$�YH��iM�G0/��>m)]�1��.�G��	�{bC�i���*��D]A}3:y� ��uY�a�#���y7*���*_�+g"ud	��sޥv�;���{�K�(՛=]�����sփٳ���ſ���M�rӢ7x
�BX�����%�d7�����@p�v���^��?j�kK�EQ3���^Ra�	�����z�_����B�ic�@�����L��;RZ#^�"K��MހQU�)mH�?�ܤX�-Y�{qVj®��v!j�.RR�`6U
�4͎�p�!��X�l�e������3P�B��"_җwrJ��:�#9��Vɀ��4�=*I@�G�ǻ�B�Eg'��~��%��S�-�j���!1�A�\U�$C�/�K�B��6Ȳ�WN:���E.)��G���whq�!%�}b ����������w�`3��>\h��PXf���ʹ{J[o5�di� u�|� Z�YӤX �"?�:?����:�rS�x ���\��~��*��۲.��@�"��G�<��;�p5��G�PY�������V�*�rOcq֑~xc/�Q�3Q9�)�R&$?>2�{�e�e��#�/~6�8=�p�-�fH-P{�s��rA�,W,��
��'U'��'zPw%۞63�c�~,$MjM���E�.mZrV�Yg��L+�u�)n�lݜFv��}��2[�B �v9ci0k���3�;���ZI�	���(L;e��
�_�H"-��Fǝ�f����=���~�P)�����h�R}�6�<)��M�x���h�Pvk�y��C��.�aM�u=�zz?�6����q�Y�����Z���}�Q�'DN??�6��b�����F٢�����R�ǵ��>�ThA������X}�F�A����Y�R�z[��"�ZQ���a!d�����/4�c.Bd��'�'�(�b�>�����Q�����_M�b��n��7r��_Wq�Ť;a�=��8p]��o�厾D���}A�#�׃;P�D.,�
�K5YS��G���%�Tt�x�ҋń%E��gF��X�]�;���On �����^�~�i�`�t����(Vd�_[I�>�2�e%I��H�������~K��4�p�n�lЫ.^�x�^�	�w�8���Z�m�A��x�jر�7ڑ�7e��!�j��b��$��w�F�� �^G����/+����EfIǢR�&Pm�aQZ��t&q��N��2����҄�49���{b5m�p˾�k�f74��2Ykq�i��-7= �;$��0҂mW��V�x�2���5�Ln�>S<��=c�������{�Yʍ�}��Y��Q�H�M8���dzj[���Κ�^�'Pd̯"�άfEܒ�D��'oȲ��=�њ6$��,}���gS��?]m<_C��4;�Y�Tx�WՔa�eHƙ`�9��f������vG�&ח�)���m����v�1���,��}��TэS��gR�������b���Ve<֦�"?��#�63�Hq�8��IV2���P��1��=d��'#�0�t;��#.�v���2
����*>O�|�A���N�yl��P���J�Ѳ�=�ݐ��|_u�nrH�_��7@�x㿗Bq|�QED]�xv؉FwGf�װHQi``���J����4R����� �|�O\"����GYͣz�>�o�N]��2���!�t��!z�(�O)P8�f�5ֹ�r�~̆�*>l{��1�U�O�B�;>��]bɗkC2/�E�Z���N�k���>
A�T'���E�����^��2t��������f,�3KZ<}4�n��%	\��y���D�4�_�0���^�=^�kbt\]EX����G]%\�8M1<m�>�{r(����`]�S��H��~���5�6t��T���J�'Az�fE:����}��0�,ڐ�?�~|�\�`�l�E,�T]cc�ZEs#nR�_���]�v���m�g���(�o� ��2��8�߁�����Hs��{f��a��J�,ф.>^[ލ���ć�Gf;�yl��k[`.�34�y<�8����Fϓ�'�>�Y��T-Sͤ�C��*�>�����D��xv��G٧ �M�k�^���G5ZE1ҒZc��-,*xƂd�7�k��� qv�wz1s�թ���O�T����`�B�0	��`��Ε���V�&O�{��Z}~~��8��60���.^16>��}8h�˸�XP��\����->{,��%� /�I�F�]��A�a}wt�10�ݭ$A���B���~p��8��qt�E�� )��(�w�I�HN2;؈�	&!=���`�����$5ʠ��R"]��xM��=��*q���x��O�o��S1�U���ܝ�z������s��/\���"%g��
�N;8!��^~I��mV�^C��W��@5��ej��@ê�{���֫6HRt��B+a�tցPKmSAc�;�n����p��_NAhO.�T��֏��L���UUY���E^hQ>4X2\9�j�5�Ep����vn�"w�J����a��p��-Ɋh��%DSX�D|E��)^�wi��YV3=e�KzH=0�Z3�'�a���`g���S�F�<z#*�pF��4�	��wNA���g�WI�o�j��a4�秎� �
fu��وNc�yO���1Å���dc�:��~0ӣH�����'��m2�633�?w��Mp�c�X��	��B@�պ�2��f���\Q�}5ޜX �g�d4/�y��ґ���	��9��ˤ�n��T��w0?i�������Ryz�]Vq�SK,��'�F���m�2�����<��:���"b�H�6�Įb4\���$a�y��୦gD����A�[�R�3%տ�����:��>.�S�]_�?���P�Aģ�S)�5�j�����Ӱ������Ղ�*ǥ��⼘V'@�XBD1�l��1$3�6�o�27d��~0�F�D���4`g���h����0�V������X��\�I���"��ڮ�4�Sm�T�)r��]�.�W��I n|�l�yN�J�'bs�qڏИ�.+��V{`��c�(���<_YUA.f�Ӏ�#f'r�u�ό۶6oZ9qi|}����$��k������?X;s��w�q��G/����
�,�&��Ahj�a�gܜ΂E@u9q̼�5�Pܳ!�"[}/V���?���P��;�����Q��[���\�G,��R���UK�af���x�x,u�8�Yk�e�XI}��5�S��*�����zy�Z�W�s<�cGF���D�b"��`j���JM�����0�j���9�F�|��d�⾂v�x/�<�ٸ��t�#�;Z��Dn?���`�[E,0�*����H~��a�;
LN��L�A������e�c��f��/J1�q~t�Mmq�1�9b�	`b/�:���SԺ����:k̢��!^���7��b�:�hgN��L�Ja]U�o�u0��3?;�)�X�K���b&��3J��������1~a�D5���dϲl�&�5�W��G�ާ�����E� l"��z4��j��RN�(�7B��!���
�9u�=bv�Ux��FĿR/mu��vu+M\I�|[)BA#]��ه �&ۧ27!E�6t����n�����!�mDYs�T�!��J��g��ґ��ekId)�6�H��i�5\7& ϖ��s����w&6Pt�J6����0\ڮ�\�]�����l��(��,��U25]a;�]v�[d=��g�M���'��63F(!�0s����Í�Ya$ם�(�8�|��edi�w7��>h]����G�&\��aަ0��0�qYo�4�?�UC����K//���[9ҍi�2y�i��y��n�/\�82B��o?�/@�����?����y#��kIrɋ-3���N6���vXC�yJ�%�;x���)a�x��w�x�M`|�\xŁ��c%�Ϛ����I<���O�"�]�(qtܣv�E1���do���m��K'�
r�@
�{� �>d+���j���ir�^==���h��Y��2v�V'.�U0@2�/ȅH�7�
a�h���A���=K(oqҶ�9Y��sbh���}4�4{H�Ր��DQ>���$�ģ�j����\���0�ƾ�r½��#�,�<�6�(8�BE{uT4�;v�
����Z��fI���r�lg���7���'���,������W����)HUrQw��,�N�!�I�=�r�T@�+d�H��Ҿ-olq�� �pi�.��4� �p�yM�SF�ܳ[��ly.���B#XK.~���)��m_E,݄_�*Jl;⍾�u*��$U)a>�n�0�ͭؾH�d�*����t�D��w/�w��zR�2m�)�4�_WWަ��!�b�<)�9z#����E
}R��΁Qh��[DI��$iw�V�dt�ߠ���D-3S�������=Xي&��k©��	Pځ#��@h+.��ڇm�.��M8��R�?;�Z���་8# �xfpTA�+-:{Z�)�����#oռ�>�����'��[�(l��N�v#��@z�=	�t�������]~��6�P�Z�)����� ٤�J������7Cܞ	t,4ټ��&����y�r����1L��X4gT�]�A���'�7AOu9�l�o�ֺ�g�ǃp5�����4���!�v �
f?��k!U�x9��W�ݲO�I��K��K9�%�H�\���^��g��:��	P����,�)�b�[�N|�u��H��M�6ԴN�x���2�9ܺ�dIKs\i3s�k���d���f�9���fm���1�������&�
�$(�+0#U�e�
�iV����&���Mi�C�x� �(�H_y�2ê�֦h��
�He�z�<W�i�j��6���U��M!nQ�[:������o���po�+te�K5��|5��U`���F��F�=z����d�L'j�T絀"Y�ȏ�}� =w�(�axy�+&��7�Ȣ�i���>��TyPZ�׭P�	�O&L�8f�:Ƕ�|sk8zy�I_�R�4���3�Ȑ},X5kơ$��d���M�R����Hb|�7�۴͑��~X<�ݍ��H��(c�y�Mߡ�D����Ū�,L�S�IOIO�9���I�����8O�f�Jx��5
�j����agO���K7Z���R�5� �o����B2U-��aW�TO�˂�+e�$$�L��䛙t�D-d`��}��Մ&��O�u�^k�&Z��\N�'-yk*������	�b�J[�Q2?.8!v��JYo�!�������yy~v����ZhDp��h��T0��+��S���%���nd�yD�񳖿���@z�{w� �`=e��a��� ���8՟B2�=f��,�0R�R��o��sO���M�t
� ���L����L�>F������hX_���N�Gԧ�g�k�+:�R��~)��i_Ue��Ն�����'s��0�f�k]f�vȉ;���x�m_��r0�K7�9��|�B5#zGMqb4Z���c��Ǣ���SZ���'�`w?6��d�}k�"j���T�|��:]
=���}��-'K��gOs?̤)�ڎ����F�=�lj�PIx�a����eBW�T��5����r��M�P�	I��>��id��L��ԲKJ��:�Q���"5�Lc@�*/l�\+���%�g��<g{ѕђ���Lˑ>l�ܤD$i�Xݩ������4�g�`^Ў<���X����оK=Ws������֚T- |���${�/ǂ3^��ΟB�W�D������z®�}8�`�ң�݆.Zx�R�J�B`� �V���J�E�A��Gr	k�sl8�֨�ӭ��DD%�C\���^F�%�8%
��3���fN����gQ���� �r�<,���%�K���GI�;כ4���"��<L�<S�3�A 9X�3��A+��6O � �I�hR���[X��n� B�'�Wͱ��d&��o$�ki��ͧeY�Lw&e����>��vX�A�	e6e�|us1/2e�޻�(ݪ��ϙ�Z6�͊�-˺-�Ű���~yq����H�� �Z�7������^��ID����T@y0���T0%���J�5� sZ>�/�'��G]�Zի����ƈ��}KE���ґ��ϼɂ��!��2o��hj�&��BO��>x].�4�
3mO����*��	ө�"��R�\��f�H0�������j���E�?��Na���qjK$~�nH>v��a[��*_d��SSW^�ar���a��{��6W�P~�`��8���H}h��3OO/�����h�6`ZGU&6i��3�AS�b3�h���v���WL+��
%�J�)I�������⒇�AiLQ� �����-�i�T40�2��Dڹ�թ\�2?�yw3١2O�k��m��E�玲SI^�|m���eX���l�
pd�5��~�^Zu�76Al��qi��<ԛQ�/���y�k�*���$���Cm�(2�  �X���\ޖ�����֞/��"�m�4:���`�B>mK;oc���n�+������\40�:�	[Гw�(v]�Of`\�4��l�dK*T�h�we�|N���e�j���+]��<ŧ"�ð�ʉqB�v?��G��ͤ�?]��f���S�#[x��Ĕ���،�W���{�)M�����-�O�Ȕĭ%"u..uX7[ "�#��^���*DO��yS����UF0��:Lx�	S��-#y����5CXP0f�����nq�8s9���qQUٯ̘<U�;2��T��?���#@A����q��씛Nr��|9�6�zg�bd��K0�Ŕ�
�&����L����A_	�����,��S�T	Y���(F>~�V
s�*=�$HN�y{�hr>ULK�%�)�+ټ�d���0^9��ʾhr�!uC8V�
�����!Cu=���������!���ۻ��mJ.�XH�4���9����k���lWY��@Z��Y�pOv������������~*74��+�F�*���p�Ȋ(��"[>���x0�l���U\�^/�Ǣ�	$ �6.���9��h��ѝ=��D)�d4������u3���ht�G�p��S�
h�'�R�D%������Ly�:<;USO�t��L׌�,�'�������>�7݁S���1ќ����� X_ř�d�`��D`K���io�*��;Or�����*>�v+��G�`�����Վ1"w��%��[�X��;3�,5b���X�$3�,��i�>�#�泱��A1��r]&2i��� �:]L�d���9��,
�Ʒ��<n����l�A�쿾�|������?�*�d撏�s}��	_�ڑ�NwX�w��"���h�0��c�Ub��1t�W���`��ͤu�-G�|�\���tng\��rdP�6x�D����y�F%�g\�V�ʿ���,1�	���;.u,7�PÌ�E}C��=�ϰC5o��k�������8���I��.	��{�ƚ���· �,��a�Z)�R�¼;P����l�si]�,��DX�0:�@�>�m$��y�f@P�4J�^"�]���X�ݜE6�@�d!�<��䗖\��!���.�3�����k�l~{���Jc+e�p���G��bޝ��½X�`�P�3!d*)�?�I�."fk�X�[�VA-�\,gRܑ/��W2� n��">֐���~MH� P��� |�1����u�����z3�&/3n�:�\|j��3�I'�/ڒ"J=Q�4�2xX�]��E�P`��Xp��0z�A� 8���C���{�g�FH�2{iaZ�F��[�-�K.��G�!-Z���=e��\J��5���}�0-��h���tE�	<�?3�b�E�V����y��]�B��'��a��[�W�9D�8�l��.�������>�M�����r���*�"�;��r��1���Ε/��M|D�8T��cd����p�G�'�Y��3!�k5�/�F�a&�NIY�ϕ��3C�G��J�!�o�]�%b�P�u�+�̚�%=1kl�����,i�&�x( ��?;b�Qw�^�E5��i���ڭmG��%��El���w�ʿ=Xu�>�5W_H>����_���+ԍb�hRr;��U���p\mj�"W�DI�Iۄd��Ai�����g�X������w�Es�Qa}��$�MR��"�ol�(v2�ϰ�/U}E�C#���G�.(�)��G��U�'P�H��b����.����0�/�|/�N����V�Ú�'9Xt�B!��+�����5
��ʺ��ښ7,مe)�� �����3EQ6(�,��E -G�2��S��D��F5�"�[K&'�H��p������,Ce��*���xN��S���`�
����.��� 0�|��>����	|�d�T���2�m���R�T�3G��+��@���=B�ؘ��!��G���A}�V:_����z܂/�J�坯��W�)�g�>�pں������&1���c2��YO]��U�y�6���jTu�Tk�{�s�Qca$��fhQH@�C�e�>�16CIS�&5�Ӭb�T��s�N��ھb�w0�w���x��}]�����m4��F�Og���*)f�,��rA��>$�.��7�3]���d�yl(,)Ă�6��#͂�/���?�ާ,l�l�Y��PB�xإb̉��#d�h��?��"�3����)`!/"c�է�q�Knڊ�����&Z��#.��3�Ψ�(���c�s��!-�G��8�J��e�e����.6�m}׽xvb(?�n<�*�P�OK�ޯ[ ; lI��[�'% F@���zS��}Y'6x���5��q����C��D��>���y<{� Ԏ,�ʁ���U�Q/�pD����>����j�⮧���0LH��ʾ����IC<I<�i��e��X=�g-䎒�FC�]^5"n"���b	�0F�-�:~�s�t֍2=yd��^���	�!$�� �����a��Q:u����t?6���>n� k�5"��'�6u��!o~�U�8d��H]�`�
��O����,�g�-�����S�A�_�23�⍊ �6�&kB�-K�	=M."@v6�<�n�hI"��\;���'��r=�`,��.%:�\��Vg���R����@uf�(R���<�P��V�x6���D�XV�1�4(�v��/��?1��m�?��]_���:�N����L�BЬ�#���/Z��(l�ד�ؤ/=a���%^�]1ȺUU,�I���$zQ�IGn��lO���Pз<(��J�z� �S41�(g^�a ���ʬy�����/�zL�q^����x�']wǌMrD;��(黍iώ�D��Q�W�fE-����c��CE��8N!����{t*����ɶpv�������>}��#�I��j ��$W�r}j]@|!)8gn���5ݐX~��c�\��U1�4e� �:l�� ��'0�,�3S^��N
����������\�D�
�reL]gV�el��A��'�����0�(N���Ό����]���/�D�$��Zw�#R��2�;�=��V'f7���cB�H�r�
 R��Qml<�/D�F-�7����%Yk~�̀=���2��EF#�g�cY>�ِ�Yr�	�j��V��kN��W����,l\h�@�)�p�t	z���k�;H5G|wagg���g��g��\y>*�������χ�ޮ��^���2,l��k���pٯ���#| �ɖ(㪹�~�Ma~�$���]���'8��ɲ"I���(/�v����WW��t��'hc�_m(]q�M2����)4����:)�q�F��f13����(%A�$�lp�,��{����4�e��i�����%��V�$��Q��V4|Sj,���JV3[x<���+��i�z���ilhH)������c�8���/�Quo�K�`�OM"��~��h��n�q�>&r�o�H�lS��)�{v��:���h^�4� 4\�G��3��Bi���\�Z���.����j��?h�;n�x3�iWp�E�}�2���G.)�%�q��4�d|�y����/�)����>��3��Vմ��m��-I� �{��a4=I]�y��D�(9[/M���'�'�<C{��>S�B�Rn$��,V�:�.t����+�2Ô�r���A�� -��k�>Ł��K
�hOM�P+�GG�����l��gQ�/���b�h���9��Ӹ��x�{�"��fo�s�7����\	��j���lEn���B��K�p~<��"�9ݯ��s���?�2Db��R�A�*)��"�Hg�����j`1�x�X^��� ;^.���h��o����d�1���]/P��p�M��(�B�u�S������Ʈԓ�~d������������ s>��nGɭȸF�h�F�ށR�c\W�C[�����y�v���ƽ'������'4Џ��f1=�-AY��i�~�"�H�P?���$��X�\�P���.^�l�B_����P�Ʌ�����rMiD�����Z��į�`^\�|4�F�
��Y+;K�OR&�����d��n;��=��#�t�眻�t�
��PU+����z@?�v�t�ǦO8W�s�h��e��{�����Fw;!�~	��1֯r��b�\DI�^��?O�:To�4�H{s1&���\����_S��>�?8s�U�(*�%�@�u���o����}� �h���,k�Em��d7�d����d�,�ky�86$�'�@'7�U��-����H�������
߲�L����Fԫr�5E���0\�ۧ�r�!%^�ɏ�n�Ȏѣ}N��!0�o�1�ܟr�o<��113P�>=}��8{�g,}"����6F%*CA
��"Oݨ{��@��qd�i]��_�~���U�4�_��P�4�|H��O{]mjPF�K�r�(T�T��H�vP��q�|-���`W:o��D�܈͉���o��z�W+\��yN��e�x�_&�q���o�v����:�=��W��-w�{��l��lņ�Ӱar�"�%B����q �<>I�(��	�ޠ!����i�r���nO��I>�W6یn��fnV��bމ:5�_n�t����������jU<�_]�V@�Ca����y�UIx��^�^�D���M⤰�0h�G g�X2S�x�<WZ�x����T��C�r�x�r~e�F���M��gfM���`<�����!m~|��M�R�.���Ȃ��U~���܁������:#�~ f�*��3��S�_���*�IE����/�����g�5�xR�����B��q�lV oHg'�J�Y1� w3�&%�����w{IPo�d{�*�`����Ԅ��^7���\�����/ŅwXI� �Acj����tV��W�1S��Jx��Q��e5ys�03�������@���*Y.��3�'%�JCb �7��E]�������pNAs�r�|��F	v�DƘ�t�D/�'G�Z�MM�:R��P��B}&��eI�Q�2J�e����ķV����~,Q����_���u�4�0Q"$��>�.Qt�>N�)��m�NV?���\H�]�<�����ܩ��-�رsk�������<J�\V�Ĉg�O�J�ϕ�Zn��[*&b�&=�Uep*����Fd5J�������gʅ1i/�\.Ի�\������)�e�/��� {B���,�+�SG��z��*Q����Td��=B?��P���n$Zn@���T�X�9p�D�mڰ�%�'�k"�q_�p7Ȯ�C�RKڂ�����<�v��A}5!%|��+'7a.��~���9����Fcr<[#k��s���KzrsP�t�:�1vu��&](�D�:��3�dF��.dz�ۨ��4ʈܘQ�D��x���B�@h,���(4*��LS���!��n������ҍ.C����d�<�´Vy�QOx���<eô�*�b���Z���G.0m�*$~,[��s�ct�z�%���݄�4�e�Jb��ȱ��?���A��C9���Pm'�!�X��a9EX��	�QRb֙���=�9��|��a0�A�E��]��i4b�}K����wN��PW�sܩߧ��˫ЀxVۑ�W���ᑢ�#Z<��@�B��_�Ļ�hL��[L9^K	L�u�ޞu��GGw5�����͹H�q�E�0!�b00�t�@
'23���mV�;��DS�J�7��A����X��M��?��jy���Xļ����J��:���2V%�Ӡ���K8�N�b��2�6])�A1�� d��3�P��F A7<kA�d!�KК�D��R���h�I�ih��E�5�mLWkt�;����4�� ��dsx�9�n�7#9�ܾ��7�%��3 G5g<�ʐtR�C��<��2���$�%H]��H�,2���ə�D�_����,��1unA�樴н��5@
Is*����`�]�=�­lW7�c)*��J�ԣ��L����Hy~�}�:�X�O� �~$p�2�Y���r���T�!�.�*b��� A.dHd�\�5�[2jAZ���T��􌰕�6_��G�����[���'�X�%�HrO��L�w�*|�7[�Ce�G�����*�πA@(���NN�8��s�[zZ5��&HR�4(��AK�?5n�c���?�@��$<y]��<�<]1��zF�;J*��gmr�$�Y��� �Ƀ�g��41q���[ڠ�(ª�l�c������	b��n�p��vS܉Ou����􌉮� ����8����~�}e��R�nc6[h�V�~g�Jq�{�DB�x*���0t����V�k݋]�����N�/>��w��̝O����^����JE�b�j��U�ӻ���KM�ӈu��(����j�`8rv��"e��N�G${@���=�ߤ��͠0��w��׉"8�<,С[̑�ؼ^��}a3@w�eb�v�;�8`!B��l�$�Q:��'j�_�/�R����OW���[���n3�����ULb�aO�uK��	|��_�\���H�0J���ð��	R�Kf"8\@�ǝ�o���4�"b�*�N���?��f�g��������o�ݚ-�I���e>u�vBה_�F|�� ����L2�w(���)�T./@�k&����J�s0C5�Q���D��.O,���h������O�1��r˹��jU~�y�����ߠi���^>��Ӟ[ĝdwY	�.Ɵ��@����b�q�	��`����B���1qb�_$4���頁���9	� J�'���������@ L�mJY��{u��Qߏ��X�x�]Q`�zj����G����Ff,���YF��,VL�)A���E�Tmn+��n��崸u9��B�#C qH������wi��m���/�d�U/�
U�q�>�΋���b?�0r;)k��͇�O��\*���4Iv��������d�O�~<P�Z�h��Re�!Qsl�7���qK�h��4����z��	���rTŀ[a�G����ռnP��z~�Đ��|{�Eb��Ʒ,�����C �Ag� k�ق�n��f�g��nǹ����J�35�����1d[ԣ������p���*���*�F��[�&�hl����:��q�,C�a��P�J7M�p�5��~���Qoi�ҏ�O����ôBAH�opާG�
@i�P� Y�i.�>m���U���>0Qf8Q�?�Hg ��S�-�b��4���&�JӓxA���\���``[�T��"^��r�[���3�<�0�{�H���KVh��u���ˆ� v\�Ei����IiJ�!���s�͒�/y��w���ɑ����Ұ��f�C�eA=;#uf�w�#x���ȇx��0��V+���ԕ��#-�oO�
Z�K(�������J��UNٜ/�
j,&���	و����_���]�+��L����讐��Q�ka�^��;&o���{3�8�[6p ����J_���G�ޥ��ȑ��|S1�)x1}qE[��в���W���.#3Tb��B'.�b,Ċ�y���C0bg����(�0��Nk�91�ռ3��/������1�H�@�6����JK�Ca:��k�J��F�)E950�}�,��^6������7�&	�خ*��*ebj��һSy��}�7����[������tV�*B1�?�� ��_���ʼR+��܃��ZWL�C����L������1�Qu����)�R�[" �1F�57���Ex:_�щ���)���bC�Q�'0�dU�|�~6>��v�����#��!1�V@g$�^<A9���:+%�C#L�j�bQ���5|�U�o��7��r'�y�v$LT
9�'�d��~nNڄ����z�m<?EԲ�1�2��.��x:�7��2�-7}���6�W/�f@4��@1�S�̩�tDJ�F��b��������73��t�A����~��[����
Yַs�� �D�3�֘��q"���I����`F�z���`��Ҽ��)6�[D���;Th�[��"oج�}M����L���π��}����,�d9O �S���ǡ�Ƃ�|��)e�}��BNzʋ(Ll ��!�SZ�iWt�����ع,.��T1��B��^į���;��C2�P��$Z��y7��h�5=������5k~إ����QP����B�X(�>��j�V;���u��Q�t�"��V!��n���nZ�x����~�׹��;���P�-}s��5�Hы���	��d%����b件�l��X?��|!x�/G��\��Xš
�"���� j ?�����|��(2�}�48\v�1Rppy����C�z�q<��,�0z{8�R�wDt�ٳ��{�n*�+xǇ��n��u�5�D�X����V���`�?��h��ڞ���T�!�(�P�1:3�E���Z+�)�+�GQ�b��Oīt0���槊���S)|�<y���8���0���[8ڕk"o��e�Dj�����e�(�"������z%R�G�7 (��n"���g,mj��AM�G�`�0D3	���%�H�7��j�VH%B	�z_7UҺW�j (��O' FuG�mo����j7KZ�e��(�W�^@�w.��\9�墌��p�NX�z�y}ፃ@�k�F�����Q3�|��1E��]*���2��|���#�?���V�<�x���%{)x�c�0�w)'C��:-x's�E�H}�C��;�rկ�
O*��G��%�R�� �\��YѪj(ř	P8*i�;X��*�v�}�����Y
e�Z�N0��"�a�"������\��4�9�,d���k�E�e���g\^���$�&�+��4p�u�����C�JoyU%��n��&�r����Ef����X�f��B��	�P#��Բ�I�ݒ ���U��t�A���Y!�;�/*$D����Mz��nD����C���,���Ut��l�<!�=1���T_:��K_���0�����u������z'���w�\�����ME icjj�<�lKhJ~%�r��BHH�N�1ɨ^�5X.��W�R���<�lBN�p'���l�� ��bb&g>[)gW=	g�4����e��p��<6Z�^Xu�޶�Ly�"��1��18���6�a�Z�l.�P'�a����)��^˔AW�v��~T�
d,Vxc��0p a&�a�[�,jS#6%�OJ����-{Ȧ`�̶��&2o��
tG��i]�U-�e�������G�f.����9���3�P��� TxTX�Ȅ���[ٻө5��Ѻ�JH���.���b�ìgSl��=;B^��%����US5�K#��"*�P9�4d��d�?���ȑ@E�Vr�Di{h��(��e�`%��j�V	P؊�����@;G���!����[����j�f��A��D�Jn.uF����'����՜���$�of�<���|Dԋ�7�n�����}Mq���t�>��-�|�:�?̾�qosC�
X�9;���x�m��:�4�K���Ϛ&L�uh�p%»x��:d���d��@}���kB"Ę|�qn�֓�O�m�t^n�����θѴ��xf^�-�����eN�n+?g��K+��2*+)�;�#c�J"�W���
0�s�)t�g����fC#+��)9k5T��6V��ӬM5�Ӑ��M��޽�r�H_)�'���3����)P��1��!&��&R�%�|��`�b�}�)e��Z���]Mx͢�q�l���w��f�VIy�������5�� ���w�����������r�2�I�wc�K$��Ttҟ���a�Fu��d���=�Sx:#X��~Kwt���N����ʄ��.����f�����Q�b�n��?��s�q���	CZ/��gz:i��2���3=r{yf������V�����i��mMW�{Jj�7�0-?�r)atY��{�
���B�yWA)n�-��X�o.;dU�6Ppq�4ԍ���婡��� ���$L|R�nu<�@�R��z��+�ʐ�0<������W�R8S~}쎺 ��G�ņn��Zpf	��>>��R)wTj13Ǹ��߫�����j6�@) 7�i��5���U����͆��#��Ț璯���cHĹUѓL�*.+��O*�;�!�4,Ig�J�:lBh��<����"E���i�e�N��ԅòy����/����I؃1�Sy�'���ϯ)��큵G���8m-D��v?��������q��t#zq�AP��޶�5%��k�G�4M�˲��X�ό|���B���o���M��ѪЁ�b0uf�D�LB�%*ao��1����xU�����#|)�u�ҏ��>)��c@v;:�h�N�s�_����|v����-�#�ء#����ť�	Q�a�Ԁ:u��O\����������$��[*�,!�y�d�G��g��.�͘��¼]F"�󞷑��:v�a�-Cp�N�0XY�[���Lg���y��>H'������3ؙ��!���B��o�z��]�\��y��q÷��OA�#��:����ᙘ��ޤB|]�U9��>6E�o�Úg���@�w�.v�"]qb�t���UC�h� �1-G�)Cܯn�Y���6��`Ms;bEu_{&���(�����ɨ�� �D�C�8h/�MUj��s�96+���vTwy�?�	_���pz��xS��p�Ǔ�8��UGm�p�O�WŻ"��S'iϞ��j���Y�c�馭�z��ҭt�p��>c1�8�[w\���O��U���Q�W���8�:�:�������rY�B;}�#�M��&- �n>�۸YFq#;^���WeJ�t����-��>)K����+� hZ��pkX�z�<r��K��r��
���=�1k��b��"
$ͯ��ͼ\_�S�ѓ��N�޽��q�4�}5�M���b�#R[p�C��j�u.{�dw=l� �7W�*~&H���Q1��� ����Ү���!B�V��Ak����[�a��4�A�[1۷�X��)/}���E2�#{�D��ӿ.p���n_o�]p�Ϩ���{$gI׊s4��j٪D����ecx6\[6W%L�kfify@��Ϫ�`��_U*�FBAg�E}](6�saB��Kf�`Yb��׎jDߗ;��O@��_|�s�6���vf��(պ��^�y�`-�M�����oz Q�7���x����YE��޸�zR�&��|�B's@����S�X�Е"Շ[�Na�'䢸tHo|H�3��q�#I��8";&z���?���~?���N��i��]mz��6O� �gh/j,�v���D��:�5UQ�Q��@���d���9>�u 7<�����^Ώ���+#�qh�_pS+-\8ώ�bE�N��"�{U��u|R="�K<Ix�Z�퀲QQ�J/����)|����-K��~�d�yw�d��1~73���6��!2��+g����j��-�'δ$�^��B��2��a�6�=��ɒ��+ܮ�u�❵ĕ���)^�\L�wH%��k���Z�D�i--.�(t�Jkr"_B���m���?w��;�}0o��>N�P�}7X ����+�`���T��X8삩��]��&6�T����|�g���'47�R�f|{`��c�V��V'D�k��<�mh���*K��LD������֙�%��� q���Tc��sM��N���]���OHN@-�bǰ�mNx^w��e�^Q'6|i���1c.���~8�/XQ+��B�^h���x�C9��ye�-9 ��N��`�R��Qcs���6%Ű<Ln�X��<{� cey�h,C��UUD��>�{JzTU��fF
���H���G`=ɠ�λ�s�a��}�c
�8��
��4��^.��.��l����������t�;�v�c�MY�+,&b;�YmZ��D��Y��!�0h @�_F�H�~�INԩBvl����Ϙ��a����h�slw��Y�YM�l���U=7G������2��oS��Dp�;-YkW����3SS��8���H���u�B�/+x*�!dI����uҝo��=�b���<i�/:齙�KY�5�w�~����*��9��i������ڇC^�Yr{��#�ɳ�i؏|�N���a2>Al,��r�a.y/\|���e�(Li���ό�ǟ'6㙐����Z����h��7��DU��������!�4p�U""BlXi�n0v�*bչ-�EV��;&��H�tfc���M���.�C&mVKF7v:a�=��~�з��V!�����n��kfCA� �Z��D��w����г�Xuf�~�� �?&�Q����E��\t�����d�8t��@�D
��-<� �(�b��`Yp��&�����z��l�ԇ��{�&�Z�czu�k2���jOb��9�H�J�Q"���)РR�Ш��&���,V�Y�>��Y�nh�Sn�� 3&	
�������(ɀ"�0��W�r��)B�7.�6���ggZ{��(��f뱼��
�3ǏM�X@Jӓ���Cxlx|�'D�_$��`����<Q��S���Y,�"�*n�،,#�g�y�Ƌ��* P����WO���#�P���̰��u�3�54��=[�f+�gu�%c2$R�����'��JGo<��4�ݸ�W"��c������ī�w�[uG#�P%XmK3�]����OW���n����8�4g#�i:��^�.���?�D�)�����W�A��D��b,�uM�5����[o�SC�~}�0�X�<Q���~F�%�
�MQ:�;��p�o���NFͱ�GL#s]�S2Oc�_j5=2|=([Ugt�2f�L�/#��Q��d./<���>��H<t��_�0�T��豙+>�Xٙ�v���!�O��Fs�#V���� Ҁ�Xۋt���yj1�����.kbp�.Tu�<�+�f>\v���.��������g$��ώ?,�V����^�|=Q��#6np��vHӴ�2>�n�Q��ng�l���K?��E�0=hS8����E>��S�(�����a����4��(O����m�?�r\����{s�iٶZu�X���X��i�o4��8	8
rr8�&�9a� ԧ)]���>6&F�XH�.��(�,��w#ޜÚxF��8�+��G����J�Γ�Qm�ݦyB8h�����A7	Mܠ��R��p�)���� ��4��Ae�\K@�$"�b5�-n
/�Pkh/��(_�x@�y+�	oןML��5��y�l�щ���6>�b�܌�h�!J�7�c�ڶa{x�r[�K/[;Y�,�*�\i/���f����ˤ�A+w�'���R�!�^�^IҊC�m�맸\Y�atM����!-i��X��W�d�R�7�-�	��P��А�ub�5��¢j���䖑����~A:sI�sCe>(0����O���CL�4���F�ȟ�`mY�_�m�S�9K}�֤ac��ȧ��l����j���7�!Dx Be���e�`E�2������:?��5Ւչ��+KD�O�=1����TLȏ-!���9?_�4"�03`K��H	Rx��������x�w<Ӥ4Md��@��4"�o�۠O����i���Q�{�^�"g4U3��Q�Q��~�b�Q�FK���Jh����"2�*����{�h�?(�%N���h��8����2L,p$��f*�d�T�S2��o�0p��X<�)W�7��|�``x�4��LmXsT���˻׋���R��|T���2<ډ��� ~=�|[�f�E!��	�L�T(����<9
L���v��(bևǁC7�~��^NԾ6�<yG"�����SQI!*7��)�/n�DS�	�G���$��"�&����/�W���,�T*��b���]�&F�0����X�(Tu�"��,]0�ì���y̿{|����R@�p"��m�|���s���sb��F/���@��
�|�����-D���(�MZz��tP��!#��_���m.ʦ�ΰ������0yu�v��+ZjƝ-�c������)�P�7
c���^�]��7  ���#�i�[�狅�ph�+�YZ�{�Y$S4|6ј�����H��-�3 ���f�%�[�r.dGs��Ų�>�N���'9���}�7g�g��j��&q�g�3cWC�=S����^ڋŎ+���@a��/�$#p��ǵc�G����9����)&�أ*��i�5�8�̥�u������YA)�4�5ǭ�⅄�=�g/�(|N�r�j�5��y��*����<+�4���Z�/3���e&�Ę#"��5C��^�D���4��>D��N��Vׁ!M$_��Ë�#�J#n�dd�i}�(tf�l۶�V+��AW��şl��
���+)m#*͵͑�)d�@�@z��o�>('/:�n�Bn��&�D���，���f|�3vv�јB��l����F���sh�_�=M����>���n�x������M$\�Æ���i�+<��hSbL�D�T;B���]�X�Y*�L$���%3�W[��B�gl"�cd	D� ,�>�w@���mDC������X������ �fp��.�C�d���!���/n������+�u��E	�!�������.�D�ʙ���D�PE�����|P����/̺�#Ym�j.��2�����T���'I&�I=�0����-ҷVL��_�E�kr��W]��&�6�`�+_��{z��Mm7R���.hH"'�"�4�v~:j�tt��55���F����0�:ڲ�C�Ip�N��'Fưl�
T.�� 3w��%P�+�bp��Z���eҐ�l+����dz̰�$u`�����)ltn�`oo%���x�W�B�
�:��� ��=��@x_�� ��C��嗍p��	�|��R����eg��/�d���xTD�[������CN����p��j�C� 2x��I�b�bOV�ݛԃ�꼑�����I4�{��/�S����N���X��W�q�o�?L�Ԁb<Ŕ8�����8����������~���܊���P�	/�|� �?�7h�`��7��4h��{��tF�%%@�P �4��{B��M.��*���c��rKc-�-�O@J@�b�	q��}��X��ͱ��K�t�"��m/���2������q�=��QL��Tj�r��f��G}�;�RZ����I&l�3j ���Ov��F�@cNmr{�#r?�r��_d�{���xb����`]L��|�)̌\�9(�wgB�T0Je''R��Ӡ�£��.�(���V0B~+exhIw1�xP����'E��R5��W���=��@�����踾.����e���m.���0b�o,Z��Q�{:��(Y�����f#���N����d�@��3��k� �
9l�S8O�ם��ٿ��t�Km,���U��y�i�^-������:ʹ��g
�nMok�͠{��P=�in.H5�_��	�sP�`�q,��SܽDfZ@�H6%�%�`(X�E�nT����\��ۉے�ۗ����6gh��̫��g�~��kڨw�ᗗq2pκZ
��R;~�gGS�Xy�Sg��qD�1��ޑ�e�)�F�����N�E����{�ϕ���w4���o��������� Q��&�~��Qq; ����p��Yv$0�9�l]q ������O������gN2�M{6�ٙ���9�7�.r�t�d��
��	�5�K�c��R�-G*��pK#]�;B��!����Q��`�8�/ݏ���K�B�������r�f�9�J���].|�$�:EyC{騶�e$'��ԝ�&N���o�d;Ԏ�
1���v��K�J�t��Z��|0����ƍ�C�c��Q	��0g��ˎ�&�6`�2�Z�;G�����(Jr�ϛ`�rGD~�W��� �9�,�Ya�/�kUe�]�0�*~-�xc�$�L->Z�k�̰�h�W���&��s� [(��,�e��N�u���#N�h���T�������Q�����d~��h�F���$tm���?.i���:���JD	ú&����Ȏ����MW�������ΜF�Y��a�?%��o;Of%�u�/`+�:nm� �<��`R7��~�v�_��j�8Z/��m��a�X).H�&`�84�� s�k�h��v�X-)T�S�LTk5b�����c���WLE��b��Wߛ�U��!��$�S|�m�^ykw����#3�l�p1��{S[�����DD�3댝y��x^�A*)��D���zD�Jp����?F	XBÆ*w�-@91�2��j��6�:G������4��I��.�%_%�*���<��v���1���>�"�w#�:�!�����󕧌�]�vR!��F�ed<�j����?���=��7��>��+�-P�+��2��(J�r��z|�,vD��`c�x�l�:��(ӣ�'��a^t��h�w�����'�>m��V����F;�n�x��`�E�@�dq����Г��E�v,��O�e�^�ρ�\��I=z�A\�-�?ǜh��_�y���G�W��D��MCy��̶#{kϢ%iD�bf���m(-Á�߂�o;�Pp�ͯ�,uG P���z}?�����/�x�Wj�w)�%,8@(?$H��2c���1�E��g!$"u�g��18믍Ƽ377�!Ѯ�J��+g+Zj���oy9hje��^N��X���uc=����@ ���yT�弁�B�]Ж�[	�����J�,�b���i����e^i�o�������붿}�f���ؘ�#Q�<!�ܭ��V���9	F�Aˋ�C���,��ZN�	P`<�8�������]4������w�{��^l��RU >�z����cٸ\缓����o\���b��;�|Ra��%��/���d�|�1�0�K�@;d㨁�'�.�HG�t�`�`�u���M��pW��˯Ô#rNC�
�9OT�%��-��*������B[� L��XM�ɜn?�F.ciq�����1�yB�w���X��U���E8��tR3Ƚ[�x93����.�0m�Qt��LAd=����%��WD��;� �ȩ��*�����?�DL�o(�^�3�f�N�PM��U|�9}-X��>d�ݦU,�~[@1ǶZ���|b�⿫-|f���e��"�����[�1OA��V_C1;�,7����]���sZ�`k����-<2��}��%\�6�$��`b	��0�w,d��n�����jBf������!��Ɩ�&�%��񗴔����0���}È�^�ԅ����Z�����^_�~tJC?<�1��B���AK���b�p��]�=�*{��-C(pa��LuXz���=��X�i(.���a���#�b���?�_q!ף�'�_̎0��0�^�d��~�43D5��(��K���&��<S�QN(x��@yf�M]�e���+�M���Ӷ�uO�FN�[�	\��.��kB8�=��tr�T�eIk�Hs�N�]ʢ�K����<(���M���>�燽�:h�w�Z8ψ��5�=�B�� &�q[�";�$��ͥ@��.��o�| ���w����ُ�a�!��Fk�ԥ����	�H���{k�"�5>Z�18C'���|g)>W����F�=j+S�JO�4���}�Y�Q9�I��QUE(v���Ǖ2*�I�����<`��ҟⰦ
0_�k�:"��`�*�_QC�~�Z��/=��ga��7?�f%:_�"{�J�8��Z;Wi��hۏ�Zi�۪��F�"�!��6�f����յ�=�
3�F����7���7����5�$Ӝ\,�x)�Ê)Q3\��uX�;Jע�D�U��u�PWa���sN�9���}{�}wcg�L���P��$Ē݁H~�$`��BR�n�Bk�S$p�a�c��ު����\�=���h�_�[]x��� ����<�zL�\���	���s�lN"��� �\�wU"eR�ƀ5��[W=\�U�l�[A��Yb�O1)j�tӜ��17J��SBj�W��P�5!��[�i�R���ϒ���{𦻪/͏���,���v��|��czh�$"Sx��li8ET�	;W�f�nm�KV����.W�n�N�p�/B��y��&jRo�-rf����Q 5Ӎ/���{�'܍�K�zS��Ѩ%v�@�� Ex�˩TӦ������6���p�/d��QYh���Hx´�Ey[�����b�y.����Y)��o�s��<�b��� y�_^�ն��h�؝0���g��M��׳x��{�|Ś;
n�5��H,�v9�������4fV��K�w�xy�F0P��O�Z��t�k�T~�h�-�x�������m46��@׬�юJ��9JW��о��HL*����lj� a�x7��,'������L����qׯXG��]%� �.����mO��q�(
�f!��P��0��T�ے��g�"��(�#�b�'�*���+w�h�H)�Y��E���y�x"?��bp KF�z����l�������9��C�]�7;�5A��/�-�/�1�����4�{-z+q�B�?� 8J���6]�5�#�`]��N������_���*��]��>Z7
L���.�਒���
W��;�����B�C� �B��n�G�����g�gj�ô��^�GMaV��#Ym����L�~��?0O
e �?<<Q��l˂=s�?6����J� ��ݹ���*!7�"r���R9A�#;�α���w5Oj��e��V��)z7o.��JO��e�SS�䆗���W�b�]��9����f�F�?ŹR	Y$;B�a������]&�ϗj�D<ՠ��A}��(R����m������@�j:CŖl�>*�oI������n�Ϳ��A:���� �2x�#���SP�&���7U�$�A���,��4T������?Amta�سRHXj��t�ֺS�j�a�d���8�'TeQ�&~�>�;r������ζ7U��08W��k�[mm[��v'��Oœ�9(��f�*�0׵]�K��u����թЂ�}V·+�X����e�1j��L���1��Lf�}�����j��ѧ�����K�����7V�܍k`���hD��B�g�5fwr`6�����{rSO��a6+�B/���s��:+� 
B��?b�^�<Rn�|0���� b]�&�RL·ax,PA�L��լ7�&��"�ߜ/x�yMߜ+�� ���L��g�\q@~�>SJ�C�#'ئ�%@�(���q��XL��8UlV��'R�M�TAh��b�3~#ڤq��$����G�x��z�F� �]��K��S:o� �nR����� {7��W����<�����Zy�6�ZQ�RK�g>Q~��b��ߪ�1d��Ǭ|���8	��z�2���J�q�-.��Ws�{�>��[Y�����qӤ@T<Ю��+�}�vL(%ጎ#�i�Xjs���!����5� �?�
[�Έu�n��	t)����t�C�0�F��Iz�Ꝕ���5����L�{Mv���vb7&_+�K{aL��X�� t{�F�����;L�x`L`$t�Xm'��^O�7w�J���j�G\C��&j2�o�Y�����֑�҂�����}0��Jg���K<-��i�Y�7�����3)���Z�BÂU6Q�~����t��Zz^gHi�=M#80����8���xC�Ln��wCk���`)��#�,��f��8Vm�3��n��tt�((pؘ��ʨ�=��7�җLH
K�s�罜A-��G�}�[���5/�������xڋr�V/g#߱��8/�E|�ʮ\S�}�$*�����*��u�L����M��X�2���X�-]�jQfu<'kVe�Pl��Ty��uk�7�4i�q��=�z�L]���Zv�߮Pv��������)��={���]�\�no8ߟ���,圂s�.��{�ʶ�
�+ ��a[��Ǘ�Df���l�-|�/ty����"P�h��"ޠ_t����H�Q���쇁LM��~|%���'ZjN`rO���Z%�	�S��.�.�-VG�J�r痘��K�{�"��#BK?��Y���_����=e{^2xO%�|4o~�4f��QxS�F�⵾K4P���u�:��G�2/����[��Р!�����V���m"S���ċ��623�����hl+i[�"�h���G�c7��M&��FW8)Cw��/ﭶ<�QKDG�U�1GmHǱ��-�{+�U��̛Ȫ�u�[�a3y�2�R��	b�:Sx�k������C@������Vj$�V��@�a�9_/ N�$0ˉP�voǩk��@����4#�c��4��Ȳ�dyׄ�q�����˖��`�"J���W��DSz>j�C3zM�����:�ĩCE�%��N���d�@*@� ����I,�v��Rw���0.� �xX�d�^��iEB��zRAû_?�$J6�0[��3Y��S��dl� ��z���J�6������[%P0Q�6�cx3�<���$b;�җ�N٪�Hv�(��
�ֿ�[�T<>��c\�q⑯�|�l/���a�53����u>F���lx�%�eU�:Vd��#�F^RG��W�������(�J�.�������@nϦ���[���K:����<�HRK-�6>Սh���,p���;fW0�M���������({��C�ܥ���.�����1>Q����)f8�҂n��x�5�P�)M��o��Ƈ�ʈϒ��t.Ԝ�.3��C��O�p��&Lo9ҘbECj��y��ه����2�6z�Q�7c���ۀ�%5�,*һ��d��]+���8X��"vL�]'qՄTi�S�1>�|�@����Ul_p1�U1�ſ܋���ڇAUW�իT����B�[���Vsb�� �wB)--b�BG�"�l��EI�YD��ݕ��Ef��a$> 	bէ����ܟm**Xʷ�'�ý�	y�'~�j�&��# ��i{�2��*�P�cw�G;�r���_jQ�|�Z�3�Pv���K�U_rt.� U��V�osV~��9���;����`ɳTl��\
��dr(cY\�_e�IQG�nn��h�$0Eb���E�$�t�;x�?"e�}�iH��
�u����^��0��w��T/�o4�\2x?���;��S�O^]���E^l��@=����/5��~��У�_E�B���XQ_�n����R��N�������$�{r��Q�Vܷ��4$7��b��H�g�>���(L�ci`���w�~��AKl��u�.ɫ-�Ҿx�e.*�&;�f�z���� �)�o=�-i���㹆}�������/�d��P�w�21��@�J�kL��r�$��I�鷔9����B/����ϲA�薾��Ō�L)��+��1SN_�2��S��.>��|b���n���∥��uf����A����J���� ⓮�lE���H���v����l�>z���1М��@�E�������ͅ�z����@��eQ��I2i��I�#辈>����]�T��`Շ5��(�o����e�;	h�B�Cd��F������Vo�7�ak�B�QKww����:���{�[z��]�oN��zc�7�7Q2�u*�ƃ�|wmeԉ�H�"�+�ԧ�XS1�Τr���s)<k�p�	p����M�\�4����V��P�M����v�9JXt=5r��l.{�*%"cl9M$-�ͧi	|��������3���Q��)K�d��A���)�����I5g�E}KN����昴�F-ͻ��^�S�����q�4ѧ��ۛ�/�Ū�c�ݐ�#:��1`�uk�<�3�����8���5&Q��ǫ�&��x�	f�y�E]Ϧ$����/���t��-U�+�g�P!\����i-ơ��d���%�HN���UM�8Ȑ<�L�=���P~g;�P���;1�J�{4\T�.��Q�"����P[��m�H�'=Hn�WY~ˢEQ{Qd2qwv�R����J�N�,Z���]�S��'���4���'/.��/���ʀB�zK$����wa��I�`^�L��.
 T|�x	
OEe�����)�0�j1k�����֏���Xo���4�����d��A���Jͱ
�L?z}��_�]C'�p!��9��'x��`���T]Tuv�Y���u���j~}?�mb(�@KN�SA�?f3�H��>}�����	o�n#u�29V�Hw�,�/�{�<�[؋|/�>�Ν����҂q��s��Zi��W+\K>�,�;��+ \H,�[N�7 ��R+�leX g��ύ����'�;e�t8��)��au0X��5�:�y�c�v�?�8#�5����xI���*�p�/di���UwS|�A��G��9�2`Gρ�����;�P8`r,�-<�=3���͟�e���ƣ6pZ�~�����l�����v$� t���ճ9�������W����Z�$r����E"އ�ĉ����O^��8�Ӏ�Z���υ��<��St��,�������}B�8]q�[��
�G��ug��c�Q�"-��u�v�����RIS+�y����!1�i��-�.iu^䨞oZ[��]n���>���%�XQ��̱�͛�exTF�y�e�A����Ps���Iy~-pe����"�����x�M
I����B�v��v��]��k$���,k,�N����oW��glP� ��a���B��<�⯊]a��ø<f��r�*�� ��:N=V8�	+4L��<H�K�mO��U�؜�͋Շ5����!�n2�qq�>�e�:䚫(�#@+h��L��>��ΐ$�w�Sل�}�;&YE�������YO=��=6i>Ǝ��p]� c�cG���xw?%�����ؕ�3 l�uU�i��.���g��֎o��+�{#3�R"C�Z�#�'��,j�%�+�4�f�R��k���h�h��`��#���T,o�;yn�G�6����_�. ��`2QY�84`JY��\e�~��~��F�7�TW�.�L�W�(�����Z̞�$p�0��%?�����^��!u�3H����O\[[nN�<���?k���F\����9�����z����}rt�r��7�A�y�����Ak��r#�5:��k�Fh=ŕ��X�J��Dv���h�y�X�#��^�pIfG�Ӑl-'P�j̀�_�w�3�Sd�h�̈́��)����}���m�b(!ƪrS���`x��� ������>j��
�җ��"dt��$�c�pt#PQ��H~Q��́]�������܈Cz���\\z|'j���3�֡��ɡ,�ֺP�l�`��	iFz�!��T�I�FE�c��֓԰��'���(��(MmC�«�N1�7l��5�0�D󥭬#���
��=q�ň�Ե�g�c�ݱ�2owQ���zwaN�[�������4�����ȃ7����S�@�'1vX0�6c?�@i\a6`0�ڋ�e�fǚ(���R B�Tk�%uG�E�� /���30')�0u{��Ca�z
�Gh3���E����eu�F�i��@�%/�J�Qjd�f&V�?�IkuQ�U���/�w��G
��5u�/��3^��P3��4��L9�s�X��N��$����<5�Ci��֩�x�qM�ʎL�q�m����+K<�;��=d"B��������UN���;Oǳq&��	�2i2��!����!�Mǹ���C*��׷rx�� F�?4�7��;y`��M��Ϩ�w��6����Bg���e�:v�&���3tW}�--���,�e;ĂL���Y�Ms�D�*�dL6�) X�;�]吵���Kr41���M��r���B�5ץ�(���L�r��5�\����*�.i��"K�1�]M�����p�*�3|XP���B�?1g����Mb���P���)M
r&�~�*g�'z�9�U������&G�-�IN�S�"�;�\X��z"��܄��+\�.
�G��v�9���ҷ�K-)��7��Me�Lz's���:��wJ^R�Z^�R#GC�X4^��|>���+��)nѡ�3"����2q�*rZ��/ã&Zτ��7���@��jP�u>��j�P�����{��Zׁ'�:�mZ9�8�I4NG] ��m�C��� �S_J�����������O�<�|'�uޯ/��G�w�Y����,� ��8ݲ��FKꔄ���G�@�$�Y�\����V(����7y��m��vr���#� n�S��p�i�*�=b�/���C�4��N�
��y��,�S{r/��)���?G�˲tKP�GO�h�3y��=$����'�=�Wv�g'F쯿C2��}.|��(L�Lf�)���RV�Zc�s���K�[����n�5�djn�YD��[��2o[ ����7���io�����X˞ g����z�m�M�dg���$�7���7�u(�6���$��/..K���,t��H�띣>�jGb�ě׎�����q���"K2G�3��Z�`�Ӕ�ЩBd���<+��u͹�J��RF�Ct�0y�`����s�V ,���/�b;
&]f����.�e�w�QS�?(�`�J�,�z^۳�j����9��ԧs����"��oD���C��}l'	'�#�Ð�`Ʌ��E*� �i����O���z�Z�� ?�Wx�]�N��lz���DTpi���}gv��"vl5���k�o*��q��T�y�w���j�0
WII�^�ǁ\i�W�cJ�O����?k;g��a^��9VRz��"a'u6�L��\�Ȉ��?�,�7E�dPb�N&���+���:�RzXݴ���co
�<	v���t��]��o&�{7�)�'eO��W�3�'����^�e�1"18��[����C$!��z�����y���:�SY�SYb�Ϥ
1�K�����CP��a��8��Ƅp�x��7�oaC�~�p�{�n�ٴ�ym�~�L����"�R�yFi���?"p��MB��\�"XR�Q^8k��Մ�S�83����ѩ/x���!2Z�ߋj!�-<�"����x{̼�]��S�l<ԉ�6��!�9Mo	��]�'�;rq�������䶮�����y����>���kb5s�xR�����4M�w)���"$�2iE�ҝR=�{5����t@�pD�Ɋ{"��ߢJ�ƌ���#c`��o4#@PxM("��N`�Ax6�(��ԥ�8:x�=��1 ͏�
�Si�R�nB�gjʉ\�͟�/�?��UΛo±�0	f��z��40B�i1w�]Q�~�~�<&9�8����!~"wXΦ75@�>�b}���IX)�ԍ��vA����B�ai�@��˴$X��y�E�1�:�yς^�cA�ڪ�H;�$�q�FCGߚn�լ���3 ����֩UhF<��{�m3��[��`����0��1ᬘ��*�!�N�I��9#p��_����<��������K;�o�ʣQ���^�&	�ސ
�/���*�-�� b�&�
��5�U�Ֆt]�z�R(�!��ů*���O��������50,�>V���M�����	{���ۤ���ƭ����s\
�OO�"�NrƩ"W�[�B����9��?N�'�p�M2gz�b�$�u
�{�jF\��t���HO쒾܍2��@Ĥ$`��?c�#ps�b��iEjZ��ͥ�DF J07>�K�N�nf�[<�F��O*��>?"^8k{cB2{�B��,h/I$>Ab�J�����ÝJ]z8Yӭ�aJW��_�
ČX��k�-V���"�чSK��>l����8-[��6}��$r83M4U�A��H��7��|�/�@�����'�#��"le�A�-�6����ձ�%�i�d�n]ƚo�\nۛl��B�R�z�j,��5�<}�X|�P8�Ӄ�u^4��إ�����������)z$�B:35uǟ��:��	t�̧eG#p�MZ�4�CL_X��&�xf�:����,��E�퇦1�8?�#�P̅[L�Q���*5�??��Ϫ�c��Q�!�M�x��eݞi{|2�r�蕟@6�>R�\��5�>x����՛�f}r~7]9���Q:�U����.��j]�f���kY,OJ*�D����� ��`���u-n�7c��g��Y��đ��2���M���?SU����D/��Q�c�\���W���h��9���$j��b>3V+1�v(�5%hD�o��l��c��43�ch=~��EuY�l�\n�6]�z^mą~I�����P��ӷ�5،]8���ߕb��ӫ�-�]���A�w�{�҆�
���ؿ�V57�7QYQ��M{<e��[v
�\C�k�����PO��'���D_޶"2�<��:$q�l�ox"�#N�ǹ��t��_�3D�4{�g���I�x���Zݾ5�mx/���l�=Ae����+\uƟ��^��E-���L�ͤ�E�3�/5/LT��ܝ۰K������lMs:Z��5#���HA�����'2B�q7�Q�mt���x�%�r֔RM����lp�I�[	�il��"�ɣ�iO���0�&���4�8.W�y���'����v3���,���C?m����b�����v���O0�U�ut�b��з�<r��Q��	����ӫh�N�6�(d.ފE�yz�Nc�v�?�;3}��u[�Z�o���Kb!��z��F?C��,?H���&��vR����MW4аV� ʚѵ��xqv������(��tvx�VP��9���`��8�WB!]��l�8D�;G;�Fk����W訜nc�>�֡�͹2}����K�?�td_��S�F�q��k��ȴkk����A�� O�4�r�T�q`U�+�%��fMb��2�ĝ'6���j6	���e�,��z��3oP-�#6F��6�Z=.������A��* �ê��N���/��yˢ芍s=oz�P\�A��I�I-�Z,*y\�a�'/{���Zn\�ǘ2��;~�55�s�2={R�:�.�G�����T}�`�dS�m�SL��O,tLp�f�t�*�J�8��8��*[�5���a�' �|e�Q�o�j�v���:K��V��9'�aØ�g����1^FDq�A�����n�n��Kd8~1�͜��-���2mܼĩ��[�6筩d�:�r��_�t�{��%@NrWm
��zV�J�4Pn3�+�;^h�z��&���M4�X�51�S܊/�ѼT�_[aZLx���v�-%�)7�$��g��ԇ	f��A���u֘`�^�Q��:��y�x���l�Ǽ��o��ܫ����T�H�B�2�?�N>�87�\9/%u�7L�GDq%9�0r�T۲2�	Qo�bFE �,�?�Ϫ��|
�1i����JY��wk�'kp����G���4�����.�WtK(��폍Ф�BX�s��,��LAD�$ψR]��.�`$���2��)K(l�u;]F�%��н�~�������@���r����(�If�f9�Y\�C�)
Ը�+��cY�s;��bI�0=I4�O�W� 绌��!#�׬���JɅ1���%�2�	���Hid��Fr=��""����a�6�;� ��Fm����cAU����ԟL���^���jh���r�#|�"�n�Eٌ��Vgz3Vx6�oR�-t�1�hV�Cш����=
U;�)a��z��iu����-�ӳ�Q�g��N٬�:��$�L5Ā--8�����oǯ]��Ϥ$��<�^�k=Tz	M-�_F����E���^��փ��-�麂8������M5��!Z�
�DJ�x��>�4��dL[9��t]�lO�I�Ӆ[}�m�����-0�@1Ɨ�5�fI��k�U���J���.N;�:1������ �c�9<k����T��أ|��L��$�?Q
:�A?:KB���ti��c�� c�Nv�J�T�wK� ����?�R`��P����G��ݱ:���<)I�GugAB`+BA�h	(��:d/�Zs����W�	�nW����2�Q����uA��vw�Կm��k��z6���b<�|��v��-\�|�a��? �Lb�n��`�J؅F���K�(�_G(�R��b�5���i�^7��q�c��Xz�M|���u3a̜Z,�է��P	݃�z1��-z�^�ƙK�.���P6�c�b��X�vx�7� �n�
����>���ߴ6�����za�����Dj�3�34U�&R�5\��?���Z����� ƴ���866iI�P#�(T������{�a�1J��3r�Y��Q���њz>��G?+�V�$%=�SK����Ȃ<xgdm��e�7jح��G`$*��l���mZ&)&�����L��*�$�g��ru0&ϒǷf�m�v��=r�95.mI�9������Jr'�@�j6Xn���k{���Uv�Z����ّ@��@%�P�S��LʪC�ى#���:�^4H�p�W����ª��_<g�/%D9t��h��<v����'��W!��l�~���:��H"�R�x�%4������_����b׊e[s���x�~L����h�/%�pU�ۈ��g�5���ά�e�DA<�7+@d����3�w��
ϓ��#
M�B� 8�����(�ClaKT*T�����b������u�o���_f�F���	(No�}%o��Գ�IM�4)�{ѯ��f-���e0�Z�ζ� $H�>s��g��&|c.����3nU���oORU#���P^4���8Xs�L����hȭ.�ȮQ�ړ��c~%�Q< J�����z�X�CE��kP��! ô����1�i����SI5��8EIoo�Ȱ�q*U��bk��8?]m|&��n���>�M�?h�V���ܾ�I��EnԞk؋���ő�Y l<�ޫ��v@�4�D�氌�ʺ즺vb�rł������檰�������Ԍ ��v�ϡ�����E.4���)�i�F+���[��7]�$�-���^���w����B��пN�T���@����(GQ�]�s�����>�g%"9xI���*#][��|����Z���}$�J���V.��� �z�s�J��<����{�H�è�;)Jm�����'�q�w·T�67���h2E���[e��S�`7�ƽ�j7{gI� P<��D���Q\����S�H�7$Ŧz�1�8�{iջ�O(@2��չ�B����}� ���7�O�1XN黑`��L��GO�L�me]�.���q{Hdg+����ܺ��L���y��W#�Fћ���C��%uuXN�x��eL���Ke�Ĺ��_�2iB�1g�)���Ei�x�H>��!����a���p *�m򰎁��.O)��j�Xb�G�����J�{�R���;�H���i��5_I�Ԏ)ySs�?�c�QpuF���� �"�hS��/Yr7�ѹ�k:�M�C0����:;Ixt�"��ӫ�)�&N�0>7?$ a��u��7�k��"!*m+��O=Ģ!s�bC��ۼ�7SA�&~B�Ǻ�\�;�����f�9��z�8��0)����D����#0�x��X}W�hL�Q�4Y��@�@����1O�L$�i�>?s ��� �ɕ���{��OT0i��W�
C͉T6�m��y�4	P�D�PU?Ꝍ��uU�.(�{��K[�!�A�o��wU	�s.-J�L; ��h��|�;�y�7]��X�o02t�~� 9����!3�1��ى�O�!-�rÌ.�YG����._��r8TJ�C������?\ֈ%�UqKh�o�g�����ՠ�B�~a&7�n���u����Ke��YA�/AS �n��l����h�`n�Ůx텿SDoS2��N���aҷ�}E�Vw�ȿ��H.8�.*�Wa�F���s�'R�����\y�L�a�����#����/_~�c�g��̞�u'ӝ�9a�wL�$ ]b.\�H b�7��򄬹lS4�|@ؑt7W~I`��	G?�g�퇢�Y�~져��1ʣ�Z*�w���u%��Ծb��UB[6��)8<;��-��J`�3��X���%{e�:K[�m�F}��<ʝ����I۝'i+����.����Q���ƴ#y43�t-)��[���ʿ��H�E(PH2-�I*o@GU8t��U��;(���r���L*C���`��ZsZF�)]�ؚ�FEJIe�/L	�]��Q���D�_\�׹�б��l�{��OVA�8����=k6K0T����i5O1�~d��6o�gN=��P��C�0�[:�0���e�D�SW*)V���
|K��kwu˳|�C���}e��3u�����Θ!�&}i��,����{��@��S��0�Hj�Q�f��n�@5�{æ�럦Y�{Z� 1�B�cOC�x�ͨ_��&�m7�w�$�6�ݫZ����<�͘��L����&h����yB�����·�����F��y������?5gA�x|�%;���3w�`b�ې�5�~^��DW�|0���Z������Ȳ�-��UIz�*-�	~�@�P�=��K2Ȑa�կx)ًPܶ�<�+��7*��F��}X��O�n�_�ůڅ��km7�)�c=�%t��q���F(�?�:��c:����m�a�m�@�N�%ز$$�2�s��25�5�,))07,�0��6Y��I���:���iD����,���Ҫ�<� ��S"�>�?��Q�
5.(lDoF����2ޅ�+yMW:+�S�P�WqK!6�� �!��e@�ӄ��w0�:�H�~�褡)l���"�_���a��ybU�<�^<]D�k�(Q���h SR�(�$h��|�<�ڍM���a�Ǵ݈��7e�Q�=������_"|0����CV8�H�d=���C�����A��cm�9F?G��G�5��r���y�9�/E�|�ژ����.<�4F���Z}!MBNJYl��ӜM˴��<N|�=�]����� p��c��\K�]$Q6~�����O�m�štһ��z��ۂC�a[D���At�K����R�f��70#����Aq42:N��ړ�Df�Z	�b�$wi�**���d�B���4sO�L^(�T�b�	�|��;�:/����j�U�;��Ev��o$�p%����Ge�c��ɐ;�}F'h�w��,��p�G	q�٩�O��r�kK�����^���z/7�躙X6��E-�tY�6!-�J=]�D�o�{8���T6�a�(G��w�7g���� TPa�q{����+��Pb$��Wzua�*jB���6�P?���^��@�	��K�{z��M��v*�+-�<�F�S���c����߾0j�F����8N�u��5����{nHG��W�W �����X �h�U3���?��;�lĬ��4�B
X�m2*x����O[	�� ?�2��r�n�s�p. �O�؃� ����/�򅅜�9t��"j���K������q��G�_����<ap�j"�
~����X���'� \�-=�l��}`�U'�u�t3 � �u [L1�Тϖg�B�w���f�{,�s*��m�j%3�-F�U��nt���k%��兣T1�U��I���d�t�p:x� �kh�m%r���\�z\��J��
eU,������dPa�9�Pg����~A�Agmwc�������a�ؔm+.O,�'���B-�c��hR)�aZ��;�j&)Ϯ]!�,��z�T�{�������0f���a�m�pg�I&��/�~u;׆���=N�4�d.��yR���r��w]�����;��Z�w�����8����E�_�������D���+)=-l��(�嘙�f�0�������rn!BS���"G&�λ��k(�%���GB�aݞmpf/_�'̜�3��i�%,�M� ٚ`�E�p)�DP(�^�����K:�g�Ppg�13�]R��?�n ��NU��\Hf+c�SrD�1`vT�=�����5|+@ׯ�u�s��s��� ��7���0 dꢹ�I~-�ĳl�,�2J]��u�����	�Äm�>��f�rᣢ��fP��dR�cj׻R�@�zAv\rTЙ����D�����l��,���)�́����B1�1ҵ[�.(mE��)M�X�v4-�� #o���$��s�Ĉ9��TF
��:�^�at�%S+�E��c��d*��<���.��M{1�Cz�N�p�"t\x����S5/��%�$_�c&����s��V���mYX�
��;/�*"k��̗����%�-�w��tx�
�TJ�7��[)��*eԯt�׼y�Jd�2d����)JM�Ja�*ŨB���:���f|�zõ�nJ�+�<x�Oc��}�8�ɋ���F�*�kY{ϙn�6����<�2:���l�]18fS�,�1�<�Q��Y�����'2*#>�UW67حc'�m��kB�Oz�HQ�+mJ}��e��D�%�e�|���Ǉn
<�v�aڰ�]'N<u��m�U�(4��]"c���%Y�Nґ��R�L\p�CVZ=/��
VJ��	����%���'m��0mDo�?�0'��E�?�[��m�����
,ƩN�x�?�M	��BH���eF��3�J������X_:
fԇe\��5~;��A��Z�Y�e���v��W�T�V�"��մ�T���z�k�E^( ��?��PA�?�<ӑ��K�6F�K��oZ(�b�̕Q�G�0��?+�c�:f\��*��{G,fvi�/�&��#��Y��c�(����mׁV�����x����!�Zʆ����u9%��ۥ��k�8����r�s^oS�ş��k���RB��/NNm�"��^J*�zf���qW뜛8p�ADT%a�|����)ęǚ��+�5=�y=R� �Zjqu	����Y�u��j���;�N��꩸��gK��EI����[�P��"5PN�@Q2R�W�Vw Q�֣u�Iyf�\�Dk���sh~�JM��Y��v$D���	�R[��_�	�8���B�]7��;�V�=���˚ú��i@.�8@�|�{�g��99���-�\-+T�RM�M�|��^�ų\�C��Q�+�W�Ӡ�j�M��Cbf�.T��t�¼��/��<?��8�5M����n���kf�_����_W`��\�S��#x�`WO7�c�,�O�ĭ���5�?09��TYe�
P��M��_R	�.������n�1dX��-�'������Y�Z6��9�3j�TyK�Շ�gc�� Y�qJY�!�4r�홃Z�G�������Nwp�8��f�#��V�"}K�l�b|fS�s�-���r|�V_m�i���V�AX�_ ��.��?������}��q�6����aȠ��x��j	�/�A$[V�ZV�$Kؐ8���.���F���=l�D��ߢ#�{k��^�ai���y0��R5�ޏ�����9`aF?��fv��>�q�.���c�+�q]�@��2���X[�R�U ����L��;=��l�=�(���l�2A~�o���p���ݓo�j�Z�,����%��R�4}���,%eɬ�z�d���ޒ�̕П{�7�{wȸ�)9z���1'f�rc	��(������:O��
y�2���$\�� ����d��qø9=���.%*~��W��������q��HWR7[q*����Kg-!�8����Vq�1.yը���$^�?<����_���liw[e� ��Se1��ũ��P<�.�ho�\���]�0z�܇��\�0�ť�0����`���� ���a�p�ۗ@7��� 4�T�L��.ΐ��i�TWO#��J]f�k[!n���2�B?�ә�U�^]F���0��Q@	`��^��ik���"Ȅ�32��V`i�+���#���s�&����Q�]ƒ�|�f!
�g�J ��J.U5@t�Efy���9w�8$��@����U&zQe.���XC������o(� ������݂�Q (�����M�3���7~s1,}�e0�F��*ey����P��r�� X�f��6~�Wޭ&P$U�<Çe���)�rV�s>�m"j'*mnD�y���-J��Qb���6��4��#�9���x����1�Ƕ��[>rľ���/b=N� 	�|J$d��<A��%~ĩx�M�UG�P�*���o���H���S.�Ҏ��Q^t)
IhN� ó�*��v��R���l�F�6��+��a8V|x���]\%<)�1 �,o�`MÆ��˳`�0n� �I���caP�ԉm�A���;�%���l�;�FQ�U�x��8�.�/fg�M�m�n�+Qk���`�Z�@=p�B)��S�l&H\c�G�򅂬e~���J�`��d�� S�z�OE�w�8�����ZT�� �C��4/G�� ͳ<c@ /�+ 5<G�D�ⱳΓǹ��	t�/� ������Rxڑk)�`+������q��c�7�{\�7M��7��)↑	�������i�@�����R�ZI�6�����Y�S�V!��>�v_�d5+�h�2<M��[���?t�L��ƵEN��vm�qb�$r!�i /�M)���ig�*�b8��ذ	�5����B<Bd�@��'�*�7��������QC����J�x^�0db�*�_��t�̚�[�^qBln` Ҽ�Y����3�5x=��b+���V���z׍�.X��� ��'�N3�C&v-��SAڙ��3�ѩMuBOo\]�������ڜ�?��*����M��v3�_�+I���^�������|^}Q6G�=,���Ք9}�f��iQ���P������ `�ٓښ��8i��7b���"T�F��\d�j8+�0�����M���t�s7��
˧�b*�Q���\߈�d�w>K��f8��,�\\R���t/fv2ت�5Xa�H�/��m��E�A�� ��5�:Kc��G�+ �С��V�C.�=�����[(�&}1�C��_8�5���9�oF}|$s��<��GU��J=�}��D1_ޘ�U�;�/u��;�`u�C�5�8E25n�"L��Ak�a)��NK`���[$94N�v��V_.�����}��Y�2���� �P�z�=cP�.:��F���9HѧVJ�Z/d���_�������ߛ����7!�O�,-���M!��|h�s�|: �����|)�\+푳��X0���&�m�7�1�T�v����Hm���@q������XЪW���m�$��SJ�& q�$��O7턒�\n���\ �Pc�K0.��g!A��U%�X��� 9�x�T����x5P#�f���L^���ˈmk�.D����~N�sH���T�og�f��.k�sE�=r�IMC��Է2C���H������K�^�s��Ғ��o��ke���mN�����(���KWM6��|[�O�����?�������[�U��"�a�53��G���j���E�7�`v���
e���'����23qf���we����̊�:K��{
ȅ)��"9�mA�T�E+{��=ҕ-��֘�]��"�_�@܊��HS�&������a|N&\-�Eo3�b��ˈ۞���p�9ۜw��H9��xsFK�n5��|�/'��t��յWfv�p�Y;�����y.�5xy��n6a���0��L���+�<F�����j��ÕNB'07/��ݒ��̐�����C��c��%�JL���T�Lr�M�%���+���a�ӥ�VyB�![�<�1
��P�7Dxʔ��Mn�nհ=�"c1��j��Wz-�����d�:㪓�K=��s1뎍�fO����� kQ���� �jU�Su���}��/�f�vPϢ��W	���=-'��-�zb��C������Ca�H¯dd�kn(��%������3c��B�ϔ,���	���ՠR�cQ�����Z�Z�.�!sbx�1t[��n��c[L6���P��m[*�I&����QRZ�Oe�.��Gq6�Ş�e� I�V\Q���9qg~:ꬑ��'���.8�hO[U���
:�K�} cN�HD�
��ۚ���-�Wd��}1I"�	�k|��"JO�Ae��G�Ʃ�s �����Qx�S�E(W����T4Z2���kQ��>��+cv14�;$��Z=}�0�ܑ���v�+;����i�<f�#�y�:��l��U,ٖ�_�ؗ������WV�i��8KN�O��eW�{_3Me��7d��'���1�� P��T�\�i�����0Th@@2���7���b��tK��0��lѻfCM3�.2:�P@���rI���:sy(_�_X��[��j$�L�! Q�`J��]�;�� c�E�T	����[�|K��E��Y��Q�BUԉ���]o�&7=�F3e)~��� �'��n	.��^�AP5�:�H��� c�_�mF,$h���^1��-�K���s~k��{i6� ��A�S`vZ�����ē��c�����N�ٟ�.���ӊ?��`�iC��U����whm�P�~㤁X(��ƛXs�]���a�����%e�*!����#��q6��}���P�nY��`4�9�{j٪�f��/b��q�$��@>����O��Nz�ƱUW\o��r�+Cr�x�8"�k)ɿ�Д��I�~(��k�QdiT�e(o�)h�Xޢ,ϐi}�1��N���y�o����kn���4~Y��x� �W=���"y�8>L�	b4yԞ�ܾ�G?��N���_^��k�n�X�������P{�Q�ޡ|N�%J��f���Ԟ��P��3!Wz8\fF���u�e�?>����v�[ͅL�"s�������B����-aq��M�'�񍅊�G�����n�Rg�K���?���c�9��o�gB���|9�9��MQG��6�b�*��!���!��n��e�����]=JY�K�Fժ���4�.����\i�J�}���
X���x#Ly�^�&VĜy�G�m Q�2� �"�Y[:��֢�b7����&(��=ը�ʫM;Y�vW����Q?������oE���+ nRܬY�,�M}QXx���P�ll(�Z^_]!��x�*dq����S��y��	���3��/������������k[�>6Z"���D��7��
��Ω8�m�S:��5�"Vk���=�N�N�B�V�"�Hya�3��)�<Y�HH�oIi�z�P
D�톖b_l6��o2��'wp� 5���љ���GU|���%���+Lu=+�W˸{sfʮ�>�'�*_`�7ݴu.Ʃ��=�[��Q�f��u)<���	'�T$~r��]M���9Cd��u:�̦���i��HU�9� �{��R�勰%	��ʪUX`�f�/.�u�@���n���)�qV����`�=r��4����]��U��zP�Y5�X{{xp zR��B�#�E�ge�.�9����ǯ����y���2��OL�/K�8 �k^���Y�SK�]����~V5IvpՓ�b0�^Gsn������-�5>%G�ra������x�oz�.�����5�4�ЃP����B����+�hF��uj+�04~�3F9\��W�����4�q�$��#87U�<clزi)U�ŝ2�7��u��I+8p}�`�N{�����v���[��Cg��9��7Y�&�'qX���HJC-�xP�l�5(�m�S�	�s�d����'��^Nk�NW30jj
�B4܍۠w-�CVmu�����F���#"�d 7p��l<w8m��v7W���,�e3plZDóY�K��ʬ,�#���,���'��^(���(5l�z��_ڽ�6\�W�7���pV+���c����R:�+ň�ʾ'��EDe:4������M�]�<���3���8SR�dbl�<��G�ԛt�kT�b��
�Φ=>6�l��t
L�W�X�pV�9���c���Ƴ$p����K%���ܷ7[�8��.��z�)�o��U΍N��h����\kБ��M�����c@5s�}n�u�sF�jX���ؚ#k4�X��{H��Tb��:FC@Y��!q�)���I�O��$�8=&�d�x�;`xZ����Hf;���k��u�O=>o��X�t�[�ٷ�k\v��tW�삥�&)��������<�^��R �
���N�i@�h!�`���x�T&_�HBlD��8��\�Ti�6~)�+��^�q=}�V|�_bf2;Q}J:D�]�]aP&�����'��E��6��������5ب����Gm��0���?�5����:�Su��m�y�?� ��#�3�M�B������U��\v[�P�����ۄ.��|��Ĳ%��Ӿ@�=kիF�p��R�x��n6߼��`ꓬP#�63�9����Q& �_�㓔7����̵j{)����}���;���B�mIm�n]��R����/#D��m���d+��>Pkyl��ǉ����P�>6
��Dq�Y�8�0O�/�4R���rػ��}�E��Xؕ�6>є`]SL&1nf���iO䥖��9�	pB	%}�ex�XP���s����,�Y���W�ЫT�߁�σ����*��O�����������h�l�T�B2���aU��tD�t�yڂ�λ��1��&a0����0P����HA���Y��@���IB�L|�I��(��`�&u�b=�=�.d������[��_�r!����*���E����q79��;f�ܐ�Ͷ"�Y�t�y�t;lp ,D^�{�l��7��gPͳg��p(���J�R��D�@k��<zml��W�=���BV����h^�~��+Qu־�F�	��$h�����Vo�<�w���M�Q=����nj̿�o�f����[��l�x���!AQV"!b��=����rԊ��Ҧ�w����;^=�ǆ�z6р�^RD1�z~������oLX�b�:�R�΅$n�Üc�	���q��CkH�<2�~ʈ��j�oN��)���=��J& �<�"K��D�;0^h����,�5H<Ɗ����EJ���8%��}�A84A�{�(SW��F)Lk&�?F߁D�/�.����:+6�@�R�;��>=P��_�P�r�Cѽ�O��@� �·��0t�pi�Qg��K������]Ȱ�G�������!�G�zQa��g
�+dw���-_#.e����:����I �$^��FnW�����~?ϼN�	�=�6=�_!m�E%yel܋L�e*F��|�O W��h��%ih��gy5'����~��3��t7�߭K9Ji>']����2�w>�U0Ȝ�1Yr�7��'#gE?���6�*V5M��5�$m�z��U�*�x���s���$F����#��D��}�w*��@��⾄���F7q��)]�Yz�H�$�>w�[�YT�y�-<�$�}�E-���D/&	�
��ָ��Ǣ�-����V���4�t Er�c�N�&u�<g�]�d#��$�!�/-҉�M}��h�d�K��$]��+��[0���Py�[���u-(�	�D6ٺ獀����w,�� �"T��Ɨc�/@�[}R2e�
�|�g�����>��ܽ�.�E4\v� �}�r��tƅ%�C�IM,d�e��Y������6.d< �YP�OI ����c�T�a*9�H�j�!яM��z��hͦ�oM�͚�7�j�2���6�VI~�tD4�j|b�c�GO��nwo���z�s�P���ӎFM���_Gо�Bh�v�j$�^����*�j�0��G��ӈ	]���?���bC֠@fl/�:J��7I���?�Z4�Ax�3,#�^h��ja��� /I0�'4/2�h%��3:�Q͡�H\|D��%Щ�Qf����i@�l����X��3CM|���iK��M���bT��}�@�B�5�&+�7!�S��� ����L%�W�:� ��}��b����8249������U�%L~���������d�F4����|p{XƵ/F��i�����\A���Ow�7�S�Ot�	5�a��k�����u�H���͎�ΆhWzz@�&)�c��Y����uL.uw��z0�~`L�'��h����Կ��g��@S*�$�b��B؀��׊p�)o���0���<�K
����v~(Z�x,�l�-�UY�#z*GJ�&��WD�	N���Ҏx�e	G��^���@r�8�*I8���WZW�\6��b8�K^>QjYu��.�h�-�i7�ݺ:�8Dǀx�j��Q�}"bP;Q��~f�3�EQ�C�����6�(�}o0���*|��+Z���xcz��פA|��{��]�./�=�J�%���^O
�/J=�9!�`h���SᲞ�BĚ���٥kB�?Ҧ��� ��Om!�1co�~�q���zt�m��D����0���k�)+�^��?���IJ�x�����u����-��J�H�7�K�C���\�J�4��^J�6�Og���6�D->����4(	�<�������z�w�1�C�~�_�R��m�Q��<@��U�|�H^�*R�����K��jj �G���o0%*�0(j�������-��[+���EtI��G�8ژ�HTur�]���Q2��t=%���&h�J
��m�+I�o%~N�^"�P�H7"�������
ۙ.�uq��:+�8����g����x?�o*M\�&x3:xā������]B�M�4�<2�9��5y*{����ȶ�x�_�pv Њrų% h���]`��1�N�Mm����8�|)�u	�8��"yx�-�ZM�j�(�d*��wSJA!ܯ�
�qފ��%���}�D�X�'��w�Mh�V��[�-��g��$��j�D5y��~\�~gr�1b}k�V�������P�a�D��Z���YY�3�k���Z�F[r�Q�HQ������ElCT:���s��%�JK���W��p�c��}B�O4��"ؼ��~�޳�G��x��A/+OA/w�`�*ED��z����O;�Zg��R�dIu�h�JY�聆�$����dX�Sp`�K~'���Q�F`�ѕ��P3��Y�Cv��P(x�6�թ�}�֗����Y�= ;#T�Ƨ��(�W�Wm�8�&�ݣ�1�,�ޙ�qe��=9"R�;(��2�~����t˨�&���uL��&q��V�vD���0"VnysiUzI����=s���s�'ʡ�R#)�b�n0ݔ���X���e��̘�	�o������@��i�ro3ʘ$�q9-i�0��d��}m�	���;$ҍ�;�B�迦pq��(�X�5{.����6�%M}�6I�Q��ǰ�d�O���5#�#��b��D1���p�����~;p��̷^����(��%�a����=���Y^k�b��J�z(?�ـ�1�لG������^{�o�)+��]јi�l_�k���Z� �n�Z�*��'�r�%�7���Bt-��3�1����Y�{(����wCɁ�f�1�5D[��_e�%(x|�pc�FT��ead3DCT��Z�젦~�YSI@��ǁ%���q�M|�+��S	%�*�o`�IˈK�J��7�vOܿRrW/��Eg^�4��1sG�KY.@ˠ���j#�&l��Cp��Á��{󰼉/��A��Ӧ>��0�{������9{h6���ۇ�h^L%�Pt���Xja��x�d���R���)��ʑ��ΝvA֝������Z��2Xx9�/_�i����#��h��{3���բĚŴ;���_H�y�K�lx��0n���G�C;M,�/'c:_B=��o��aʎx���p�"_��M<�~B��ƞ2+[ƹ
:���埪�����X�)��y�'X0��:�x3>$�{��� �m��>�����߀�゙�ieȻ�]d(�\�� �YI)�70(;g�xA�ޕ�Ck�����t��`��f4)�#�����I�3�͚�z~nڏv��GSB<Y�˿�E�*0�P�)o[U�>u��,X$�j�s�7�ս��z�cKK���gG҅��hpfEb�A������%�E{+~���H�[�
F�S�o-�v%Ӂ������Uq��g]�+��3J>5ѩ�7ǪM$\X��#�ә�7�2��~j�����:ǫ��6<�1yB�%�����%���ɓ���-��#72��7c����$�>�c��!bMڽ3�4�e*��΀U�ҷ��˹��}�����#�������'�� ���0C��]9ߑD�>�v�r�^[��W�$6�SZa���Nrb�~��U���ݢ@f )��D���=� @WP%�E��ƿz��9��������i��'L��t�>P��T����ilE�)热��=�/Mi��h�[���* �d�h?�)H{l4��g
�c�zDp����ZU���s.�T�s4�X�C��ZQ�WE�!\�d*����]/��*i�p��8�����:<P�=z6{m4x7�)�"N�J��V�~\	�W��\l�^z_wXݖ�߅ʻl��˺�Ta�� ��/U�\_�~F�xXd�G)��sFDV��h�!����U���nv:��B�>������S=I�zF��)#�vH�7sU��m��R�p���ǚ�Y �]�~�x���,i֐��=s&�[f��#��8�ůӆ�I71�?x�����ۨ4NJ}�iDzqD,s�����!����L�H��ͽ�KD���򂾴�e&dH�>�4x ,1h��?TC������qg(������m����<"����op��
�Ǿ�N}�7�͐VF�߼�r��)�j���:�^�N�� �,�2�&�B��~,�`�'2~�g�#�6ns�+BL�Vc0��g徇���1�^0R4�(G���\%�(��aH�]�Bq/�`Hݛ�.d��{������{�s[�n���G���q���SG^�3e�M5k2��[܇��iP�@�̙a_�\�Wv�-�{��ըO��
��*ǽ�"y�h_A�e8�0u�E�ٚ��p5���X�JIdl3��߇��u��a�T]cr��œQ$h��A3�X)w(��yE���1{G�4�a??y6�D[2T��S��֦��4���4�����-^&�lgP,��噸0>��H�c~s@�y�!b��X��+��gE����U�����芍�)t>��W~�p���XJy�u?��FEI�HC�:��j>\�k
��{r�V�'�jP5������*/�$yq:��E#TR��*IN��2�Pv"D�!�6� �wz��U��h��Cv����6s��e,�W�N-�zt>��]SpM��6�P��:��q�*f6�ll��Cw�$�I�n�2��낱���$5�#�=��;*�Q0�u����2d��j-r�h��y�F�I�Z��(��Qz�UO���,VK"�^����EѠp������:!e�t7�6�<��g­�f'�zA]o�ϩ���S5�n:�q��"�K�=�c͗��Ts`�f6��ܨ�`#��y����(�5���-���l��0�5'Ǥ���$��8�0ְ�w��um��WY(���F$t臧jg��,��J��I��3W�a]Ebi�v����zf$2�s�0(��6:�?{�+s��	ON�z<&�i=���g'��nڤh�Ɓ��Ęv�\�\��	�;b��<��i�J[�>>��OCȬPoݪl��X��ux�6�{��h���`9�2�E]�P�+��(����)ʱt*�HV�8��~�K~/&��󏫲�h�D$y^IC�ͽiڇgHH�iʭ�jxU����'�8~���W����ܟ�Z ����aJ���(DV�v(�$2yEI׏˿}�|U[	Q���Q���V�S>�gn2���k�?����9�}o��I���������k��﹍7j�2����*�d\/�zG�=��zXDX�yi{��k�����b�S��q�2��Խ/�/�����c6�XMb��|��$�y_�m��a>�PV#������4��ۘ_�����@��[m�I0X���6�ȏ���T�,g�9�3{��1Gy���_;���9ȅ�� �����@~�z��B����`��v9)|b�׏5� ��wK�8x[d�mi }�ƍ���ŋ��$K!%g�d�.�{}�uΛJ��M���`��j!HK�=�$�x�6����ySu�#�c|p �X�H~q�4���31�u愥V�#�p�7oz���聰��\��b�ʤ�q��7)d�D��}����c?����I�h����_1�2����y��5��R���*$�<s���Kp[z��M$>�,�6yS1�Y?|�戜z^e0�t����E?�~��${���>_E\Mθk<��&��R��M���-# 7��"M�q������UU�_i� �2�������D���XW��gd�RJq%2E�����Rd_��ʑ�N/Go�E��v`Ν�L�Hz��Z*а�U��|D���r��pd�Ί�C�F���dx���\!��!�>ۺ��߄<V��j(�<�tB �D�Yh��]�E7	<"���/�c=e&8r�.�`��ġ���[
�jǶ�����d-��aisW��2&�S�ֿ�ݭLF��*.���$��S�e�[C����$�]�z?��q��e��<'��7�ԑ$�Ɵm+;W�%�I�{�}��Щ5���u0������	y䜛QJ--�&|Y��*ۧ�a�A�TZ��]D��Aq�kF.p�ڷ�����C�<-*��1 ��y�^��⦏��Y���v�ZH���X�=����3L���JPt
��C5D��_�a\��mP��F%�`���YO��_׳��^J �����E&wqR��8X@��ۀ��a~9� �7�D"�X؈�~�7�O����?kݿ�L�,ņ@�v���b��T!�+�S���W]G9�H��?æE����ZYx���J��N ��[6��4�TWC�łY?6c���ƉoB@�Z�N�Q��4�����c\ɤp�X;Bю������%s�A�)�E9zF�=h�3��N��$�%��GV���7���"C�m6k@u��$]8A2[�yџ�!�r..������W�.��hƍ*-��X�i\�i����
s���á�s]�5 5{̚�u�o�o���� �P����\�6�!=�$7j�4��}\�'���� %l����Nyng��SoၖňV��&ã�tQ���l-G�B��=ҿ�짃6%氼���{�*J՚�O��^b�&�ݓD��Dۇ�X�b��'�_o�ۅ��mO�-��3�u��GJ�ҟm��[����������tƠQ�{%*ŲZ��xr���	��˛��m��BPmC�8���p*)�*W��?���)ƦoJ�-��������a��/zq $sz`t�v���.F�����������7���UPQ��uH�'����Ю��N�ԏ��bx����t
"��e�!��������+'�C��p7KrD�9�0l�P\<���:�L�К�%n���D/��q��Ț�^f�Q�^�
D	�[̏i���<���+�������?�?'<���\Ź�+��s�����[��Q+����ʓG��Xؤ�K���˛��n� +a���r1��Zx���a�,�Y�8襉�b��e �T^�dHvWuE�+43#��OQ-��Ď�EC�l�V�d
��tO"̠ia{��C�	6?}t�������rG�+o�Y���"a����}�ĝ$��U��x���[C�"�g�-yƑ�� Z��[��s�PJv�2u��b;'��ȥ �v/ :o���Z�2q�'��L�U*�}�!��N�������orI����1���@+�x��n���� �`�˾�(�&B}�f���	�^r�g���E��Ŧ
J4K#�1����L�P8�L�b<|�[�z6֥"K#����ţ��q�w��WT�+M�E,3Կ���Ol|9�O
���Y*�H�0��ׄ@{��&��b��,����X�ӠV���E��d�tS�\�D���?�:�;"��1T��}�}]D���bKg��9N���Q�VM�e��`�Y�e\V͈�KJ�_s�k3˛7ľ�tQ�/�,�a����v�
yε�4�s�(�q�W��qa%
���RY;�����*(GdBk�OW�@',�ki��5��fDd��T����P�s�rʖ����f�������9>��cb)��э�=�]���mu��\c��\?�{j�#�.N�N�*�,�����ۖ�r�\q��X��cN��Y˗�vU�ԏ]��[�K
�M�����ʙo�{W:�����Y���늭\w ��.v�]��Lc�V� ���{}˳���a��R�f�L'�Y	b���#V��WN)"�8�^��&���U[�(���y��ms ����a�#; ^��!G�󾛿l�}�oi#�j ��߉���1n�A�2���ۮ�W�~BR��5l�|��>6�Gh�Ĥ"���4n�h�q/}��3t��aֈ�7�;4io�z��lö�b ��"|XW͞���S$% �� l�܃@�ƤY�j��
}����?v��Դ>�'�i�48L��RK���ŭu�o!�ᛷ�e�j���q�
������o��)���tҎ+c����K9`<#��֌`ԥ��yY\����zy@ؼm������'CYL���1�Yg��e���+u	#Ac���d x�����`���b)���	{�Q�޲�|x�e�/�`��[R�����P�X�Ŧe׮HƅZ:ݣ��^z��#��d]��V<$�}�Gd�t�Ԇѥ���U��iB6���%�gAU��F��xQ��P�W��e�pmJ}�As�V�M��_.$®R���#�R��f+��f�j��'��5ܸ���'�?�y?��BH G�T1���T��%B��ZW�^(����5kg>���G�~d�Kq��U�8IsU����if���^��?�'(�t��P��Ta,���7d`���T��Y��f}��JS���$1>�.��+�`���2	�D���@���Y��o��Zd�m6O��]�Hb:���4�ꌷ�S�H����h�@e�ϥ�=�!���aj�x��T�NG�V,�ǋg[�V�32���pp�%�6�,9�'��)_\a�h]�<�� ���s���b����z�z��-��P�:�,.M���c�����$o�꫼�"�TB&2'���x��Pqf��	�5n����n�?���c��Ȋ�t�j3�"'����?��۝t5�E�t�;�<��_Ch��>�kJ��b"��գO,-�!��"2���[�Vg�%�ak�1�(k/@n�~��$7�r���JdVxF�N�)׮.1F߮��7܂�tJ����:����L���T4�`��\,�h�` @�O謸��O�\�؂-׫O�߬�5���9�'%X�ݑƕ�
����ZG����=���G����l#L�L�d$�:)�h6�!3Pޡ*��.�\�m#�!ݗL+�y��#�T������%>�,"�JkU	j��#U�BaN���<\��BV��}>�ד�S�h<��a�����hSo I���^�`s�olMh��R���?@,Qz�NWͫ�V�R�j<AAGK����9��0�*% ����HI��D��H��W��P�� Kc�3��n#������"Y���8_��ޢ]9s����sՑ�[�My�@Q��e=li���(��i�X�������ž3~�~Z��A�K$��ק]��!�"-�$ѧ��^��[~j��:�B��j�<U�R{C,�����6Bk>�+f�!��B���R���O���5b@��;��%��Ey��y9�F�:�P`��H���@w�
S;��̿~Ph&-��w�(�ۃ�.X���{ǉW�a���$XL�۸2o
b��ĒWE��,�#NQ�x�g� ���dt�N����!���NeN���?W,V}@*ۑ�R���>�h��	��=FQ�=�D���3� �;l�{s�/7�f��y�����'�< ̛3�TR��u<�2ؓ�8����b�w�_XMc�H��*�	�c���ir9�>'��I���sem;y7��C����������B�M��ϛ�o'�"OR3A���7��MP7N�ӿݞ'��������U�3���m����^���ؽ�,t^�r-�[e݇��?"O��X'D�;Z\���	�����|��#��+�4�:�7+��Uѩ��|�}�_��K�c)93KR���=(ȫ@���0���eנ	����]��M}�A��wz%��F�nj�������Ֆ{�/�w]ʭs�ĥ��/��y�,=p��V����cgQ1׈峷�]�=����?��wvEE^�	*�x��~6��T�v��cI��9��W�t�D��)�р���K,��q�rυ&��W�n�㍏���^�h�%�pPpۆ�!*8�^�Hj���~]��6_r ��J�?�6�r=j�����NF�i�=��� ���&�ݓ�uR��V��9z�C�?NM�i�����K�����²�,z��m�pg2�iY�9��72fx��'
�(�p�p�iv;��SK!*9o`�"���ws9�:-��T���)uE�|��α�p��%}4�fwB1	���Hu+�<F]�_�ql�n�w�����Dݜm� =�c�������.Z�΂"��<��tע3�2m�Xa��7���!�:' vp'�暯[$����Z~�x�ʱ�R������/a�����-s0b�؍~�/2槸�b��״�����
R�oE�J8�>��"�2o}\�Y2J���D����N����7����#�q��_<�6�)lN�ZW�r_-@��BGo����c&�Ͷ�-��vt9s�~H��v,�#S�P+t�h��!�@-	h[��~p�ǰ���d�@A�!�=�l�r�9�*�9֢}T!�J��v�x�9�
�ms��������/�!0�f$����6�L,��7a�E���^{Ɔ��T��l���=L�P�/�ܢ-"�v�P�d�Y�?[�#�D��g�<[+���R�|�Y��P��Qw��W���
#������14��&����.���t�0�����1�������S��/�;�o�Jy���7�'�R59]�ь��Ʀ!���ş�:���K�6 D�tEhfb�%5������!�� �)3sbV��#j1O<�?�,�P��L���cf�8��P��>�(�9"�����DJ�7f�6R����QЇ��/Q�8U
�KnYrO��-�vC��R-`��g�޼	#�;��Y������El����������K��]m+F�6`��i�*)Be�R亸�(d��a�Z��(�#��|J�%!k�p�\�苿ޔV�=�#<�>�SZ�TB�D��Oh�-T[�>�gc�t�%��־����#����\��"S !�l�u�$VOg(,zX��D@~
��D����f���6���ڳ��Ա
V_@����Ȥqc�sK�:��m���&��� 	P8O��RxJKA�,T�������?aK�f�mo�%B9Md��h9Ϲ�8�p۲@K+��5dk:��]�Dc��Q�{���7��F����ۼ�'�-��*�:F%��
;Tiђ�%����T5;�ӽ��Rp��^�ߪ9NRew[�m+��>�ًB4���ϛae���A��s4����5��w��9ol3Z��@�$ٕ]�!�7C��[�-�v��:騃�ҽp����>���X|b�e��9� p��rs�w ��oiTB�i
�����-�h����ޘS�P�w3\}�|�!s�m���I�hY~t?C����������M��Wc��sOw�J<t��hwN#�>P��O�G��lo���a��tU���i����gߕ�'�M ���G�"tm��ze�T�:��0�W��^��I��1l�*^��(F�F�ƱN0P3��3�	��-���Q<�h��t�=�l�"�37�J;?DmS��_n ���O��E3_��׿'G��fՊ�H91ә��+�b�	(���y�^�k2�xֆ@W�B����
X�v�7���uһ�j ��T$�f��i�e7+�pz7N�z`>���6l�Z��p��@~�H�{��b��EL��$~
K��?�Q�pPH�b��w�W�(#��^��������{tM�XV�%�ԷR�J0Xq�r6�4\8�����A�qf(������_r������W�^�C��!j�+��� �V�"����vר��˱�=��a൹�[��c��U���gD#�Xb�`��թ/M�J4�}k��^�[OTt�+���/�:)�e�Q�����c�<j�]���n4��/y�����~�ي��ͅHps�:'��7 ^d��Xp0�n�7ޗ'��Y?I��\y�����'8�ٲ�u��UȌ�� �\�o�t\��%7������$X{!j �J��e2��#�����f] [yq#}cѣ�;o�xj�jt�PE-��F�鏺�Zv��BM_6%�[p���0	yt�L�p��X��p�[�; <ϪG�ϣȼ�������D��`]-����  �汵䐺rh9{��:8W&��#�]ݚ��f죀�۠x��q;I~-�`�P2X:�6L���i;�7��⧷�Hm|�b��9ׄ"#��H[�k�4�k�]����cj�#׫�l���Ⳬ$���C�>~Q�a@\nO_H��߬1 4��e�?�%B~�m���O��	�@}tӤ�����K:-e�lJ�W��.6�*M%u�=��ʾ�����D�Q+��{��6����$�i���dr�q%4��X@p�	�����*�n=�-l<c��6����*+W _���S������+����rbm�Z��j	i�0��J��<����*��x�3!z������(؉%\�s��)�mh�5x���S&�;�(,e�*M� p���Ao�	t�%¥�	ޒ���u���_��5f� ͱ��4;� 5%����x=���[��f�5����a&7�D���;5�u��i�p��2��R�6}u��F�[LHzKTx�Ẏj���m�����n�V����"��@�|�~�8��slԘ�[@�}�h��̍�������l�s����\)D�E4f�(�P��u�OY���ꏼ�0��=�t��6���e.xl2 ��d(4�g��NO�Z�]���
~en�o
38��H�͒�D�D+<\�A]�D1��6��h�9�Qb���Ѻvy�q]��"�f�K����\��0�!4#�,�o\�����2.� �.G���#,��u�Q��rg>j#��,�U�T��,�A8��k��ӳ"/�y�y�4Cg���{Dܨm�gI��űT��U^l�a�Z��gKmc�"&���t�qC��:aP wS��v [�
�9W���ssتR~�־q/͢�B)�Yi�{v!O}"�j����bpB����'_�d���y����hu�o����щc�R�j�o8���$=3#�A���Ux(���* )�g��W��~.����X��X����6'�����P���u�E�T�����
$��!��np��R��ˈ&�g�P"�.X+����ѿ�R�t��O��j%�+fVQ��`&�mo���m0��.d(�xe`6��
a�`�ͳNM.�
���E�SV��A���f{/������b���`�u����0�ץr�<edA����:R5jۆ�K#�~G(g/�����[�|� Fl\X�����S�p���6.�Q�e���#@���W�~��!�r�Y�Ҕ�H��k5��U[��#T�O���|ޡ��z�D�w�$� �V#q��~�(o�{4��Y$����Ё�eR�!IG7p&EՍ1fdU>'pi�b�A�r�4����ם�t��%�N����ʢ�2��� �����3����w��&����.y&3,=
�q�}�$�<�Wi��jҏ
�ϰp�ȅ�uw��	�^"��M��~9XON0��0�t��-��J������\���}4�1���c��ӯ{�R��䗐Q7=���k6���NA!��+���Xb,�z�V��Y��/8�洅�:i������/[�a%&���C �y��������� �soI���"ur��b�\��?�9��� ��2�J��!8��>o�j8�E�v/V�1�\s�
�u����6$�M",�
�>�����϶��x!l[��h2E���o�B�d}��O��1G�M+-Ba8���NP����%ǀ1|2�*F�8脿-������-�ܪ����J7�L��٤�۫�Ci��-e�o��JѢ�8c��
[�!�m�v�� ���{|u���C|̓��NT��bS�+��D6�:��
<Ϸ@�sV�*�Xv��Z��F��f_��E���УOT�Dnz����:�mu�� Zp_��A�܇��i�6��@~�]v.*f��f��|حG�
#�eE���b�)�)�U}�j�4�����,�H��ܠھj���ƙ�vshm|^X�c�l����N�>�[���TP�y6O,��zYr������Fe�n��)�F�t傾as�ݍ��l��c�͑�����m睺b����J�w喽r�&/���N��Mm�,�m�f�[�'���)��y6zT�;�"vU`���W`�ۀ��bs�2��"aH+�E{�2���-�ۢl<�̷��]qK�Q�X��'�ybR�-:CR� �KYȰ���وsV�E1�IDI:�����������ҝ|NI��_g�%��Y��l���R��Rҵ+	�eY�*!צ��HOH��l�0��?��J�'A�"� ��s��������z3O�DU�+7P�v�iB��P $)@�P���n�#��ً/[��ŕz%�¦0Li�b:��)�R� �kA����pDPu<66H��P���~
FV��[�b6A��ᶜ\>��9���W����}Q(#���}*�V.���ZF�kV��8�;;<]ݥ�GT^�}2�4�s 1����J����aȍ�p��ߐ.$�ߙ+��Ӂ1��)i��� )����:�����ῄ�hB�ʇo�v�Зt̓Jl7`���g��rԓ~K?���E ���U�&��%|I�*;G�����)�iif��CZ&�/F#3Z�_/���Ĉ��B8��;5���R���p��`�D��>d�z*�u����Ǣ���о�H�W~ D��=LD����;ճ����=�^ȝ
�*d7P,HJ�81z�H�g�k� �əF��+�P�)��5�攭���y4&�Y�a�),�9^�^�����hH6�2	��W0$6�R6��Mܑ��֧`�y��?���;��I��Y��	���U2�c����9����#+&9�#V��r�A��V��(���_�F@2!���5z(�HΏM�x���Oϵ��؅��7��0�S[/2��M!dy�z{/0�?s�Ȑ�фm��%a�x�
��R5+�ɂs�v6��h���)�~�E��V�����s.�$a|��D�5*����es�r8�6���-�!��p�<����*��p���/�I�bp���I� �DJ,pP�CR�G�w1����VZ�=�<i���H��n�^h�oicMH$z��`r�s��:yn)%��2����t��]k�[I	����P��l�0��S�!��pc��٭�T��,(US*l�ʕJ�6�RD9�Iw�A�%ř�W��7����#	�C%��x�heL�������7u�i����N�8���U�\(S'	��/s�)�9��������<7��a�������ڏ+�>��%��U� � �ݩ�M#�uv�D����b����d2/H�UT��z��� ���}��(�]��B_.HqQ�B#��pG4PbJ6�7'0 ����e1�bf�E�����~r}���e#�\�?��@�.Q���Zz9���"$>O��	�� ��אؽ������}�y�}n�+����S\��%e�F���+��1��FG�1�3������Nm|[dI.=�������#��m�r8���D��wG�ay�DY��n�{�k�wn�W��`�&�R�M�xm���]/O�2�{������3�d��PK���Y5�� �J�-�@��_̦6i)NQ�;Nh2O��w�5�[�]�����?{҆�/u>\��ۜ���{�(-���َ��4ﷴi��{ �����ļ��"N-���Lf �\����@�i"�L�l����f�+�,XGv�EFslL�З؛�y��k�]�8�V�drԺfEUۺx�%���i��f������^�v��|�����Z����2�eI�l���һ@C�@�w�K�}X�?�8�	��f*�l����4��#l�7E���}a�ۡB��a1˄=Q��_uM"��+��b����RM�N���NV_��>(�P��xN�^=�����(M:V9ڲf��Њ-�u:0 zT�P&�I��%1��s�����_�߁�âUU�
t�qe�*oi��h��Q~.E��{�����s��<��}�dB����/����N�nY��1\��k_����9y����.�L�%o�Svv�=�f�l1�G��q�v�ނd}Dpus͏?i�D|0m-��u�~�&Z3X�V�"�x�;�K-8�}���Z�������r�^���{[F;OŃ
8o�cC�����:�Vgz#��������A���;��Y�4
�ϰ�G�7	y�|\�0m\5���H�n�hk��{H���{�s�Й���Mػ��_t�1�0�^�̢=�Me�Z3@կܳ�!�bg���O�`�\�	�`��:mVnzTG�Y�NƉi0s]T~&1��&:�5.1Y�ѡ�cа�F�c9u�N6��h���,�f
�xM�p��Un�k�⍍3���2O�;������"��̣m����2NK$�}�|�:��� w�-�&�i�4�a`����.6��sB�vmE�� v+�5\ZE���ִb��$yGE�T��a��� m5P��^��T]W���/}��N�>T_����z���>I3��`v?A�͋�Ww��}��No08_��8=���?�%xxO�b�����]7άk��	��\�V�bx�9��*b�>FL�,��t;����Ty���*�{J�Zg���EӀ^�r��Y�Ww��u�A��Bu��2N�N_`�Sl��DA�`���"CT)b���\��@���㚏�Wp|�mr���]=�8��bo�k�� ��/~g꘲B��B�u�}tF}wGk��r_�Vc�f���3������4Δ>Z��v�����5�\PW� _4�|���QkJsL�E�����1ǃ�+��}�;֒�r�io+�\��W������L8����{�VJ�h5r��h��͎��c�D���&���O5P���$[�meQ�X6%E����<��^"ބKt��/,�۵[��E#��y1O�a?�i��^�'�K:w�@WUC�����Y�lJ`��n��DG�����ޟX���o��
ԓ-cw��{3Ł�ٍ Fı������V�$o�W`ȤdeI�����	F��C����f�E���&������0B^*��|f!#��x���Y;N&;�ˣ�´����ؖ�וX|t� �Q��K:v���, |��1k/�&�~�lO)�{ ��;�����`����4!<�!�=G��O���V���C��1�D�2:V!���Kʨ��	�6�<Aˋ�Jק��Ǵ���L�Ok[z���s:vRܘ����C�x4��Ξ����ݳ��05c��b��u�C *���n���y��`��	��>�>�:�����,2�o>�� c�%��e̦^v��9��D`���?TKR.�}z�^7���di����{	fl\w�%j�dp��9�G�r3[^V�),�:sY��<��]�£1OQq�A7̓�n5�F��Y,vŀ��P��N<6ﴗEE*\k�{���"Oax�a�-��B*����
I<��u��T�ȟ�йn~E�M;�#�q���=H�U�DUg��K���!�L�J�@T��1�e1��?��W(z2����CY�cpx2up�%�?�)��B�L�zv��	�od7�J���<�p��vwA>��Egj�H�j=z �����g�o=]��l�L� �af���-d~\���] 	fLQo�G�Y�����i�ԃ�L�M�	��<z�F����u�ipX��)�Y���9	y
/r�N��{NvX�̹��V��]K`�}F}�z�T��4c��9��J��J1�.J� ����r1��ML�`.zL3� ��y���k���b6q�4���X%d��K@B0œ���^���Xj�>�'p�f�x��Ϛ����\qd�_=��'"јj�<F�v�����i*��*e -#��{�'�6�ֹI	�C��ט�0~�O���g>���nj_�Ԗ\od:`�n���u*L�tЃ1*���\r,�����e���	{ٳ���$-�~��RY�:vb��ț�Wc�HCL��!���$"]�-v�]��9���*��_��h�r�ѿ��~�Wq_��gg<���ݷܰ�c	�N:�-�-Ⱦ`!��.�	�{�����=�Ò�ᧆV�T����"��[5[��2{	ɣX�h�o�|�.�&�����
�3):��SA���i�[ �@Fr��5ٿ�-1>5�c
��V�p�/BC���>��̶��-ƿU�����hI��C�X;J����bd5	H����}��Ev���_V@F�!h�50�s�=�Qdآ�h���qX�ԵN�,��f�/��6w��L�)��q;VK�Ȉ�vTN���ۼ�zsIx�kl$1<D��Us��1J�A��u��͘M�$�����˵�!C�MH٘쏁$�#��q^�(3���K��-�5/�F��X�����~�
=��)��4�l�5��5A�mE��w�I VR��M%��/V�t��m]�E'Ʃٟ���ޠ����2�v؈$�0[i��T'w��P����
O��Τ�qO��s]���6ǃ��.�n˾&�jy�3UM��&� 0۠痜+e=��CZb����A?�����@��9�#Ѣ$9�y,wo���y�B�!�/-J�4���j��Ɗ3z�sju\Pny�EL���@�X�}w�v_�Bv�MK�ބN�S7�N�?����N�\���� }��qj�:͓���_ZPO�YWC� 6f7�?���_p1�?���/�;,�E����h-^��j��,AU/��X9��y �E���A6�� 8�r.�'��u���Z�қE ��i8���uC������U���<��:�'�e�b~���.2;3�D���@�-�No�R=���\�K.)�2Q���F�hTrR�|~�kr
��*f�2��0
���K�<�m�&E:��k���ݎ�8�|&�껜:M���r���w�;%"��?��)�W�o��q� *M��Q��||�����)�lBs|rT:���U��!�;��P 7����ָ��M$E���rq�H�"=��A�����Ѱ��}u����ڷ���g���h=�#.�KwVK۰�' ���[�~���������D�ua[2���1�{I�g����ə*����d5��gAE���8���0�T
�'�zf�s����~���_/�ʷ3���@`��%�A�}L���w��"�IA��!�����j����Ȗ==O!�Z�$�7��pY�l��ܞF3�	i6mB�$C��<e���rC���%����v�"
�;�L�,^�w��Wbt�q�((k��zF(�Q1�m1��Ͷ�(>]/�}Þ��re־x|%�1IOi{+7�w�
j��	�-2�i�&��h5 ��]��z�U��q=�]Ci���,i���U(���
ò��2-`)�ׅPG�ߒ����?-n�F+��&v�s�!=`�c ��O���y��tF����/Y�.j����̃粟'=#$gX�fU���4A��}k:�&`ˎQ$̻���~�q�0�}8E�֋��� GL�!ΆO�瞓lS!�
C$t�5��)M��g[THl��?�V;q�rJ)��wU�܍��A�>x��V&Vt<f��Ŀ�\�&C>jw��d����!�<�l�F���>���]�Vi
�C��3�a�~��n�@��n	o��$�3#��vd֫%��#���'�Yn2Vc/��V���./���l���0�2��#=��Юf��4l;Lٸl��K���Ey�vo��&%�A$�֞x�e�%�
E�lLy�-��s[ �&�h��jHY,�f�1.�{��:a	`ݑ�K�6>zwd[M����B�H˛� �0ymO��͝��h_m�1r��W��e$����(?~�
X�B����ԍ�'��SqS�M+�G�\0��u����^��E��*N��s�y6�j1�1S�A؃�
�����6����y�f�:�LwZ�f�]�[ {�]`"|����S#d`��v���`n����M���4J��	x�PvlL��(n"��eX��o�������L̇��������s�M��Vד��Q����si+� ��w�	�&�J�ô���K�(1-H������#�Z2�T�s7��ỉ/Z���R��R(� ���Xhm=9�#���g&��d���&�}�e	CVJ�����?���2�7��M����a��@Sj����c> K����ę�h�xϨ�G��k�u�^d��>�i����O>�1��~h	�;O$oC���؛0L=4�
�Ae�ښa�V�|��K�7��.K�s��3���u=N��&�����4���Լ$h�h��hs�����VC��\�qz�����!6��;�8��g^��M)�0�'�hH��O�������7w�݆�\g��rB0����Iz�-��QP�����>ȍ��X49��fQ��}��=����G�k��eOpON�q�y�����7� F$�	K�I��nw���0G�qp�������eR���W�/^���ޢ�;���H���3F+7�TW^�+,Җ"A]��	��6h��Ā���N�C�t�+��E�]��Tjf�9-���	-����k�K�_zg�`��NP���׫��-/�{`23S
�w�t���)Mzw��b1v�����q��]�v�����W�\�V47��H�vƆsPɵ�����;��+-݀��y3I�	�<�$҈�z��
��(G�$�ҽ�F���D���S�F�Xx������N��jl�f�Rb��i��9)��Z����Wuϒny6��S�/������7�h+MQ[�;&Y̨�oVM����Ѱ�ѻVA��p��j��~��=���l���K�E��:W��&I:�h+�2�zf�����3���*m(�Փ�眅����_ңeM���H#���baq�!ux�a@�hPr����-�3Z{I�(��ie�`��	�+����C�Sa�%�m}·#o���,���G�Td�����8@��?�rVf�J�z�i�y��b���������)��h#���LHScQ�r�n�q���mTG&�D��p1�ՉA���,���$�����:b2&l���h�Շ�9.�M�{�}��#V���W�׬�~q��f �uM��P����8o/\�J�%��A��T�'��\�CB�)�P��W���q�Wd�GZ��jI9n~]�G�}�K�p暁�S�-�6�`��RJ׀���f�Ø9/*������',ơYd��z)ħ����۵FAԤ1d������z��&��h��rwic�?4!���%@��H��/��`�#�)l���b��!<�!�旰��L�Л��ڗ���5�$��\��X%�W�o�L�2H�.��I��\�q��X�I��&r&����->1����wg�Fh7H�*	��	��=�����X�f��]_F��wc.V�Z\,�	�Ԃ���P��OÜ�)¤�r�{�w�N�_��D�i1�B�N���U����E�V������W�g�$���Z���h	�8/|7�4ԥ���5p{��Έ�a�v5�p���� �?5q���7?��/�T~Vq�|COuΨ�(M�l�*jX�]B��K�1/D��TpHlu��k��<缅�����¸���|Ç�&/bU�	Y\h+K�f	�&��U�}k�ĵ�8~\~�jx<�X�j䐫�?�*��]��2[CށHR����<>�=�g�#���*h��!AZ�حG>�)�Lo�X,^��✾��>�`�p�i��H�ehC���*9�x�6ڠ����K�qO!_����q���k��/P�5�.�=�����|��8b�S��jl����LS=X���SX1�cG����;~�Ϊ��g�-���jnOv:BApxky	�&�ic�2���(�M��\����]Z֜���nO���c%�W�d�@EDD��r��aiMpE��>\3f(֪��P`t�c�E� �E�mS�3"}��,�G �dob2TL�4�C�B48�ʔ�����NAy0�W��'���i Z��^O(E�:uY��!@�R N������LT���yˆ+c3$�n�����b&�����h�8�.f#t�M{.7��'�I��l��̈��I�ߜ�ja�V��>��kEk��]�Y���&����-w��d��Y&,���f�e�dԔ�%���G��.���{���<���R�]����5���uo9#��ǩ)��b��pl+�N�v{�p��*v��w*��^=�	ۊAlG$tc��S�U����PT��}��=AC¾���h��YG���w04��B�,a\}��B�&�3�\]�&S�n�����4p�����	��{yU
�V�f�!� ç�8��U'�?�ۖh��,��J�����z!Ob��ٽ��a=�+	��s��=�*0a<�I�%Ӷ�9)`N0g�Wd�YE ^$�i$8�Rl#K����!����vv�|x/\`;CZ)��Ιb<}�<�4���r�n�È3h���d�腹�㤵7l6�J���/򈖴=E@P�T��B~p	g��5q���l�NA+(��Ԕ��ܐeEqnc(��mAS����ЗS��&��~�����\�mj���/�xh=ev�N��{��a��2�q0�\��z����B<�b�L��k;7�h4��'y�od�C�������n��S��=_J�5\T=|�����Z��CI
�éN�.}O3�D���G�[�cD4�S ����j�����ȀO�v\o;���Z����=��I!�z��)=����!��f�]g�q��y��L�h�ۇ���&K�6�Ug�t���)�k��9u�7�ΌYm�F�L�RA��g8/�����`{�>WP
}�=��L�+f���P`E����f�k���^&iFͱ2�v_jG��	YT��~���[FVx@�m3�A-2��H����)�.�I�K��1�-PL�܊�PTю��uH��\����x �����ِN��S��Z)D�J�3<~�I��Y�]c�]�}��}��΀aN��ViA��׺ˌ��q_�%:��*gs�*w�nؽ�xe:U]c'k�޲�����Ӽ?(\ͮ�����̹�¡@I魗��8+���O�:y�_�=�/�B����E֌"�Vc�U�(��7#�:ߣ�<M�)�c*a���˟a9j�p��))�mC�/�����[Ӵ��쮦�T��oS7 �"���|>����Q8=|�z7�}���a���Lz^w"�Hn���H0�>ÿ��6�\��SL�$
rFBat�|�r�n��������iz/��^]�.�����m*h��X�Ls�N������`���7��8��a�g���bf�:5܎2'�T/�?ѱ�=��b�2��V��)>��|w2浥>ɵCs2�f���x���H�=ylN�Q�N���<�%:��yH��܈'�c�
�o�t���|ȶ� ��ö,�Ϫ�Z�#��q�3�������i�%�(T w�ӏ�+�izW��ǎG���et��� ��w�ϫts�D�L���C�{U���^�T����Q��$%U�an�2��^(�g��,�S},��+��yC�Og?�u�=]0��/�I�C��R�
آ�9�;k7Dj�P�s��� NG&@ʾv4d��[W
/�bG��
����(D/�Z(R�|hQK�T�mCv���O��j����*��۳���@�WE�q3��i�@�_����G���c���O $D��+�^���T*b���#�R��{�5x*�$���f��q�p~>x����Y�ff6�ɸ�ߚ���TP���;x�=t��~.�{��2>���i����Bj{�b�{L�&L�OIOY��C���SS���Sx>]�q�	sr�g�!h�w�<���{,��7r�Ph"��.,��t
�JS��`�;�^p�Џ!o.�Ὼ['mY�v���~���]��W:<�2v��?�7Mi�n�1늒��ɑ��TG-@�����ѐ۽�y��Y4E�(�\�/�
L��G��WM.�LG4����韉����H�}1q��fl�f�
̚Y<�4��;��0hy����������Za2@�Կt��q��P
gs ��B������rI�M�i��C����J�Wo�9����y-�;U^r�R�����y���֋��7�18h����D�>��P���0���d�M�b��*��>~��?�$�e��-ת�u"WC7H�2b.�Gkg�sO`-)%�״���0�?���,g b}=P$�>B�$���a9��R݀�'�z���������T���7�����[�vcg%�T���ק�ͪ�ϐ������L�ٟ��cn-�ㅚ0���]܅��#�߲N{�|;oX���_���pw�K��5#3Q���
IH������J.����0>�)����6���;�j��o��[ll&�5�ax���qP�Wy%W�$�hO��G��)�6��bq-?Y�z>����=��U���*
�p�����o$u�n�w��&���ci�#���'�C�i"�Yl������f�2�5�z#�r'��r?t�q���\wX�p��B��KB�V$Ւ��z�S�NC�Y��H-4�T��/�����S
���ѭ�.�m
m�CkNKГTg�	;{�X�6��"��\�/���F�ԃ��t_$�LM����#��� 
���-a����#�F^�<'�T0�������)) ��}+�22Qެ���6k
R���O��t��h�w��aC�v�b� �c�zL�0wJM�|M2B�!�)#2|+ޣ��ŋ���|~\�۶ofm(pڀwu�[��^Z�q2|�6y9<�D�{\!�y}h�iD����v��_$�#[��`Yk��bn(��5۫�}$W�놼���x`dB�$tc=�$e
Y�K̀V�	7E�V,�&f��1H_P��*/\�f��TK�G	Q��
/*���7�a-�	��fHLL�t��o�"�I�����7/�>�oP@$���Ce9s<�+�W��i0ƹ��䴁��W���}yf��5!~p�=�`8���s�M�z6I^��뚵�4��H����׮����f��[y��=a��(�:p��h��`���k٥+�+޲��1�6��my?6��/����^�~�yl��Q�8,c�.;H+ȹ+��d����|vo�v�L_�t���i��(n)�G�6�V�6(T���M�C�lV�mܮ]��[�P�ym@7tҧѲͱq�߸����#N�'儝�W�'����c�9�|G֠Qb�vD|b����>Hj�e�tp�cK�-��
���xRt��hi�~/j���6C��`�I���M�e/���3���1/YO�C~�;�r�q��S:%�obќ��-t���Ғ��K�'�s�ҙ��
���5�+�)Aۤ��򷚫��2���s�N��.������m���z�=���1:�[8e�c�G;<�/|OA�X�Ծm5��=
r��rl| Y�ifo��F��������Hu�X<��]/Ҧ��}<�$Ўa1̿ֆ��}NC�����%�����_��O��iS�(���'~rIz�ߩ�������M�sZ#�uJ�2e�M��Ĵ�.F�	�8	�ׯB����3�ߤ�\fP��7���5��0��'� ��J�w'r�n�yz�����.�{�'U�m9Vx� �Q���(��E5���n=w���D"�Oh.t��r��>�(PJ������}�`'�+�&��1� �i��A'j%)7��E-���&yr���*��&�D��7JN������&Y0��Y�K���UA5�M�9�8A��������D��<�P�؅�p��Skw�mCV��T(
0?��9�DZQ{yg�(�;�x�r|y��+{e��&���|�{�����$+�1�Y�!P�7�d�Ia0��j�{��C�������RB]mJVZ�����g����\jٸ�ط:��HB�sv
r(5��!�+"`��E����il�}ɠZw�ޞ���͏��-:�t���C7��j�� ��vy�셲Q�u���i��,a��A������j.�G�D��'05;Cz��H8��@�2$�^�x��["�����GT;�� ���|2�'��A�@�[�_YMG2�(%�kꇒ}�?F�8�}߸r����b�9=ڴN˴���"D�eOX2|h%
�	g��@��N��i0<�͋�O���ȖX�]+��'7[z[�@�ɜ}5�9�g<ϙ�ea�/��xO�tB�,�9��E��BШ[�WX���E�v'�O�� ��ñ�l �Dj�� y���G��n�JR�;U����Pi��Y���-;��G��F����\�Y1�h`�F������رX�(+�C��"���k���)�ir;[9n@��Q~h���n����F5l�eK���mΞ'��Z��{�-`�r�+�� ����Es�`�l��˴~�F��~���Rs�m�	١n_��?�̅z��\��i\�H��������$P.8'��^���?�Itc	�6�����-�^,�7 ��T�G�%[�[6|a���]������ın�_�D�e�WA7�/��QW0�1�a��A�����r~�h(H'9� �^s�z��r����K���
@��:�ҬZ#M���nU��*ס���G�=gZ��N���#�٨�!:Q��,i����E��'���d� ��[V� l>�T�?�;� f x��G�V�S�9bʥ$*�A[��3��ą��A��[2�-"4ׇ��c�lq���ƀ�]5��U"�x��S�0��n~Hl.A�U�aެRt��I�
P�V�36�N�|��A�Fs�M5�}�f0��Ѽ�A�O���yŦ9
�����Ԛ�qH�m	�i���XC]o����D���!�ֶ��m�"�H>��.Ʉ���w,i2��ӝ\�HSu��E#�N5�O��U�P�Y��h	z�1��2b���
�2\PF96n�)�K�$�
�1Ez%m8_YOf_�錂�J���`|S˕�zZZD�φc�����7�Z/D�%�b�=}1���W[Čl'��P�����7�Q[%Jsh�9J��x��҆oV�*�k���i0�*u��gJ4������L���F��H�l��N�4|�� UG��]�M�#ظ�ؔ4\A�G��+��x%��_��+@���a"j���Ʀ>[�%]�'D���B$��e�{:@s�Y��F�:S�c���Ā�i-��!���y�甐?AAC�uPߘ�'�

F��vԩ�a��76��y��~�"C�O��Չ'�v)V�D��Q�R��ΰ��k�W��I��=,�AM�<���
6z<��Ŝ(o
��W�n~�%����{ݥE�sqӕ�2v�{�Գ��$�*N�;�
������H�C0R/TO�À
7e��I}<�`)p�{�`Z�	,/i�O[���Gr5�� n�w�A�J����,�2>�xRf��&�ƥ���_�2��Ո7\P�-[[U.�*p�v�-^%Ji�!/
_�:���%���i���"7�@��pɒꯐ���Ù��RWQ��� gX0s��"����WB��Sl���FWo)�m"_�}-S���y��HR����x��A�ɯp�'qy�o���/��i]�����z5p������-e���Ze���W�y��foV�0ߺ����W��H5�������v�߁J	$�9Z�L�)��V��6(��ݘ�!|;�O�K�=�ot�"S�$!!E���׊�+\��W�6ItC���a�-��A�y�0֤W�}T�]�!;�{�^Sp"��~@�!�ty�̇�@�S�����D�=!���z�ק:�� B�47��eJ����r��5�+uy~'QM�_v�)m���D�,u�7S:K ��I������:J�5TQ����w1I~�8�g�_�����(�;�U>k��u�P�ȝ�������hX���EǷb6�ʹ<e�T1��>$�a�Bʦ�R��7;`��6et�\��tbs�m�����rÏbB�z�+�� �˅�yH ��l|�[,�����֬:_
���������V���_,|��s�Ԑ�ǆ����_c+��3�n��p��|��`E���5qgkkv�޾%� U�
a�".�Ec�y�0h�ٕkg��A��Pgh�q ?��
Z���.�0=*�9�4�lt�#��)���SO1B��bl�c�{M��;��}��o�`I�p�����W�B'9%��,�����^�	�[h�u,�؇�*�0e|(�3�oa|�����Z6�� [��ך�ϸ<^�b��}vNNOz}P�]�>�F ��y>En�‘W���m^L���?��=C��
gM�`��9��m�e�ls�H�'*c�xǘ���},&��DCtL%�*;]�]�t(�d�rݺ����y���hR�z����t��E���DB�ΣI�'}���f9��_�jIaA�@����t�H�8���d�����l��e=�;��"�I3�n��Y�X>ўZ��O����BU�CN���'REQ���� ���{9xĈ0U8=82("t	�WFŲ=[i��]�R�`�i'��V�u&����?ڋhks�_yi�7	�*0�>A�h��a�9o0y���"�N��z�W\Se�������������x=�~��\&���2�~�{���!g�Ǆٱ�4m�L�O�Hc�d%��űq^\��'��#K�T&
�⎷�N[s~ D?�=�Q�pi��eD�Ns5A:�N�H�yZ��hL4S���Q�i���+���Ǫ�4�,LsYW#�w���۞�������
����M"�ô�9�����↑��urh{d�ο�]�g��&]$������Nc�z7.�^�j�&��dpc����he����9ǘ	�XCj�'�}ή���3�B S����-ꢨ�hbU��h�������I�9M�Qt�3W�H�@(��u`��$�����KU�ikC���$+ꨖ�\�4ca��(��P�-�����=��Q>8����NJG�h��a!|���e�l��8��E��=�]� iʈз�Gɧ/�&���Y$z,��L�i{�g�ز���e/���"([��6��"Y��s�`D�j���C!rp�N��`�	Ȍ{�Ͷ5�X%�Ue5?Fꚦ��C0���6u���@_����Ȃ��;���D�}ẕ�mNx�5"�Nʷ�/ϩȯ*d|��������nL���8�O�:�7m��s��Z�Z�LP��g��8��M�c��<P~Is�D���?D�����~��f��<�.x���I��)x��co�b����/�e�8X�m�O
�X��dΒ���fCLUĭ%9"0�v]����Y\0��}�c"�N������u�`]�ă�\� ���]��%SԚ�Uo��~%�ϵ���}�q��9<�2��Ur-��m �o;3�tc�2������Ƙ����yP��d����4�������@�膗|�2~Rzz�
�|���Sfr��f�W��RJ�N@.�������j�܊l�]:�u,)?��9��wP��;$����_�ѷ�a?�9�{4��\Hx��c�3~�̬u�s��Į����:�������ծ����������_G;��d�V2�{)�2ml�],��B[�ܽ<h��J�^�8�6A����l��3�:�e�������V!���g���e�[����R�Ӝ���3�q�U/ǀ�z|>K���Y���~(�T�Q���a�Gu�D8q.�1�Ã������UX��(�O�?!��)���*��A����U�����#&wY���	�9'�c+�X�/+�g��d bi� ���SA9�$��0l��h}3`x�y�V���!�qoW��/3ע�<�N�&�o�:�ab����P�v]�X����+�+��Ebg�9�銇Okn�!�}G��~��\�13�}�G�'��aX�W�0�H�����".���.h��$�bWPJ���NM��ع��U�MS��Z!F���}$"Ha�Q���-�7/&K��La`� ��\�D����j��F.%v�R<�>���C�r
(aR�2�`
�1�\)	*rƂ�`��#J*,�V]ip�IߕUG�*����L�+�1�ӹ�&��pc�u1�F�lX���t��՘=�9ԃ`8tx��I��ԍ�C4���ĸS��́�H$���9y�ne���w��=\Q��\��1�7n{���Q��8���_E�(�P-5E�4���;u���w[3�vj����9�N��}Q�7$�l�v�c�a���L�V��s�⬄dA9Mr}��L�:�bI��U�G'; ٙ&��(�ҋ���Q��}̬�nT��U��쫆�V��'b�?Z[�!�!]�gm�4�E��O�h��9&ҺØ9�����h1�L��s����~�&W�p���X���[�_nM>T_S�ۤ�����p˱U!6�=t�u[�0b�� �+t�eED����\�f���<���� ��S54N�+��.� �T��(z�5��e�evA�[^x���:�K�A(�w+��$,���r�>�'�t70��)SW�Ef�勘��� �&y�򣏌 ch�ܾ��&�GHD�#]_�#%ߟ�N�K�V����Y���1�S��k�D�u�d����'.�:(34�M�2h��*��Z!^qڌ[��Ě�Vt,����.����餷sO?���`$�G�?�и.z�%�c�)��?Q	s#O�!���j}A(s��^Fi��y���0�x
'��3�n�e
�����m�e^����5$w@*~�w~�Dlü��QJu��|��7�B[�6g��(��(�0ȼ7�z��ˬ�Wg���>Vi���㯒��5X�$�I�o;�벓�4��
k#0��I���K��^�ԁ/e�m���x�u���T  �:*����+X�/��^�e&�ͣ/�=;�u�`&Xy&�^�j���,Bv�޻Eߛ�axNyv=������/B�YO:7�t1?*��%f�����wVüYq�8\%������ٰ����B��P-ɥ׃���T��T����� Ljp}���O1��
������N\y����lV?��亾y�N��Bi�/A���-�	g��@�K4��Q@��^-[�8����'o���?t"D;�����B~����Ǖdr�v�\ʃ"�M�n!���DO�?�|&���j�<���W��GU�?1wc7*����y���A����Y#�-�z�0F�S�46ݍ��vZ�9�}l�>�kXL����L@JH�\�*q���31Ӧ�#��.�����ⲕJ�l�c�`\��xZR�kX�h��ª�rW�Y�3�R���j^��<���h���2q'�J�Ԃ
���ުh�'���o��,*.7���Dw�[u�Dˁ�KB���S���9�+悮�y����l�Y||�u���+")��>W�2����.J��v
|�e<NA{�s��H�7%a��_J�Ӛy-�d�;��,����s���v�%��`wS�{�lT�:f�=T=�,�#�����t�:�S��é}j�Vvɗ�`��$�����$�f%}91ݯ�J�$���̔�	f_)|�������tmM��rZ���xx8�_��$E�����q�/���,Y����7�A<�[l�V$�U��m~J �jHLn$����׽��U�,T٩�i2l�_|�)
�Pj}����F�0���(��/I/E�e;1�*ߣ�y���%�\v0o�6�&�g�*+۟����ᅉA�5JazV�dXFP䴵=&���%O��G��H2�-E��4�������>�j�d��e�	̤j�i73�E8#C��Q-����XR*9w�i��W�T/�A�@��L��B�Z���Fb�<�)�eIC_�D�U^�š���"d�v����!,�a�48&0��=1uu� W~Q[o����Ut#��}d�xz��P� ���dP�i���~��<�q�r�2e_�_�ӕ�e�<ٯ�y���8��.�^�4��3��ԻQ}�/���QK����h���y+��K�H�FvC�Z-|߫(�`N���ߗ7��֖�9��b?�>��������^.LNhr�0�<��6�.@Wl?�q�i��7�[�k5�Q��`	���Loq7H�����D�쫄�����h6罍.�r��x�w@4 �ծ�uv9��� P/���]���0|@�)L5�;�`$�Tm'��F��3�3_��NPˀ���({��p��'F�?�;���&}2hs�|�}S���^/��>��@�O-L�Hb��<�����x��	���8�� �/����/�Xהb��W�a�9�ui��}�,��O�[�U��hk!��d��=�Ѝ��!9h��� �s6��0��w���
NƼ�I�R>���F<%�ȼ���h����b6Q++�9 �毚�o�[*ߛ�?��*K�G��Q�����;����$��B�zm*l��7̔~E4��8S���Ux����PFD7%v;�Q��OKg���|��¢�
�I1"@43ok�g�����l����G�O���ΰ�h �ݙ�df�w�|6��K�f�2'�Ó���A�T�O&9;��ɚp�`�9g��^8	 磦�#�M������y��sCg�p���g�B�`\#��ߡ�pN"��jԠ�� l�k��|�����.�e��/h��qq+��d����v
|�?.0C
�~� '��q-:ٯ�	��LX6�����O*��g��O��l8�w#��� v�9���� TBg��g�m<#q��? (�`n����D��[���6E&����ZUQ�����5ضCɮoF_�\��,v�.�rO��Mf��ҋ��a�sۘhwϠ���{q�>tבּV�zr'y5?T 
�/$��6v= �[�����l�E�	y�p�=h��Bdb��N¾�)�a��fD�0�9bOXlF�T2WBT��}㰹���#����#N�����F��a3��$���׾�o�V�[�ܥ|D�l��ۢZ�j�Ss `|Q��.y���*	�#'����b��.0O�2HjW�#�������3ZURs����C�����t�`z���vG��n���}�U9}v��o�vH�/�a�lsXv���{d�2������d��$�Bq^�%L����w��6t���U\r�a��A�Y���@�u+u��=���߈-I��V�Q2^ʈ�_?����ED���B�[�|LKֳI0N#M銙��x�l���¸fs�O$6�a�����đǕ-=�.�:���J�j��3,�d-$��J�Tӝ����t�2o�L � ���}�yq'a�<�ǆ��$�rV����MB����+��"u�o��BR�~�;E�I�#ŕwՍ�H��{�ѭC��Sri�㛡7�����?��ÓyFh.@�Q���Qk�c������b'9W7I�VÑi�kk�_<_\�;SQp_%�K��<J.�����a�;^3��a�v�� �IG��b�wgT=0��j?�	Ė:	��-�`��ת_�:uBt����ט�rA�nW�ƿ��B$J*1�;�.����Y��.���)̙V��w��	j"��!;|/.;�g��Iё��0�N^9n�� q��m] ��9�a#_�c�qUp�T����!f���b��v������2������%��i��`N ���̎�m��:lPyf�Ğ�e����o���!�ԉMW�M����k5�q��<�45�7�t��q�1P�T�U��3�R�|�n�}u� E���ʄ@��˭S�<�i �hm�Eg����yQD���;R���!����a���Y0��*��d~�h�Nc�\
[K��b�YRֽ����'�bf_Y�_�2�qOO���k�C�z_��cp������>ǌK�"�M� �$o�M�|XB�e���ݔ�����b�w3�&+6�10�;��d2�G!�NR�,�TS^"MJz�Yt�+��>댰]�J҈o8Vx�D�aǹ/>b[�� (�0����h��ٽ<ܙ�}tbj� W+GݎV�����O_i���'y�3����E��
z~0�\�8�c���@�8����Rz~�˜�jYk�{�+�Aj^�M6���4¿xXz�B����mX�ˤ�|��nҬ2C�o��A�$ת��+�IA?�J����ԄA+^�C)��r)C������9I�:�.(:��dĩ"���K8�^�������u��[*��v��B���ĸ��l��ӣs�4�
�[�E)�
�o�%2��Lb�1#9F�3�����,W'��c����l5��!rX�PD4½i����'̀�{C���o��~v����ūС�&ρg����O��X�J���a�/��v�1��t����:X)��ڮ&�&�D��9fc��,�I�:��X����\ ���q�^��UmYlV��~�`�e�;��Z��/2n�:�3y�=1C
��'� �Q��S:2�q�|�f+&-Bp��t�e�����O�EG��,�Y� ��%m�[�!�� ���5 � �8Ku�~�!*��Aem��i7m����8��7[���M������u���ۜ��eJ2��\���>�tK�7�A�4@.C�*�Y��W���,�����\�B� ���d��6�P��5�E�崻v_�^-���	�	�z�"�"m�j�xs�����1���Ʋy'_VFELѩ�鱒���K�����(Jh�]� kQqph��|\�d�0���<�R�)����5�(�o�j�,�J�����@mf*�c�MMj;p�kj�<qzK�_��S֥`H8.���1��=�gͣCnۜHFrrA[üu�,��d�d�O_�-����QQ�̮�2X�ʱ��ȹ�<���?�'G8��u�ʺd�Y�W~H�ڤM6��P8 ���c�aet!��r$Ռ	X�.t�;f�FWѡ?p�L����*o�����9
�Hd{�?Ԝk
������3�7?>�S�-�Zi���R��<B9/eu�G�yӟ}�:t5_�<s��\�L �O��s�#�l@�v����i�f\ӍH�X<1ZN��!��
R�+yG~B}V�B~qW���g��G﹒�C��@��8+����oA��"w��9��xz��t`h;"n:�����`īV�X��o1s-�D��.��x�pO����w�8��Q��v��k��A��Ռ��9��e����'�t�6:�_JE�������Wy�(/F��%Bҙ�P(��L1�?[��*��%i���i�����*�M0B��e�t߷*�6��j�Co��h`Z��Z��RKq�8X�Stoܧ�O�z!���ί�4Np��;�����J Ŕv�i�S<KB�,��cX�Ƣs� �<��'+b�\��e�x��e'��)'=��\1�5 �w��8s󯣿6��/�A� ��'��N�Y-�5q</����~``*eŮҿ����m��]��h����C�4�7LW�0����ք�5����؂�}�^�C^�b�߇R���;��06�#���� %x�U��~���R>ꎀ�Z��L%��{v��x\O���P��h(�ZfE/���(U@��B˙]d��{ �,�u���2kꃙ/���һ����
�_����?�ڀ��Ev;I(C�~1}䊥�t��N �i�U�nw"v6��#g� �F<fY�G$��3�tR����{�/om�5���P�g̵��x��ꖣ�Q���Q���q3'sl�>&�D�%^k7�_�D~b�:2Z�1̍�8�,��=��
����q{A6���#����ҫ��/�v�9��4���Hp��p��T�#sI����l�f�s�{��XRA�� ]W�@���D�0�B6D;�&��&�5�m��Oµ��>�8�ܪ������DDp��K�Z띡�s<���`�R��4�k�����1}܊��C�K��{AY�GP��C �fs���U���b5j�eh�X=�ت���A69L�c��?�Ӂ޷��'�m�5�+��%����C&V�Ė��T\��`�pK���ڇ�����?�ұ�w����w�N��S�"��N`������t�ml��/j��?Ê'�Ƌ^{�^�EʾC�Ю�w�R=v����a[UG��T馧a-�aIMj˕���Ĺn0� TmA�����bj���$�GT�_�~_F��'`U�H[J!l`͏ ?�<�cU��%q(��Q�f.x��GJ��GJ���J5Sa�
L8R'����O;��Nek�U���^�h!jA�,�����h������+�:��Y�u���H̑�������ud�j<]�#�SP
ty�e����i�'�ОԸ�5�=��5����&(�� �-�9L���B?��?2q�ъ�����ҳu��%����,�K�T��ӑƂ���u��¢g*��l����o���FZ֣h�>�d)�b�4d�s�k�%�Ev ��
���w�hb���Jh7ed!'�<��
�6G��_ v2^\	��T�Ҁ1݆�n��ߵ��#�L�tv�Y�#I�(l6�,�W�cS2Uqg3��(iY�۔7�xK�Ɍ��OO.����T��"뱊�_<Hz��AE�:9X��8Z��U�ld.DS_Q����bߤG���\̸���Qu��g0�{�|ᤰx��[��h��o��2V U>���H��3�j��؁6U�������p҃c����}��*Y�.oS�0x��]X8�@���oGUd��Y��u��yH�3\*b�ĝ֎��P�6�c�}�"QGK�� �%?��NfsT8_5�?��Bo���̕�b�#u��ӳ�F�0��mt�[g;Tn�!���$0U�����<椠��gD��T��V��A
�3�)������@��7O0b��pL1%�D���.��̒��C�'���^�⟷��P�B��G(i�m���ոd>Ir�����* F��i�ё��)�3� �~�����ѱ��RD05O�<K�á&v��9;j���`e�[�� �4s�0���e��5�B:�����ZTꚁuf^�{3`��)ަ����IL���i�_
���۱���bx��и�>��X�2^\x(��h�KU��Ğ]/�bnˁC��dI ��_ |�]��c���Z��z��t ��JM$q��iC9����HN\8�f����i�>9�j��	��QL������Xj�o�ߴ���.�J(�Ǻ���q;<�pJG~�K!w*s�c�S�ɽ�:�Tv�nT��!�~9Ά��
.A�����L�E�x�va�0`�v#�t��Ly��i;���2:u���Y�')�dB��Dks2��$k���9��Jo[ڏ����W�Q�JA=<v͍���
^�T�J������4�<�~��f�6z�Uq�kR7�R_zȂA3������/�������rO+�`l92n�_j���#���F�PG=�1C� �S�~���Y~�C��������E��� �3�O�oS����qt%��H��?��W+�ߕ��9����a|D>
ڌz �o_u�.���{/r��ћf߲�:�x�&"�s
΄u��� `l�14�S���aB�G{���t�'���1�.P��e퐻�Ѱ_,�$�[հ^M�M�,���r�R?�:	hF�-��hC=;t�+�{��LKs�2*���)�K��m<�&������M�IƝ2w�ɷ�7�b�5���xf��F
�S��E��ѱ!7��kC��|杖�����Q&T*rщKX���2!��jL�I� �i�y�4Z�[0h�s��?�!)=AC��Qp��a��_�3��RI��C��f@�'|�>@�@��#6�ୠ�鈨i����C���gc)PI,�@R���ҙ|�����,g���7���Q��s�0�gŽ��$c�ZV�`��2R�6��wV���^ ��	��<B�(B�8���4$�E�ހQ)�gR�%r��R׆-7X5;j#�Vh�F��1ֹ!�>vi�!qc���
��%�d7�A�X��NO�߱�P�O�/ڦu,���)�b,�2_y1��ks#�|��r��I=Q[]��,��j�E˙��r�}9zZ������c�ʤ|ʉ���*3� ��e�#"�J0������/zJ�Q�?�|"��}��TX�;��K\8h^���4h�:�~���*e���Ђ(T��eO�ܢ�ܰÔ��f=1L9lq�9:$/������G��It�.������{�h7�B/WZ��D%?H��4]'��DC.eK<���-:%+Zk5S�r�� ��ş;�q��|�, ~�?��Z�C����l�jj�Т��T*�{nG��E�pH�{�����h����ԭ���]*�"$���B��p�Ys��U�-����(:.�kG��c����K��%��3��p%5�4E�~������TvJ=$�^�Ԡ4I�Ǜn�\P���-1r�������#���_�Gfj#L	�O���#I6����JN����!ۚ�����B�+��L��I��h�[���g	�����e�@l�%��[�"ř��+T�,�հ�a{}��盻@%���ȡ�<��R�ԃ��ަ�u�1��rX=������E���nf�I�:��i�a��TH�[
�
KVx,Dl�!L�bw7���P�5jG���~��cQz��K5_+�h\��\���G���q@�r�lWOm.�	����F�W=}8�
i_�s`�db� j��*F�7޻ر�-��6�6WD9��t\���o@����νx�4��� ����B��lXꅹ�	w~�M~��v� 1Tl�c,Ӱp�6u���)I�lB�ߠq��
�`��N
W՛��]h���n����S�Dbv<K
�0�:���
Ӳm�<$�����u]^ǟ��L�𐚣�d..K4������I��M;fŝUr�U Ǹ�&_�H�P^ѿ�����=C�Rk�P�j�bNeh/���x���I%qX�ţ�T1�c��T>	*♎2	���qÆb����zD�{�HY��*���x㪹��$��JRV��6m�w��$�]�8V��]I�'�
i�����!�te�!��=L��O�\]cLσeSK�'�����ޔpc�xKչj�vo���":�Hl�v8����4\ʀ�+���,��8��И��g�����w�`5����y��B�"?o<xK�m=�hL��������EW����58�A�U�_���QnG��n�ͣ����Ԇ��k�R��HdsY[xJ��C�t��M6}��	�6��
�*"�պ�%o�U����7����x'#5�?�su�r˚N���'�3Y5	��!�|:��n���?�=�Mʔd�N��ޚi�[�{��e����GK��?��K#I��F�O���4��TÂ�,��l�����Z���^�'>����(�3�C�
�>����@��T��F�m8?p��I�>Z�}�m_Ws�i�{�#��?��Yb���Z�s#�L�:p~�9q���.?����M b�5{��`���c�[7	B�B�UU �R��EeY��O#�R������g��g�5<��KL�����Ց��හ�,�&ē��c�s#�9Q��G%o/j
ڶ��6R�ln�B!
�x��or3����#�IO/1@���.�w�;p,JX~T�pAԗ�  ^���=5���2��k�&%��@�9����B��m�s�`�����r=a��������$�l�&���g�j�qK�
���4��C�k���s�썳i5���э|9�z�;�r}3F�[��u������m�%BG��>��Ӭ-��u�P�/�	WE��A2آ�ѡ_��V��e����C��s6��G� ��3�`oY�t�7N�JTCৢ��?�Y���?�z��si�l�nQ�QT�scj^�\��>�Zs����F�{m�W��v8�Y�����)�hJ�ѫz�u��7���td%���=E[x�5*�ad�T5G�@���	V���ÿZTC����AIC��4�,����܅�C�����]�S���q�\�~<`fS0�t�aB0����`���(?=p�F��]CV>�@��R���?�|`5GXc��eŝqE?�&��z�1��� �8�k��ft�ܡ��\��g4�����
�	O^/�f�J]'����ҹ��FJ&1Ԩ���9�dw�m������H��rP�TQy��r�J�����%�'	d8����*k��_�� ���T).D]LBr6�?m�FF"6vS�~�~����qAI�����������38�̹����d��c_<-.٣1�Nܥ+�w���$�b:%ӻ�K��E
����JWp�>GQ4�O����M��.�4��Z��E��eV�L�q7�.�d���>r��ک,�yj��|�݅pb�ŝ��<*�r������:�.�b�*0������Fܳi�ȲSr�엦��q�γ���S����o�TBEáܣ���r���b�|5�>MM^�)�14��V>��5��/L� �}W���ڽ�-�-y�����$��
�p��\�X��u�a�^h�45�SKYj�/?>@3����}��)ò�KG2񔟇�cv�_҈!PLé�s�� ��qӸډ�@6l�jXh����Ҙ��v0�[8�r1ŏ�/��C�_���,�������r0N�d��\9 \C�J�*����f4�8�G�)��r�1k����&3�Sm�1�8N8������;pe�:�j[���{q��P򉋨���VC�k�3~^���Ks��MB�,@�J�1��$ץQ'�8�����
�b�sA�ڛ��#4(S�7��oc4���N�>z��|���0-|Õ�N�:�Z7�s�{Պ<�r��hQm}GB���!(U?�Ӎ�r�xK�z�ڕǉ	���m�QY��� ����(��o����{zp������ihXjs��!�1�)������S��c䭇���NT�F�k�ߋ�KC�2�^pr�M���9�w2X�_h���>��Uۓ+sF��y���V�i�ǂr:�i+�g+4�K�԰_!5��6���Oa�%���#����Xr�G�"ƨ�5PRTV�ی��l^r��S��Ѧ*
w��%K�6�^
'�R %4?aL�ɞ�H����W�|����
@��F�AIOp�����W�K�g�;�`	m�4w �߯kU�V�聁�(�+3F\���	��옍7�+f�\����(����
�-��fL�̑D���k&ω�d����E��ם�@�egR{�-,ɱHR-Aȫ�D|�jޣܵ\�u! F7�4&�z�"
��Л��z�vK�>����}'O��j>���TZ�b!%�T�Q�{ݰ�8�c�?*����-P4#�9��O n��xZ�ayW����e���"�r�����<߳����/Y��nn�6zf��n5vD�o�aeL².Fk['���%_@k._T�P#�r�n��=��yr����6}�<7e�V�wzhY��b�úD���80"�*m�5% y��/tb���z^�&(*ȏ�u}��T�%�I�#9�e�:Ϝ;�B�}0p��l�_��x�O-D�@�A#Lk/芭�>��o����=�#��w�,8.��|�u��Qm��U�2����5���ǧ}��4�7�H��b�^+'Mn�1��r��Gm1cӞ�Ʋh��>�=�#�]�0�e;�c?�v5V��q�Hp0ߨ�%�C��(>a���qъN��&t�RK�����`b���hf����tl��O��*�'��H��)��)\��ZpZ������|�F��`��M���3hg�f��B��7ǂ�<(P���9B)�j�� 1��:#l�Uj����^z�
�@6�����{H��.������|xu���o�	T�������	>� �jp,��&��u��q�F�CԿ@��@��K�c�U� �����s-zrf�)�Ȯ�>s���W�\� �H;��2J⏽OZ���|��8Wݡ��H6Z>k0b�_��( 1	�}z��|B���9%�'�X5Ysc�����S�mJ۪SĲjb ��w@19ɡ#O~�\S��Y��1wS��F]am`�=E�H}6A����"�)o�=���y�ߡ~)�I�SK�&�M��\��C��A�N��wՏD�E�X�(����/�H~q�R����2tr��Lؖ��`*��n���5�cfchȃ�g� (����H�d��Ք��'ۥҙ�D�g�_y��d� K% �TJ

<@�����E�ا��j`�@�8"�M�����5�%�0>G�������d����'�Q:[V%��%�V�6�l�i/��FG�eFȉ�����d`�CU�uI8�*�g.kt�(*�,h%�o�� #����(�������GR��C�/�����ܧ���f�hF\9���J�Ӈ���cK����n`��6�&KM;D.mS*�5�l���U:v��d��ʫUqd��:A�(YE�]�Z�ߛ�iEl����]�+�%��I�`�˼Q 31n� &-�c]�O�ZעUU��b�Ǆ��#�ɏ�\h����@i�����|�5|�l��W(�cQԠ�+"w�#䭸��W��W4�-���C!G�0��M+��h|xF%I���W�CG�Q��m5^���1�{$+�D���K�d_V���u�T:@+��$����%�d���ɬ�b/��d:�:��z��K��"�b�/�Jr~�n��KWZT�*z�ڸW*�^Q�p��%]fZ9ڠC��k���8�م�k�'��Kg�Ʃc���1�f�.�7t�GF��z6��0!X"����'W�e�s�.�2G9���-*�M_S�v��BP�p!qsU@k>�� 5��@~ȇ&*����:�^�7f~;�T�d&�Xek�@�}{�v=�����f��yt�8��IG��i�|��Oc����U�	'm���0�fӯ�д�c��{���巜�I4_���+w�T��Vfqm�_����|�S��V�id��Wg���f�ԋ7hN�������H���	�2@h�ج�Q�_�V���b�4�ļ���@��s�ˌ���n S2#_���T���I���1_��)摴�������!.�Vʺ���,Uލ��1F\�==IL�\k0b��}�Ʒ"W�T�jt���k/�5�S�\_y��dl���Ė\**��a��lׂ!%��^�l6�m� G��n�I���xi����پ��ȏ:���T`2S噙G����Q�һ�Y�p͡�b
��, ��l~�!tF��8>�M
��e:��<k.�#���� �)#�8�C��f�e��#��4��(j����xp�����^��Hpzs��胃�5+�s��a��5ձp@�+�ȗ��I���?�yZY =�_����w��@�m���4�5$�`���P84yA;3��} t����Sǚ�P���V\=��o��ܞR�=7.�¯�X]ѸR�g8�ev����+T�����wc2NN�%V9���;)a�����1CSH��6�a#�|��y[�O��5���_�=;g�W�]1#M�5�9D+cB�}ˌ^G��PT^�,F��8&#�p�3�8$�E� Ѓv�uV-5hG��R1ti3��\x��ȗ�5�M䫛����F���/�SZ�$ǭo�&��)�8}�LV.�E��2n`j�j�ʉ<��K7Z6tV
wD���O�	z��K�&��Q�_�![Lr�h�Ⴑ\2�ؑ�ʐ��/������c\�{v~���x���+D�}bb(f�fP┈�ׅP���H��r%ū����3�E�{=^U�����>�$QE��RR+����R��7�|�u]��o��������!��<\;��ބ{"�/���ۏ��*�=�L����B'.�"B��2���С���Z0����_�;�����g�$!��*x�2���'�N
���-�?\�4��1Y��,Ug�8J��c.~��
l
k��J2>��6�&rX�˼T�ni'���Ug.%�#P~A������.�J�A�n#�T�a)�� ��ԟ�v��nYqA��$͟Q,6[^ .��#�l��U3��Ii�/�ۢ�7;{��y��j�
�a�T�N�A��fh�	2��3q��~s̱fD�,z!٫ˀ�3Ԏm�B��h#�{��A,�w}���!1ko���7@���!��2-!I4��%\���������h��b���u�H
�X�Dw�� �~ud��G�Pa�>#ц�թ����x�3��E��M��wzubK&Ⱦlk�<3�$� �&0ȝD�*��]�ƳW�+��?��UZ�\��>���U�����w��]�!���ީ�qu����(��d��^�ʴS[���A�}�IH{��z;D���&Em��k�6�2���/�A2	�^�t�����pP4i�'�ɖ�O@+'k���R�'<_W��-������w�o�ˌt�@��t�*E�`#ՠ�����4]@��y(ď���9�*�>��	�jm�������l��O�\��Ն9p�I8��k��!f�9��Z�6{��"2���s?��(G�����)R+�C$�፟e���Xl�1�wU�I�H���U��׶nb�Oa��g�~��
��P3�����>��3?��8�>�9杂2�|zjix?~�inx�!�	�mGy 㞘��?��>��I�w���g9�"�%&0V�ik������T�X�ٚ�X
� �4_�p�b4�ȕ��P5���9а2���DI��>b��d��_^S�K�P����%�HAou��=�!P'y�3��=�BQ���;x�=�'4�S�-��Q�9r_�z���=�����%E�60�'ؘ�[1�V�<d[WGo�|>u�'F�ˢN�S,��
���ď2y-i�z�N�w�T�f�!%G�C�jae�l�|si#�5�G�W#6���3o@R���߉��\�����x��@Fl������U��+m�z_�"��|�A���ҚSx��F$	>yz�{����'g�`Y��^+lNE�SS?*�g�?�
P��.��R#�⩬ �I���c������ZE��{���.h�X��>=|i`�TƷ-���ˈV���G=`�H�,	�����:��+x��>Q?�&� T�.i~\%��-��;�(/(g�O�I�������)b��ҍ��]����UvJh�������$FG�������/��3@f��l�I��9�3Y9����3)��蘼�B��-�唷��\�6a�W
���!��W��D�y0�+�$\ǖͫ*d_"���0Bn�D�V�=�6#}3�P���i6sKކ�����Ǝ'���ynCq�S"`P�� �?�����}a&���,k!�d�o��"b���L��[���|z����{�pyH;G��{��s�E���#W�%ǻѠRJ:/�Q��8PU�z�o[)�.Xt�3�;�����3��pAI��F�Ĭ>	��8� 5�9$��Sh#GS�)Rq�#�����P%p���F>i�E�4:z�>�4�N�iy�|kv��r�>n��T���IB�*�, p�L�옣:ڎ�׈D[��U���<�y�z#d9�O�i�k] ��B
á䙗�$6�Ʃ7�q}��Hd$����C�g��͐e>�v'���=�kȧM*]CP��S��b����eg~�2�X�Q�Um���� Ȼ0y�}��h^%N�=�4].)'�&~�,_ೌ���y@S�h��Pߒr|����u��肿���P�&[�����i�,�]������V�8UBn�F�&Y|���Ӯ�:*v�3���]��LoV����$�{�~X9���9��~�� ��AF��U$[R�g����3K�wQ�����+*�e�t*^�����LCJ�+��r�A����&d��Rk�v��<Ƞix9!�m��ww�Ya\�ϖ	J��t�i��L6��r�2�ncQ�%"��)hv�i]���X	�#S��z�d킄��ktA��kDaw~*6`��x�gY]]F�Z|�sBc���/s�*�Sa&��#�Jn�Y��.=a~���mk�a�Bm���|�+Ypa�0‧����<{�$�D�qyj�����-	�A����G���'f�c!�A�k�����Ԁ�Hfbܩ��?k������?I�k�%��:��		r�}��6׵L��.���+8iQ�],쩎�Ϥ�ԫP+�� 䢡%�wN�-���
�`4���&#�:�t#~]%*����_�@�I#�ҝ/Y�X���5mڃ�� ��aP��9�6����dk�a���j��]�$������ɓZ�����K9��X}b�`t�D�Z��e5\B��Z ��)U���]az��Yf ��E`W&G� �ʸ�l֫L�65Q2~�a�����8�&_.Z�����\�e�:��-��5`�e�1Ŋ?TxXo$S܂��i7|�p�K��= ���ߨ̌���}�|�	�(DT,�����$�z~nb� IAE+Q���z�
��W����bm�1�rr�E�㒅<2�مH�w�-30ȿ�m�-��׽�,^��O�p��zH2m�k��"��I�<$�҆��f.3�����fp�K���H����,ā��Fz�Y��.��]�MO�	��

|�{�?��+5`$0_���Z�_���t�[�~��y�{*�)��e(�Q`���y1lM��3h0ؗK��RF~��g��$�R�!j�2M2G�.�u@�%���WtA1�m\MìBo�W� �J��Y���)C߀�$��8�
��J�?#U9�0�g��׭��,���3���{�M���)�Nd$fm�Bt�X�K��s�L����J�T���J!u�5Z�G�7d^�rM���̈�	����[�����y�	1���9��ɠUD	R��n㪻�:��I4�'rr��T�k!��&;�D�E��L?UU��K&Ȓ�O�rϐV7�N��3�R�ߒKk
,p���� \���ԕ� u���!H
���oۅG��髾H*�_�nH�|�6?�*�?��a�x)O�^����1�~-��[� ����8r���/A�Y���P|c���ѝNd��֫F�]���k�L*���@1|oi��ٝu)
T~j�d8������|�=�|SF��9�EzO�tZ�/B�"�� 5a���;�J_�J,'?w��G���5�P8��p��������\�W�L�ԧ���<A�0����Q��p�O�����2�3N�;@|���W��z��V�mk�:��X��3
����	p�XjZ��>M�s���_�����DTW!f�ɨ��+9��n�ɹ濿�tHCv�q��d��T���x�di�& q���Gi��v�G.=�"~�:@ ��T��o��>H$�Q7�iVZ<"Wws�dO�1�҈�no�ߏ�*�e��%B�Ȣ�ML�;���-L䞏��MBﴞE�,wDGf�C� ���E����%QQ�}R�O["*�������;}�!��wk�K�Nz�f�jJ�1�S�]���(��8���KX�Oui,�$���:�\���~֠x���?.��[߰5�2��٨���|L"v�ޓeFƢuX9�sj'�	�G���t<S�g�?�R���4G�r|ܮϨ�B�o�{�����R���̇[i�f���a��ʐ<$}6���Il���"��Jw<����B�5�WS��i A��ў���~(�� pZ'�AL1
��* &�V�,:
��)�0$H
N����9)��@����S�Wg����F�Q�)G�i���St��7G������S��}�1�n.6U��P����Z��a��	�¡j4��� ��uP���f��| �N*�e\��0��vӯl��v%�����ƀ�~U�9�C��������k���k˟S@�QZ��F� #.�ù��v�+��ٸ#���8S����#��e��#}�;�P�6���en.�'�nzK���3Κ��/�LNR��9|��럖����<���V�f���a,����A�|<��O��U�_�c���n.M����7:o�Ŵ�,���!�����T�n.M~ܪ=�Վ���k�3z8��{�����^ �E��pK��Lw��Y}u������kE�M���q���9{w���P��zyՃ�F~��q/�t�s�����g�;���(w|���;xBH6�L#}ot�s.`έ���yo��X��'(���[�]S��[�ߕ��`s>�a��'P��R2��KZ� 6?���1B��l������-3f���kN���]���Xz��biT�}�{8�0�^>���ߐ$-�E�h/2�F`�� �{��`p���QRuwQ��~��k���#�1Z
Cfw�2z�W4S^�)����*9�����,~�,�Ԩ�?��:���$��6�do_��XY��|�R1���FBƁW=�a��,���(��~m�	:*O�/#�FxX��B�	���m��pSq���]���P8~5U鑿i>hL"�P$E��W<��U�A`��E't��J��	�}l��e0?��'7�>�/��zc��Bà_������q�*�^�"����௶�g7����&�d�_��`	,^Z@Ń��ZD��0��
�7'!�yK���ʶB{/A�2���)T�̚�)����1����/�l��aǳݥ2*����H��=��&54�h�>�5�/���)oD,f4e��!>R��w:\?]��aG֫�m�<�ғ���Mu��.6�qc�]e��h�0
I,��+u ��<:�Q��Ԁ4���C����L�!���״3�>W���6���t:o�\ X��Ɠ�4�-̋�{q̐�iLs^8_��l{��Tެ�Qx����C>�.�E�l��0u�V۝N��`Y6M�ׅ�{�J�8G>,��Mj��#��X�"3D�p�qa�o�f7hD���B�����mO]�&���\�l��n��o(�Ë�|�~.7�)�SG�����7dr��Uu��a�]��^<-��}�|!HL䖪�!�Ü�7��l�O��@B;��h]��W�����UL����s���걻����͡�E�g=x+6W]q����
]z������ [_��F�����~�<�>��ح�'�O޻�j�:v��;ow���N��l�����&
�i��5�VKU���k�K:��g"]x����������8�����J
*M'��aO����M3#̭��5�+��'����q4�$`���f8?�*f���A�V��wk�����#8VW���Nj۰�H_��-޼s!�ΚESC]B�c���$v,ElGT���Q�>�kw�n�������U������bj���6���W3�������B�c����X�D�$���%�{3`�Vz�,���/����dǑc�no���ʱ���n���#�ni�o���K���@��"��x�
�Y��Y��N�B>ת9���+@���#��Q�px2`GP���%�39�*IG[H����1tA`$�������=���-N� ���7�Ȭ��w�'��S�M7V2'��p���:�����:�̣�(�oa0�
)��ߍ�]�B��G�0��{x�q�X|m��I�2��M�@��� vQ��v-mPLOk]�ʌ1�U3r�ǭ�������\���	sy�?}����2��!l�����	���hyo�)��-�e�2~h�H&Td)и=x��3o�V>��}T9�C�8�Ai���\�p{�B��;�R��V'n�-�J�_ă�Ξw�QP�JX���p���W�o������ ]T�h�L����%[#4��I���4�i^�=�%qQ�A�><37+|9S��r]ݘS �ճm!�`����%��c,.��$Rv���D��T��1����L%\:�{�p}���x ��j�^��Tx�C��m2{�EeN �����������&.I��M(bhgl{��������.�s*��'�ڢ<V�ְ�B���:���22�_��\nF��O������G���! #�G{�P&���a�k�bkJ�.�¹���-�E#�o���Jr�eRb0�>��ҥM����S�w��qC.��w���޵�v�K�#��<Lh��f,\��̳�NIƫ��'�Ҍ�OT.5J���q=�������r���?�	��۽8�9�~�Fʩ�2�$�[�U��v�y<f��o�F�h��ԣ�;�b�L�h��9��_�~�G����FQ�pG|.-މ<{B��"����4��I�0zp>ݢ��K?�I���V�س�'ƗPl���g�u����h)-�TRj�� �|�F���P3�?+ι�5@-��c5��ja�
_�ʲ��%e�HN�`Q*�V�Y<�v�8+P�Y�3~`��n||�g��*��(.�Q>�|R/|,��)�?�ٿ{M������䠩�C�P�˗p��MвӇ�_G�:+e�	%{A/V#�	��'v�ξJ@��L�!��2��w��ș���9-��Uc>�`��Ϭ��>���3��ՂB�lŵo� �<_��'���!L��=:l�+LX��������-	fy3���Ewze 4�J��R,&�B�y�����Izj�*�ǛM���o�>�&��]� ��6�Δ�ǡ\U�	��{Ϫ�r�\�Ln�ɐ/��tNvH�
wā�{�y�*�}����Z؝�!�$��(p���Ci>���Z�c+�8H l�E��^֙!��ig��4�L��}D(d�*S�\r°Ux�������x�����ؔ�JV�xH!v~>Ʌ �_�	��Jڭ��[ѹ�J�|��&�R�C��k�"�͟2�D~׋�zZ\;�ܦ/����@ڭ���ݧ,\�������y�3��ٻ�L�MC�X��Fu��(����O>�lH��6 
T�H�`�|�Ȁ�-Q�櫹�Ep6A��O��������9����By:� ������k/l��|��@ ��.�Qk^v�fz���)���/i6��w���T^�`�9��Ð`�uX�Δ�/:�c�1�Q+�{a޵��s�����ZD�3���A�T���]�Iq^�/����2��~���{%QW��{�1e�i��\�'��#�KX�Qa*j;�-.�`���QfBq�J��Lcp��)�"��ԙ�p{�����-�iEVa4c��>����cq�ZSQ�~���ҀBH����'=B���|S%H�Y�0�e`�t���N����~{+mL�*ebqI���+�
v��+��R���K�4���i4��WGx��q�yT{����U���ܞnzw��oQp�b�y5Ð{�2h��]/�TJױ=�ߍL��mv�7)���Q299c���L�K�2ͦB�~�U�r�C�j�Sޚ��dt\e4,l����f��k���gA"�����D�6��S�Y"�^`�9�m���,g�D�ذ��6��VC<���*��O� ��uS��=_��6"��!�Ё�c,�ӆ��#If{���n5�J�$�b�d��9�&�)Q�o�C��(���Z>��0'7�=5^�x�L�YQ�p�0|HR�K�.j���>��O)qp��!�Ç��pC	<fq�`)VFZPT��(B*%��+�j,x{ y�z��,�DLX��#K%Kp{�
������`N;�V��Vר�����+�kց�^~&36<?n��d�8u�M?Os�%Ꞵ���F��_Tizz��0��<��>WǱ&����'&�gE(������o�,,u�h��W�[	�6߬�ʖ���Q��A>�K�U46i;Z j���_w�<�-ͤz�M��y�	+�+ �?3v>�πUR�< \�P�I�	3)�0��$Or~��+s��˲x]���"(�(*�G�!��s��Ҥ&ER�m�/W��-:Va���p@K��ǉ�%!�o��_ݠ�etm���ڸ�
��w�D��?C7���ܦ`GH��y���.�%�Q��I���B���G3�)�l�T�?�w�n�! \1�D�߶��|e`��*;,N���s�
��5�/�U;3��M��4���BVm[[��g�����>d4}k>,�v��!�x�KZ���پ�nR,�
V�tj�g���g@G�����k2B*:J�E)�D�>�l�k�-�C�S@Yζ�h#όe���d÷k�!ǁ�a�7z�����.9�����0�rd��e=3��[:����􍀝v��y�_I�1��H4Ĕw�t�h��	+C��z�/{��;m����Z�3�+�ۗ��{]�YR��rW���^���sU�8ݕ��8���<�c�Ew��V��+���΍p5���AK�G�U�n���V@��-��C�q
 R0����R"��\/Z�{�}٨bצc�g7�����}���l��+���<���C�f����ʶ����g�1-�f���R�"�jR$S�H�͍���а+�J	sWi�у���=�L;�}���"^|{�3�]7L�,��qg�}���b��f���	gE�8���'�7��V����<��U�Q��N����ʓ0S(O:��\��z��MI�rJ�lr)~�:��n&]�f���k�j�`  {����`g�t��esD�-���ߪ\��c^����IU���g?�X����I�h'��w腨0I���I�F����Uk��Uք�g�
�67��I���q���<E`�"wK�z�<:�ق��5��S�Ġ]g��ܑ�b�VkmB����u�]����D�D��m�em�X�f�߱t�SA9���X䴛�wނ�Y��"<~������!���n.M�{�� ��'����FvN���{#���.�.�'��kk�_1�lߒ
�u'f�dU]�}�Uav�[��m�E$!���	Ѷ� �M��!l��f⤤#k3)|�^��.���"�}��̪�q�}�-B1��I���ָԜ4���m�u#!8������~�VF��T������pX��9���ڰq���,�D�M51GaB����n(/�A(�����H��7���%��a�]|/������,�it�����GZ^\e�=��'=]���8��E��F�_��BL���=x�p��<��N!{����h`ؚ��3s��5K%w��T���)7H�!�{E}��6z	��>rs/��,��#��Y?�i$>A{l�\�ְ%����{'%�d��j����r�`&.@�+#�z�0	��ԤMM\F$V�	��ìh�B��f'�| r+������N>/�3l�CR�W�f(g<������C�
��>E�U;��k),��`p�$8�:Qa��W��=����Hu��t��(Q����7v�?U��/�c�Γ�.2K�O�Q0\2��G�9���
�cu�䀹��+kr���N"ꎈo�`�����A��r���;s�L�+ڼ>����|\�/$��$��ֹ��sw]b������H�u�c}�n��3��dc��If�%��������^�!�\<�y�dӖU��r��k�E��4�πR��:J4+�^�%i?n�|�<n���g(ي�!��?n`EJ[R���"���qW9P�@EB�4"S���ɫ*�T��ۙ��fXYX���+d&�5���+m��^	���m�s=�R�	il��*Ե��Q��@j�%�(.�ZAp����tKdh�i�',/dW2��7��}8�F��tH��Ȫ�4��� ��,�G7�+,�L_z~�~�(�8�Q�t�`��	ߘ������-A���?��#.#�Rp}l���K����[�;�<Ӓ�v�H��A	�3k�^'혍3��0&?�\���T���oPB_�<P�q�����+P!s��
J�����8�h����$��a��/����I�?�yJ\�cc\ZY�B�����w��\���s�����S��7�?����\,��J�+֟lD&X�p�u���qX�e{���@O�X
𿖳!
��F\� �s�)������U�Y_�a���N��z��*�RN�u;��B�Sl�u�=6:��:�8�|k*�Ss�ޟ�a�4���S�s�0҈�k���� ~EG��I|(�,�um#�}(}N:L����OҾ�?��`Jcn^
+Dߌtm'��T����e�.(8W�����FR,z��Ypb�2i?6eP�?��ub)0�+���m��OZc)��������!a���`�r��c�1���;�1��n���K��OU�Ar[Ĵh.a���݋���S���;�u����Ф�`I@�8΁M�$�
��KUf��R�.x *�+/U��%v�;�%@�5���*�����kN`� D�l��*	H�|erF �K~[����sfJc����>�G>�����VU;�,�t���+cd�sY*+��!�m�c��^\�ꐨ����ѭ�Z>������Q�^7m���la=,���ǖu���[w�B�+�',E���S| v pD�Y��\#ܔ��s���b�U9L�e�3�o;���N��7�*����]$[�U�N�a�񻥡��;w/*�<9�G?�Ԗ34��6NE2�mIP��m%MR0�������Q���{b4�!Ơ�����
3vF��{&�o4����]��G�7�*��)�/z���� i�M&�Vid��yV(�+N͛f�^=���k֍��	����p�<���� � [|1F	�+��gsh�]�^7�v���a�2���Ez�S��3����]�*#�N&��#S���@�����tHR�{�sO����1�BX��%��IFV:�ǉ�h�j� ��&������J_L Ǣ�ʐ��p2��p�M�|rGx�0�G.*�3�l;���7�H KP���ܡ�\r�e�}�:7���Y�.�¯襨�ݭu+H����Mfsǈ!9�$k�j"��U(V�{	�i�a�K,���4��8��"n�H~cצ�e�'�Gj�E�[��>���Փ�mˡ�j�`7F��?�2G�6�
�j�j�#pom�2�ٶh����gR�@M�C�r�b���mɤ�:�2҇�		GɍK�Ӗ؊c�&M�R����$j)�E�l`xf��� ږ�t/��	�=أ������m���3a��"����j��%Ϭ,�5DҪ�x6�*�0~���}����=xtzp���yL�B�aZ��<(яu�����P9��!����X����f��m�u?<r�N)'+����S��b#:z^����!J��7<�&2;w�_;C�څF�~!~�6��"���GptP��Tv�ߝ�Qu��Q��ḉ�����;�V��w����Ξ'�*�0�N���WP[�'��"�>��q�@�N�ݚ�^��a����o��eA!��e��Q�Ұ'���H����·#΋�> k+5DU�;��ܼ&�̈́t���ܯ�CC��<ų^<[�*�h�&Y⢚c�,�K��yF��n]�~�u-�s�<�����P�l�@�C��nE۩>�h���k1�=�kݤVy#ھ���&��<(��++scǠK�i�{��-E���W��̕9�v���hi]8�Ps�=ӞD��M�d7�$>�0'(��@'Ղ:�o�%
6��S+$n'���TB�Kp?1�	ȷg9{o�Jz�R !-����P8�IU���Ma�=Nv��Y_�e!��� �ǌX �q�&U���}a�m�,� na;�=`�p�s^0�����8}���ǅ�ץ�����O�8�qUV:��6�`��(C'~$3wo���Mۥ�#����ӈ��ׁ���bJ������`���3?���M��aG���_e�x\c�J���Z�E"��pP�&>�ˆ��:;�J^k�K��=�������+�ђ�)��D�T!?ޒ�~B���#�vj���#[,�݊�T$~j�?y�l��=��o��"�C�֫�䦎�M+���l(�ʨ�~
?V��n��d�{ܦ��V��o:+v3g�iU�	��������Y�GV�� @���~~��B��b��Y�Bo*���~)(#�����+2�_�j٣���&y��(��݃bC-7Nյ�ž~���|���a���fӊ��pcq։�1��~�ξ�!x��PT=)5r�r��X�Ű;x9/�4P_�uk�"��&!�[�� S�L9f�G��t�ȂBO:-$?Z�N>��}q9���wZxb��P�c5&�
b�+�����H�q��������,�\�)���j���T�ׁZ �����@�W�/�zΙ�~�W�uB�[Z�W��d�`Eh2�k��	�+��]�G}�ǈ���?�7j|���H����:�N�e�R�����f��ق�(U�։A�z[�;砡��;�Βs�y�	,��d ɐ�{���r�֧w��ӣ��{�����)����gqѿ����7�L��2�t�����fx�_�w5>X�'�������m[b4�-}�)jx#���w���J'r�Ͻ��]1Qޑ�]�L{�+���GH�Q��jF&�:d֯3��L �W� �Өb�ڷ�5�+s�l�u��#$�Q��&;!b��zߛ����b��������Ʉ&1�{p/���ѫ�/���~d�γ��h��SQW��8�g����co��8����d-Dz�A�3��U�(�,b${9b��E�*+��}�H/�+�h��O�g��V�K&����4����1w�3��bI�/�se;����L��C(V����-�������*��q���E݋T�]��/�j��$ƺW�td�h|��YN�����/�B�* ?�9���Yȝ��)��e�j�Vj@�P�<<�/x���U!��.�:㓾�_#�Jg��w�I�����L�þ,j���T���"�0
��(��V�\��G<n��4]��2ݍ[��ь��]1�����=��Ѿ�$�B`CKb�E-n�IF���q��,+��1>���_Cj�[{�����͠�]���'*��(�9K8���3!Z�� ��g���d
W�U�;��U{���"�޿I^�չ�.� ��V����^�赭_\h�.1(�t�]"��-������E	B����c͔4��q&�^ljmyi[�S^����	��) ��,���l�6g/_Ś�.�w�C*
61g��,��i5x�fW��s�9�}�:�����2��c���@x�c<b�\�X����K�\�S��;�^ȍ�9�@�ږ*A�c����֒SR�����֊��4,����Z]�#�k�0��!�,�vAKx��,?}+?ܐ-:�=���);�^�vU��>��Ԡ�Ѓߊ��k���iG��Эzfa�*�@�C�q���J̌#��ER���p��Ap4߃;5U�k#�9�/]�a�.���gu[x�:�!�D�I��V%;3�d��T��;�=X��lp����j�I�1^�[�O��8&I�����a�=1\��'o䙓�PB���i����۳����n��Q�WC�:}����[������B�����I:�;d�9{%8�z�0�����Y���C�f$ڭd���Fz]� K�N-���0C������?��-<�acs���J<{�{P�HS�씹*�i�����֩6�SQ]~�;yQTg|�c�D��k.��('������q���I�gJ�}m��pX'��ưS�
W�@+�*
hZ�F��w��������D� ����P�ʅ�溤Ӧ.l7qG]�vu��ϝEmWMj[�u�#���s0�ݽc��D����#�*���n�N���؇�*n0�L��̯?�)?k,D�7 HY�Pw=����.�[��Q�i�PS��c���&��{��WR ш�As9��ff��ݘW�&��B�f__�������C�π�9����c�5v/�7b<�4xq
e9��z��|�U�k�`����t�uh�΃	�qv�c.�n��f�.����Cס�|
j�E7����\� O�P��onR�`��V�G̥$w|	X\B�É�US�M,\���Rm~��JfF3#�T8�@bQҨ�����W�?g��e��[mL<�df�@�/�E�x^S���U�C�k�
�,�����HϾ�p#�V�T�YK��+q���އ�����^�oC�H�շ}���t�bf�W���\F��	_Z��r��(�� wQ|wd��#���LjR���L�%g���$݅i�t��xS�va��	�,;MҞ�
{����#�y ��Ғ�;�GyB��P�,���+�iN������c�ʞ(�СZ������<ܥ��_�Q��J�i]zr/���wi���&e�ߑ��	�>"�J�
3��C>W��2��W����Զ�:���5�9� ��S�ž���K�|�R
�r�'�:� �b~8��X^S��ɪ� 3��,�Z��~"j�o�p��/H6F�C�%�B�A	�"�-4&ǿ�K�nt�;���`P���t:�:���Y�8��8l�#�������|b��D�D@��}�"����w�g6��ZXwqP��wSp_�z�pP�`�Č��ۚF	�M^�'�[����K�*M���S�p��[�
�?6�F1O���{wt��]�ii����H�h��^{$}�� .�}��ȼU�����T�c�x���\�'`/ ��Mѩ�����~J0b�7�.Ɓ��c?�҇TX��r}�dM���*���F�L���Z�/u׶M��	t"�g�s��|��Ճ��;��W��8�� �$P���������������$��vBh ����u���!-��Q��~��	Ӹ65�{����~ȱ�(E����ή�~�+��roƛ�þ���vl�Ι�w�D�T�X��&�~ ��_�)��4͛�ѣp/i
�f�8�c���N��6�;=��Sͺ��Wm���O8����͚��:�o)˫Fɻj�N2�{	��^N���\�uJBf��5��#A;U�c��"���GS�u���� �.6�-T�J0��{1�0jʠg���	f���S�x�qW�mb7c��I�f[�wh�~�֤2��*����ሓf2�5/�a9Zz}g$UP�U� *�9��6�y[�.ik�~N�`ն�}
�2z񲘈SM:d����ܔX\|��FES�齖6�8��8�.-	Y_����<���w��٨b���MﺚeŰ��8@HUq�T���LdB�)�ӆ��R약i�甝��J@�"��p]��c��}���{D�=��V��o�Kf��F���u��*�� �I��{� \]�
�o-*=SK�}�sl�WE���*�	�XJ�K���p�zV�+?G���%L1�ڤ疬�<1���9B�J�"��=b��^���y��6y�_�(�;�M!1�Dr:>�����]9!���f�#숂��\s*��}M0��-�yN�re�w]I�>����!
\�����Ԗ�$AD�ӭ�F9(w�ܽ�hԴ��$�U��F�Z:�r��fxX�n� ���*Y�VWԙ�z�<�&9�K {k�� ����~�|ߔ��@�mD��Rj�����Մz�6�$�t%�!f|0GۚP/��J��T-0���>`&�\ \Z�SUP�� B<�?�C�'��g�g�jeBc��ɈP䬜u�D��W~��O�Ƃ��`-)>,+Fś �G�B�����!�7�M�)��s]����f�?�}�`�x��o�,���і_�Zr�G�9�)�X�3HP���+�o��d��;�*g�@�ߜ$NI�
#wd)gQ�)N����`y�bh4xW���z����R0��D���7V�r/':���],�fma,��r�����*c|�U�T;��LSG��0�5S(�H���t �������35��Z���9��9N���bsT��!����n_�zև�b�yx��Kى��+l*?��8Cl�g���
�F��.@m��}CR1��Sv�pe9�z]jq�F@TX����5h�9��f�2z­u�D��@��h?a̵	C%�DlȪ�y` dt���p�)@3]k"�ɹ���Iv���x�7�����L���(4S��K�����@M�TL��L�$!A{Q���~�w߮��e�vo��=���֜ܙEtr�A�.����6s�J�V�j3�$1�+#h��e-G1��ԃ��R-�I�&8�ﱌ��!���Α{���'%�vU�� �Dx]�3����˘'O&���*9b)T�k;����튿����,����8=>�+$��x��=8s�h�_hAX�C�>K�gd�+�xtY��Cp���9
�cL:#�ך�e�k��4��U�&6���
�MWacb�ʅ�H{�2�.y��蔟�Lz�����Yn��;�q6�lT��[���P��D3HnV<dɹ������O�a��I[����Bd�3l,_s�3�U֎H�����۩�i�͵�Ĝ����&k��	Ǝ3�5����hư���h�T��L��.�
L�}�]��],��{��D{�-�*���F�6��U;�k���"G�-�C'��54���h���eHS��@�J���x��SlB�醆P�:J�V�����X7�!ٚ� �ve�ƿ�_�o��3��������"1��
��g�Z�z���lgn�v��'Y��l�k������r-��!��e�3������n�?٢��g���o}�+�[��V�۫�3�!kh�VK��&6jR��/�������$���7ӎ���kie�8�s�vXL�6�xS,�ZQR� �b�@}�H>ya��������"���Đ]%�F�n,�(�u:���������_=���? "�=�����Z��eR�އ�z�K/���W<*J��Ճ �A�倄�7"g�>�;�{ H&R��|��d��Y�1	�+-X��L�pn&7�z)���G�����щ��֖eLE�HA�i.�������L7%"Ґ�QnT��8�����r��7�����J���O|RG��o�k�>g�Th_Y`|�󤍒f�=�VG������/b9����ʞׅ>cp��Y�;��ʴ!xF���V㋡#�6�hQ<%n�&C�����Rb|CtP���:n[���GS�v�.cr%��b�!S��s�g����{��W���\_�m�<(�ri� 0���)=�J6Sg�64E4Ѽ��������H{�T��Jt�攠m�b}� ��o��A}��1IZa�e������@�_���ApU|���Y� ���7�b|���H�^ܘ��t�#�=��,�c6gZK��#�=���1�&��`\������2����\ $=tY��B~�i����/{)��# ��w��OdPx��{0���Z����.�v�r��v�(������e���.)6j���	�]�7e2�X0P*D�i.Xv�'r��"l7�X��D�������ƀ=�����.�T���K�x|��`�R��dɨ4_�����/��Ӆ��#�*px�D8)Fx�]/�%��JS�}�kC-^���Up���f��T��4P��32�M�u��9s�be`���Z5��F&����h46���'%8i�J���e{\{�jr2v�o`�̺��Q5d��%�u��C$;��Lp�%o�_4���;�/��ԝ�(�����YyjEp VU�Œo7�#�ﱯ���s�f���.�O��/���^�S�0�]�������5�a����a5de��y�݌��i�c5E56��{U�{�Cݙ��!I�t{C�/:y�6#�~�n?�l�����/N_���::(��q`{Dl&�� �q"���N�3�Ϗ5�9� �0�˄
���T]���KK��Ҧ�fi!����l������v;��h*�+�R >o�A�����)_o5�;���2�]1��#f?�����^����_�L^{�js��֨�\��е�G�f���8��0�@�T���t��}��)�_��M���Q&�r�G��Gс_ή�!L��wF����H�	2<�g��c�G�$2��׎�&DB��p���R������iۓ�z7q�-���3×���.���R�C �O��RF E|>+�o=�=�'�Yv/���9v��`q�n��@��QQŖ�T�m1�C��+���ѷ?6	�kK9���j��U,MQ܃ep9���;��¾��y X㧳N�V�0Fj�K@��Ѫ�N�������W��ݼ|��H6iu��2:<޶�5������y�얘U�B����pH )�"2�O�]%��/��{���@����N��˰'Z���^�5�����!5`�X����U���pT��Gv6�i��lU('��7���8*2�iD���s���o�*N���%��E���F��dwQ�J��9��K��+j�&�ǥ�e�-�r;���>(�nb�%ik����>2ѣ,[e4���%�P |��a����m]�L���Aem_�@��A�����e��0�9Lי'��Ӧ�����	�/���}Մ�[}n�H_����l�;�5���b��W�0+��]���[텭I�L�#d����|Gc����J�h$� ��:�����^*��OO����V���+JS�C� J�ST@̱��ʌ� i�����G���]6�?�e�zt|<�k�k]8ೲ6SD��6;��]�"���}�#=J�e�c7�����?���מ�B��MF�� �}�<���4�G ڎ����I�/<ym�8�;�ec��jU���3�щ�����{8`*��P��B�N_B��yɉ�m��)C{���&V�A��^�*��Y�ef(�v��<��>��Z?t�Wy[�
�$	�o�����8�	:�$�?�����q�u�'HI���ă���=ˌ}�N�w�z�K�L#��5uː���~��^;M�٩��uu��:�CK�$_!��@\��e-a0��=�G��ݍ��U��p������Sf��L�V݅�Hw�%�fY�<��4��Ҵ��90����g����Z�M��7�	d=5ʴ���d���/��Ak8$�V�n�VFx��D��?�� �!3(�3�����"-���\��$�?��-���b�����'��� �T��Rw�kiC��Ϙ����l�6E��?u¬���	m��L�!��R�%"
����l@B��\L�u���T}D���i,7��]b�V�Ab���~��q�3\�M,�}癏��ɸ(�8�G��C���*�>:�Y�b�2h}{t�g�9~0�p�a�H�\�v>#�hj�F%�u����;�_��	� ��I�/R��hl�SP�S��w5�g�ŉyĜL�Y����k���6��u�݇�O7�W�L��ڽ�ļ�>�t�pXIz6G(3�鿟���ޕ�B�����k��1��ܓp[3��<%���8���7;X�Uq�����|����ϳQ�@���?e�����+�[a���1+���ht|(M���<��k�ZT�y�I���I۵���^���P�m)�J��5�����ȷz�߭�*T�)(ۍ�Z鸪Ĳ!b'I�a�F4<�T�a���J��d��P��w	HqI��n��(g���wd^��A������V�/2_Q&�%�@�Z��D�ƞ:"���x�5�E��F�Up*�z����(�%S�(������� ,iA�(�K&�zB{���`va�@����9t����2�	�^<T�Tt�[�d�o��$"���O�!�3���T�FP�T�h�Ev(1�8ڍ��A��UzV��u����m�u��֊�D�v��E����I����!V��d�Kiw�톮7P-��m�<y�J��t�QN�ћ�k���[5����|����d|}��I��Ԗ���.��Q�,:"���a��P
�I��t�2����XArz�	�/YB2~65)��KY��P�1�kf�o��s:�&[T���jȼ׵P�_W���.�����FZ�&*�����8y�N�]b}
q�䰇�6��lZ��6�g���TR�'�I���&�h���6�<s�Uᠵ�Ǫ-�������J_���%F��C=w�Q|�W5�w�v"!1�I#��l��j'!�z%T�:I���ıdV��|f����7^��s���<-�t�1��qޢ��=�-�cP�`[f]7{~�TOQ���-�5�l���w��;��6�_8L��L^��;�G��Kn�0Q��PD�+�D�~��i���0*R(~�I'�{D��̢m΃��mW��<�g+�x���B�
�����hٿrT[bf�q�\:}��eHZ�eLɓ�ޢ�I��%8�#�F�~��{���R�-��1�)4f�%�sR��z�B�eD�u�s��D����6�������bl�6��r������Y��Ug ��`ųKL�Ν��	&g�I�C ��T6��{�F�SL��?�fR�8PՄe�7tE��Bs4�	s�/�I-j�B����՛�ڞY���4�DI�]�ݨ�*�r�H�1�S������$��4���*yBa�d�R�ZT�9lx��N-[8�������J#:�gڜ�;@����ՠ�]^vj��k�hO�k��H�!5����Мealy�I?m��$��'a�{"������o�T|�.�\��Ɲ��<Y�@���s�V%n�v�q�q*��K��wٹJ6
�����.&�h�>�r�zU'$LAÔ��ߍ�:|3���Ƥ���{(�C]v��NO6ǡ��d=2�9�	�1��J�&;Y�!�Q���$�w��J��b�ٮ���R+fr��=���e�kT^��e(:,?�O�^n��}��F>��(�ϒ	� g��e+�4��Q�XB!�"�"��e�k�c�$rfx��#;E��:��p�I����+-[�^q�I�WW���YE1A��"�Zh�3��b4��>t�������5�� ̂�7_�a�3����6&zF�)��-���4��'����w��r�T�m�Ҩ/'�� �M��>����S���&n��ӊ�{��)v�S8����묝T sW���k����Ct�����b�E��9á���X����h��2�R�w�.��)��P1��a���E�io7�D�wV���Dx$�����sSE:��:߹0��sp�E��F���$����Q��)�ɶ��d�'����	��5���̬�� �7����`\,TA��
��;t@w���S��H8/�~�qiK�ef �0�3cɞ"�qr����\|�t�]hی=��g�����G8k�K�ʼ#id���KG��pX�I�8�6 ��d=ܱnY�0r��1�iJOES<~��A_�Tx������n�9�Q�M*��,�Ѕ�4?�ӾW֖mK�od�z�ӂHݥ��)�N经&ʲZ�?�ʯ���ӵ�SuY��Y�ҏV�34g͗��3&�u�5��=�,PC��.>S��j3�28�;�TA�]��t�����C���R[J�)���Z�VA�TY�b�Q��,��d�c�:�U0������H^U�XƱ`_h٩�-�Pgl딩�ͨ~��G6^�-�QG����ڼr�Ĉ+њ����S1���,�-�*Z)����@��ڃJJ E�nP�ptZ�~(���M��0%��w��T��fz����M���nѶt�G�r�@���PtM�#��ϻkzj=�i����������7at,!hx&4pO��W]y
o�e�}E�\��:�#�H�]�x�  �	������9�����d�u��"��޽ZMh��|�8u��t�R�P|�y[�D�_f$��1���P�c�&��SW�G`=@.7��?)����������s�Z���A�ZW�H_k�A)����;v���v
��v��J�Oc��{MT��z�י#Vc0�Vl:Q���V�7�2m�Z�w~d'�p�#/Ͼ�>������EC����e�27�����"�u�VN�}2��H�'��~~�ϊ�+��I�H#Z*�ȬH�tBb��{M������d��5 [������� �w�q]������/K�s_'%$:�8i*�\�1� 53�C�̥�Dhu��+
�]�D�ؿb���v�n���U�S��blX���F|9��y����2�l'AwXg /uZ�8���!pE��h�Na2J�c*��c)_Mdt���QCm[�ۗ�M9f�9)�jj�L�
z��X��S�̵BY!s�R�����E��m8F�s~��Y����ܒ��H�Q_ݻ0K�fp+�`˴"+&�Vlٓ�P"��9^Cg�Uҗ�(���(���iz0�c�2���Vam[=x�)��� �A�i��}@>
j��u�k�fHw����v�Q����59>�%:A+�?:āCo����U�<�L��<������4��I!M��"<��\t~����ٙ�j���'�6�f4��(�Y��y�/�J��y���E�r�BN�[r��S�Q-�t�=��~� R�����!�矪� �c<�/I�Xj��~5��?�1����Hs7s�b�c ��ӣր<, �<=�F�ZK�O��pa|��*�#�{�_h��le����|�|���=�Ԫ�H ����̝Ix�q�� ���V����]{�U�u|?�jV�pk5o���(S���՟�[_��e�G�֕��K�=�F��;S�׏�1�~>���{���u��V�	akG�΄�&���&QI�����s�%��d�5K ���{K�A����/y�1��u�r��������\Jl��Wq�@*�X{�F���1c�&vp�wL��V���(R����w�ׇ�X[�û�˓�=4
TT,PфB���W܆2wF�,-��A�0���eٮ�����k�(����һ����ȏ�oÿf�����ѓ�Sj'<����#G�?��fF
���Ѐ���k�|v�c,o��2��%����O;�~�_�EJB��3ٽ���ݽ�����_hnE�����<�pI��LⰲC�lav�]͚�~���~���&ᷩ�<"U�B���Ƥ�+��R�8�1o�N��`1x*C?�2�f5.�=4�e��A��SP%�h:K7�$��4~�%��chgAD,��4�AD��������yk���T����t��rJ�A�*CF�B��/��\���W�I�4Z��y��$b���;������rNɩ�(�q`_d��jG��
��9��a>@]���,p�1R�Ŋ�{�A�u�?�S��L*J��/aĻoc�@������QC`o�����M�M�}��&��X��&��D�wQd��'13�&�?+���B��VNt�q�������ua�%c"�G(zc� ���[k,����Д�B�ɑ?b]��T�)�Vs�6�ܗt�>��H1�9��1Κ4#Ql��;j[+��m��tL�I�t�a\��T9�~����4�!��p����&)�Dq�Jw�a�@�O��6Q��_@����Vη1O��4G�8�\]�i����A����c�4q�"f���m�}�x-�xA#5�Ñ�?��(ȋ�a3�ĩ�}v�?1�+"��RZ���V�D2�a���~w��N!�;}x	��m�s�ՄTz��3��~��� ݽ�%A�O�7IkG �cTv>3
��=W��e%��� �[�d�5�(�a�5�����˲�I������W�lb@yѾ�$�Շ�ۛ���MԬ�� �Vu$U���T^��K=6V`��Iy��]�f��3&��e�5�J��WUz�P��M�Bo�.��g&	�۰2SQ#z�W��(�t��3��ֳ��)!}�n_�&=��*m�iP�u� CG0�d|�洏xx�.3@q��[��Z�X6�n-�����s����y�^
C�h"m�"�$fj VUt}m�ܮ�r�i3�*Sښ?��9��A�NH��$B��OQ"�@7ۉ:�A|�<y�bk;��H`������������X��L:AV��� -��E��Xџ,��3�I�{(��J�����7/��� �d{5_�nW>W?饛�<�
1�sj�(r&r�U[���/ἕ4r;����7���0��Џ�Tn���d��!܀ư����G�J�dj��:��;�u�7��VG���I=�0�ۊ�T���'����t!tP��f���<�+�J��R$M	�J�;���&���7�q�� ������E�Jg����@	X>֗�(ŷ#�!	ڜ����?Q��9��Q�=��,)���(��fr;����(�C���?4���At�Th\�.���`���Ȃ�Z�Ϝ���_2A#�i�1�0�v���磶�@�Ks�~ 
@_�N� R�`n�}|?M����I���jR����`iw���Di���Ԗq=Cc��AU4ʝ�$������Wf�E%�o�̵�R�c>w�S�-\i�KX^`8�KTM��n"��zX�t�(�����C .�r}���59�z�N����BT\�>�L�A���_nĐU���� &f	3j����x�`�#^�X612fz��4�ݏXq���4�cmwh������b'�ћ����\*��i���9���\�~dPraOv �8�oDL��( b/������ޓ��[�?�s��Y{+2l�� �yݐ�M|�7����:G�V�w�2q��X�g�RSdSA���O�(и�{]� ����aI�"C�v1~tB%T�X�w�-s�9H�\�J  KQ����l�f�C��u}(I�i��f�A����:b�MaO�*� �����H�&5Lꆃվ�@�����J��-;�kv���S�f�_b�1gf��������-�͉K�R��h����ՖBk s�vp՝gz��@c��e�;�(
���.�H�F�E�;J���7�u+���[�Ԇw^����V�!vZ
�����pM2s1����N�5�B��(��C�%�b�������1Ū��SH2����ʘ���"%�_��Mf�fn����U%�%<ҠKU�_���>h���G��}��|CqI�/�%+��Fb�fF�F�p�v,��A�F���ܠ�P%,Y�\o�?��Ȧ� �=��_��cԬJ���$&%�m�65��bs5A� �G���MI_!���^�����E԰�mQ ����?_po���mrIR{�L /A@��(>�B+��-�Ff�˽;����K�j��&����/Ag��R�^���!�:�K�q�c������w���	E����Z,�޵������w(g�;���Ѥ��֞|�6F�٣� 3��e�-�d�H$5`
r��#~0��)�������1&����z�A����^)�T��������^�v�d�}�y��)��4M�%�$yP�y$;fn��gq�w��5ypr��U���ݎ��B�`+M��¶���D�	�ph�-� ��(,�
�]0� o�Pzm���W���zUֈ�/��9���"���X}�ϔ���1�ڴ��K��4���������R���pj�&T�fz}˻Ow\���ׄ omob:�.M����D����\c׉�� 0{��H_`I�2WM��ƌ�L�����F��.!�_c���0๑��^����kB�Y5���9T*�S'L�(3uTu��0����%����HQi���{����%@�l�؍	wP7�e�i��`7��G�
�x�@:�:�P��Jk��2���"�4��Ɵ�3/�1�(����=��E9V��� ��02�\�B��>9	��]�~���v9
��bc��[9>c� ��mG���`�+�Em��3DRȍ.q7O���j��yG�L�z_���6�Z��xa^�H�k|E7����K���٬*gEoAF��C�H�y�f��~��3M )�����F��H@Q�K�k��P����D���E��kxW <c�K[2�u��.��6]& �N�o�S(�	l���J�L��=e��U'�C%� �O�N�U�5�tnW�}�=V%�$���*��pa�q�q���讼��P Vrݎ��A,�xs�\�q]�?�`P�qh���f����_]#��%8�@y;�O>h(�<���fe��e |��@"ߏ�!�}�?��k����H^I#|a�p`)=�ʏ&���R������ΔP�����)��ٓ��q*��HU��d`k�$ ��K_��҂*^�'I��M
%?E��-�AB��j�5��%�w��Ԝ���`���l�>��v;���8qd�%��6Ut�r@�O���'��T�pXX��	Zq-�'d�ܺ�}�� �{�B���D��Eg��M�}�x����$�� �{�i:���������Ɋ|;)���r5K�7h��hZg��s�.��S���ψ���[Lg��D�ķ�J�*�Σ�ČǹA܌�L��r���璕�Ķ�������EM�o��>��7C�4N2���Լ�ܡ���}\��$ *,�2]1�|�pND�y4^_��8���-�3Z�ވ�U����[w{�{6)Ţ�����%��FБ֤����)���v/�N۽������^�vs^��qܳzy&!�n>9QjX����mҾƘ�W��YQ��$�b�.� �C��� ����]普�Z�U���KB8���Y�	�oalf
0��R��^��1?yQ?c��oO@2���z:��,��QiQx��Z䉪kj�7�}�H�"+�Nm(�s�|�W����qJ�a�{e�Gm-)�M�v���CG-xFYa3�"m5̠R��v�ȑ�E�� ��N�����J�LF�ߟAh���i��n�ӷ����Z#g���D����\P	����p�H�jjǱ���Fx�_�92z�陽t 5k `���.bߒ�W��"�ǽ���������6J��i�~讄��%�\��<.����3r�rCD�d�s�3rI�d�X�����գTwHpY3-��*LH�*f���/�1���qmh\�t1�z���f2�[�~���zƐ��:��a���Wt�v�	��I���i���Sd{�p������
��Ei5��>�֔�?��=�mG����`k
`�����D$e��TvA�>�'=����>�!�)f�K��
�aW�� �Qn���?���[����5o����9֭vw�{������'��{Cc�=���T�4�_a5��5.��ɨ��9��zR�&�+�Yn;$�H��Z���]��Ze^��Kz^�gX�|ơ}��Σ�
'3X��Q�u*=i	�+��M�܊`l���]�i�>��j7�8�8���뚽��}��+F��]�&?u4����G�a�8^�r���3��z87K$�晤���z ����txYt\B��9i�5+���C ǉ,{�J�_�nx}?��/o���'kWp�.�לi�P�f �'Iя"A��pٳ255�������a�����~�7��3�%aCE��%B��-�[m��U�;��
:>�M,��S��R�|�n���|��  �M5��%/9q�7�l��nq�A���x0��n��V�K{�����'�[u�X�DҋF���Mt��Ku���nK�Ӭ���(���B�b��ZL
�paj���(��$ȋ�^�7oT��Qa��L�OA�#ǭN���(�T)Z��;�	�Ԟ;�U
I�]kF���c���<C�K���]�aؠ�vɊN�	 Wmd�c�F���H�g�  ��.|qu?y�E�
̓=j-B�"����wJ|�R�H�)����nY���!DW�*�]�0��H�F���W���۩��� Ĳ޽	4I��UI;��aG����.�N��0~�ssw�Xނv�m�H�6Wύ�i�����#d+	��k�=�B��ٰ\����f	2m_�k��"ˡ�,�P������|��v����o�1m4�f����gl��b:��.΢,NI4�Uڝ��֥�I$��Q+�f�h��#�ٰ��k��n��2L(�A�.���6��D�HoVbPd��m���
�v���[;�`Ggb����ˮ��َ�O���(�j:����Kk1׊(����OӼ�Ԗ�Sh;��q��x<2�ķ`_M����K1U�j��q�q\�nBH��9�D�y�o
�0W������Z�̦�^%��J�L�Wp��ѭ��)6������\G��T��䩱��7#�oR������M����`Qg�f���z��fG�3G���k2����$��l�@��a���e�G� �싼&�3�M+��i�!-�L��	��:2��G|��i�!�|"�-gP�['+D\Ht}�<=�,>�$�TĔk(-{7}Y�ݹ:��Ĕ�C�W@ �Gsr�8��(�r�q�(�2Z���/׏n��k�UѬ��t.��W�-�H�;C��0����8��zv�^�F���<'�4�W\�a�i��@�D@R�a�im���
���\.�=V��k�_���+��2=�%k�\��������� @�NUu3���MB�Q��z�`����n>�v�UK��|�F��q�����&!2H0��PJ̟�֩�>Z��"ʂ0�ii������J�r���5NĢ�AU�<�W��o���OE:�/�o|����~�+��|����2���I��B9��:Z9��䓰O'gX�'�v�ep�%�N�,��H��ħ��A��&.r�Ւ��!d�S!�Ӫ�3�ϑ�=�}�^#��ib����^?0.φ	^PSUa�;x�+���h���Fc\!W�%��+KH�0�����Y�������q�[�=J�R��ѐ�R%~9�vAXKl�����֠��z�@4F7����C�SA�KF*�:�I�V_t�8���>�r��T�5|vb"OX�s�bL/�(��|[�x�
�L�!�蘑H@�.�$������P8L�T?ذ)8"ǔ�����[59�,$�Vw�֒{s�R�,(��Ќ�U��Y��L����d��V$v�xA�'��kg��<,��Ͳ�	�W k%j��Y��x��ָ����Q����l��/���~��10�ڊ�tN�Xyi�4�_�c�b��ys�;855���@�A�\�ĆK�ǂ�R=����58f+�~�-��mK�����*Jfy�ʦ��p�q*f>��/�FYרi�#b[G.�o���#��&M���Hj�ǜΣ�rb�r����@�b�ұQXj��R0�2��Z#��K�Q��p�I��T .��@�:!5�D˾�ܢ��<Jo?
��&��&����
���@��_�-e�JRp9q�ʡ]#'��m���u}Ò��k�Mr^vu�*��9��
���?Q�A#ZC2Z�m�
h�<���>me�� �.�X�w(�vd�?�l���%���/�zn���/��ʬz
��*\���غp���ɡ�����p5��"���CFQ��鯳Xm��@r&�0?�Y^j�|٤ݾj���2/(S�}���U�K� n��`=6?.�e�Uf���9��5�viQ}##NH;~>9����Pt��#�ç�*�],��,˜?�ĔI�h��_�x���*��՟�e���r�.��f�S��	Fe
ْ��Ik\N�̷�{G�"�.�Mj	L�W�G�G��gO�nLU޴cg�~���Y-� q�)M���\����w|�9�!���(�.&�L3�>�.��͝�7��cͬA�i��{���0�Fn����h��X����t���L9��}��X(��Ue�mG( ��re9��4o%g��W<�e�	�(��Ԙ�?�n#��I�t2+�1�B�����1y<�� B�Z�N��r�2�k���#H��N�-.N����ɽL!'����
���DRK�/���T-34�#�H��������/(w�D`Kΰ��+�|�h��ש��"�3���S%��Z�ΰpS���>��&ٜ�Q��5dq�P�"H�yՖ������Z��^?o6p �)�B86W[�ިBa���&ί��u�X�3\5t|��W�:�CVH�VNA��?I��r'�aUO.��be1T��!�-ٝ�"03��7I�;	���`c7}�
1���M�X��Ri!�c��6B�0�ŊOm����_�Y&=#�\Z0�����q7PKB&5��<Y	��U,f�T�~\0i�l"M&��k��h�H���Z�d������s �M,m0�4�Y>",G�x�M�=�`q+��,Tu���D��04��h��Ǥ�{��Ҽ:���[̸���pm�[�9��yY�����/��ǥ�� Pp[>���f�$-.��o���N%�B�v/7٧Σb��%�=7w/@�?��fX�$Fk�B~�ds3�k���wY{������&F)��ϴI+�7l�ס,?�b�~jl�����2����V8�	0��o�e�NbC�i�7�x 끅VN�7���#���K9!�V��N=Vg��!��SBtP�~�@�Z��-�*u�W��=��[2
ss�:O���|�3Ǧ�r6��%��s_=�-a�|����q�c)9쨔�簏L��}��~H����صp�E'��K�D�8Pgi���l�����?�+]�?_f�q�T#�����ʮ3bF��u*�V4S�V�i�X�Ľ���}.o�?�Y�?�<�T�`�6
|�x.�����atY��"�J&�
�����������.��t(96��7P�S���=%KBR�On+�4��h�M�!�Q�����_��#��F̭����m7��)5�� E	�?��_GY�B=��
d�=��pK�Z�x5wi5VI7o�+���\�f��y�[��DYRu��4Dy�i���i�X����H���+
^�u<\ԟ�����H:p
;�P���H�ҭ\���P�wf�ӟ��rl���Mt��͚�jYOp���\�7V:��yD%�g�X\�ށh�-_m��-��	��e*�-��h3V��ᭋ[��l��ݏ��-7�vM�.�aY�	��0��q�p��l��s�	{,+U��*O�! EAOaСe�]�j�|4����W���p�s�KQ�[����K�I��GooB�qb��0}l���c�p�������?���(t�mmP��`�c�}nG��}b�ci���Uo-�_Z���c�3ȗ��_���4�<���ڮCyU,UD�E<8���jo)��	Ӫ��r����@�T�OL��#����ʉ- �����C`���޼�YV����6���R����T:�ug�ȶ�Lsm��Q���$]��i�~M������7 ���2#Vk�(�յ��U�r�SD����y��1�5$G79�F�)�Z��=���p� ֚*y078��?�V�Н՛���k"�ro�t�h����N�$X�J{XQ�l��2�7�f:����������2�aP�|\+3��gG,��p.��k��HqXJ�oV鬝C=����F(*����s �)��$Ҹ=U5��	|��f[N!F�B�y~KJ���U���[��iJS|]�ǎ�]*�opa��ՃW�4s���傋��w:t��e�6���ǣ�����T蠸d�Xɓ��)9�l��"pq䬗ʽ��� ��踣@��C�K���Nk� �H�ߜ��=Xh��v�m�͊] h@�(�o�Db�S-f3Z7ȫ�$���+\������\""m)�aoo^���HB�4(
F_ܞ���LV��(��ϩD5:V�ͣ��3gOn����+,�g[г�NĊҫ�x��n��x�˂=�����n|�`5
gP���3�bS/�`��)f�\j�Z�+���_�ƭ}Ä��2N����tu����[@�o���D��Cb��茒��Q����|�W{^
�b E���I�S�F7k������e!���}V�㈡�t������fV�����J����{��w?�`���ȶIۥ;3�vk��bx�礴��N)ճ.6�k,�����";������ND�F��$���瘸�7���><`Ӣ�x���sj��^�9�EI�W��m�:��H�:"k�kz��\Hs�G�d�%����Iԯ6��&�sfr�I�H����2I�p���p9:�F��w��`��r�I����B;c��ϛ��%C�BS���* �=�"C�d-^���L�aA����+H��y���zj��������O�ଭw>߫���25�.152��S�~f͉��,�@�2��n�6�4�w�t��mS�$�B3��uD�|��<܎Y���j�[/�B
��m`�;:_AZ4�'~��綜J
�L�����I�(�4A9
)�Fw��z�N��kGUU@J�Q���u�սTd�^}���Mŏ���j���t0��T棝y�SiN+�
�5B��ބ���md0�1I��UYyc�+�8��t�h-Dp��˿Y1��f�sy�X]� �7"dDz�X��O.����R�^;/��v5*{�$@��M.=�h۔A��F�M�_��1�6i���a&�e..^ܖ֚]U��v�]E�dr������ �P�1%�$ښFx����=�7b]�+6G�d���N@G� �U/�;�G�.fz
�p��H?�,�bra�m�T���*f�f#'j�?��a�9�T���q�'М����n�%L�E$�\ܚok�FȆ�B�h�/�$�5�yu��=Ց�˾6��~��@vaN��,Q����G���S�a��Wu:!i-]�3��l1;*	EeI��<����Em�F�ܸ�.��j�Ÿ"
|M�;R�L��"����Ġ���kg5_$��j���7��`��7���ѫĆl�Q(P�������p�w�<o�f*	I>'Ai_��P+�'r:�y��� �pI�������Ą����"�	4�z�H�x8�U�~��k}�6f[n��|=XAo���s� ����׭�?��q�[2�J5��E���q�.w���	^��Q����TJ�:B(ri$e��w��S�����,�>� :�[G�P�q����#q,��}�.\���������(T 5�d(�+ɋ���|ޞָaq�P��'�u��;7����z������̊j�A�*���H�'���y���N�t� ��#��%A�_\��s�ꎚN�C�	6���-`�;�a(uy\�>�����@h�2�.��ޣ0�i6oU�z�}朱������������
p����tb����X�V�+�3Ȅ��Y��u?�R<Ye��XU�[^Ǹ�Gw��=~|�����`M �Y~G JΦ#�L4�mcFhnE�Ί�����$ٲ3IXq�@�_1�����-x�������\T�h�nC,pԨaғ��5%$R�J�)Уш������i\������K!a��Ӓ��q�&8o��"���GP%)�>��D�n*����,�B�B�v��\�֐6yck-Ģ\�<����O��h>]ۃ�bG�����!�N�&�^��tRg��YO)}QV��\)wc�i?Ep,5�Ҩ�~wc'+3�s����4�M깅aq��v$~‏�۴�����v�wb��E�������p�Jg ��1z��+��Ar�iz��ʹB,���gB�k�o�a$)�Moy�Ĩr�@��P$v\�'I>�w�P�,�I�$��W�T�	[%s�R\�AUr�p�^ǉ��_�u$]gfHa(�{�٦8�&c�=]���g������^G$HGMY�{��M��G��w��<��6�R�n�[3N�W��A�#�������O���Y�P!��	�n��5j^����QS�@k*A������	RW�l�&�����>��%�@�!�\�2Py�ئ�+�8 �&/��-�!���| S��>�O�u�v��8�Y~O��;h����w%Ο������s��V*��=T	�	�u�y�g�1�:��c�,wi�7�'�z�H�i�딽S��ټh�?���їZ$��f�D���m ~Pi�e�w����  pX�>�9��V6�l�m�,��Va`x��A��K�`o��(�n��ewQ�rI��{��-���7�G0��"������P�-�I#�]� �f6�б�rwӍ���H��
M-���X-2��\
�ep��rP���S?���;7���(�\��y�%rY� 0q�B
�]��Al�E	�G�4=ZL]~4C�N{zۤ��vF�d�g�ߟ���K�dO��7�Py}�B�F��p.-m<�QB��l@��΀�3��#)e���p��F�����e5p����x*teحе�H�M�h�/�|l�.���,E�l;r/�?.���{����_��5�k-m5/K�f�����仩fG$]ܪt�u�3!���g�
B~�C�����s�SN��v.� ��͐��^u�9Su�"J�?�]:���+K��%{B��@�\r(4诞�}w�{�v0�Y�_ ����F�߼���~�6�_?��&\9z?�¶?��H�a��U!�Mv��g���N�*���$�>B�J��SK�[��6�I@�$q�zDB��.bj�Ϝڱ�,�R��PH*^AA.�eW �d�z���at�jSz�kQ����e��2:�ƞ�6�3��Y�!���U������|��ϥ�M	L�#�P
E����陷@\�(	���'X���K�U����g�1���<��Xs̓R��5��w�Z�?Q�BK�v����F���:d"�(�j
��뤃���4��	#Kq�Bγ�:�JR�_��H�/�����q���1 ��.0���2^�$
�aԕ���$}��smWL�H1"}ޅ�6�M�e����Vз���m�t���j>��"ID����SE�a�͗��|�c�Ԛb=Oq�dZ�ԃX�v�����)�7����m���׿�,��My����F��������֥z=��w)؋���Gqһ�$"x��¿��!�)J���-L��������%��I�p��S��5v��V[
��2EK��mأ]3G��Ah�%|�.���%&��`�昫Ʒ��%�֚�7�zp�hu��'��c���j���
��>�����!��܃0�d��Y�d���)���;��f�U�� _-���u���x ���rA)��J��@�Pw͜U��c��Ie�	6����v�����)�� ������T��d��ĸ$*��בdIT��yϳ`x��۫ږ�-����Q�:h���J�1��	h�(M<a��{�.��:�������VqlA��0v>��N����by�Jѫ��ґ�HY~'&,���J)3�S�|vrf\��6��� E'�!���<����&���4�����Nn�G�tۥ��v���n�kAjK�#t}}�D��5�5WerU�?�ߎ�G��VD.}�(�p�sblUE�/w��2�c�n� 3gBA��u���Vc�\�;���d�#��P���1;�<��*K�K�0v'Ŵ��Yt���S޷=Y5��zx���(Y	�٠����ٲ!�I���;gR���K��+�9
˷�3=��[?Ԏ�B;��P%���G>mv/@�=�33��f��v瘚�Ie'��w,�f���S�}�O����hR�cf���e�ԩ�ډ��9����\���lm����ɊX��J��#ԏ �Z��k�0�9�M5/�wL��7�	��}H��?jM7��l
��OޖJJ ��+���~?� լ]}��
�]nq��#5�~�YI�&�sn��#u�U�	L�n��J)%r����q�
`C�{mp�*F��,)'�Tډ�X�yԺS�Mf��>!�?)�����j�L���kC�v�&��<n�tW�4�M�<x�&M�4�)*�~�_Md\7ƾG�,�f��`Ty�8d����Br@y�V �P|��C��~���^�D�@P�i��t�1�<+>�7�(��BB/V �p�ذ���
p3i.w�w��)�f�_PBp����{"Ɏ �(,حB"��P��̝��V���9�h��pe 1{Y�6t��~!oI���y�ץ�~жR�PRT[OX��&��*�U7�;��/_^f��{b�Y@�;���V�EfG@��L�F[W��D�,�6�lC��z��,�i��L4~fvމ�OV/�Ҕ+U�� ���L�~���J�q��3x�	Eq� ���~>pTo�Ѣ�4[.�I�e˲ֹ㷋�A`G����hd��� FB^��yD|&P/��cD��M��4p����%0x�W�<�a,�Z��y0���ƨ��l@�t׫��!��Q�"�n'�e�	�m�����ɚ iUd�7;�c=����EsU�15��7
���ԓN�[�I��U����� ����?���r��a�d��0�k?緃� $*Ŵ��i�Ė�g�q]�%�<,M#��7J����H:j�אX�m�zBصu�W_��e��iT���+�g�<n(
��>!LrB~��2�(�Z�Ҭ�ۼ���������<�KjY:0���0�i���E ]%���2���9��q־��W|��S��bj��j��c�u{W�ě�g���_9釽'�)vX�X���:��5��YIkȷUBp�?*Ms|�� z_�x�=�Ĩ�i�0��_$��}]�Hhkj�.Bm]��}CÂvȚȒ��%�0�o3�W�4�jF�*��$��d8��@���z|6����\m	0>��#[�A�N�	�Y^�l���#��u!v��TZB:�������8�5���[�E�!�9�K���i��z�S?�"����ÝC��S�/RK�����In��:'�_���K僐��`Y��.��d-b�@g����'�y��<����)��װ�;�A����l|���=��M҇�K� ��I􂣗=�đ�߸~�x�͇�������"5��)�+4=�����B�xl&!���EVW����XI�rر;�iT���[�TØ���}�q�I��ؿ_b�ԃ��o}F&-��B=�>���iA����D��Q��A�K���e���l�V�+{_e�����4`ר�)�d�aXϮ�H�!,��\�ae�EDh�ۓ�? �b��I;Nq�u'�	��>�`��G�����5X�����}�a�n:�"����O�-!�A4a�x��Ď(�sk<���(��R���P9u�20��"A�kz������v�Z��G(,vmṜh@�-R'� q'.N!~u*�MY���(/5q��CݠKCk�E<��j�����vv��ɜ>�ڍ���ERY5�_i�"Z=�Q[���l���vj��p�IS�T@{�)xm�8?gl��f�7B;�o~{n�W�u�u�R=��0H�I]"���n�Dqx����`ݚ���J�0�J�����B���t����M��<y��T�ZKw@t��B�0��*���1I����Iے�A�?�1+�@:L�o7�`��\K���W�{��$�饢G8�	�ͅ�(��7�8�AV�O�c��%��>�-��lw�P$�����?����s�3�����jC �� }+�<|+����%�\J�3ԭ0SsgY̐�	!�ϊ���f�� B� u�&W7tr=n�F�(�Q����8��.��d q��Q=��!g|*��y��Q��a	����L>)u���3�{��e�F3���@D��G�D��߮q�7�\����4Y<)Zx�}%_�mz��i1 +[z���0��,�C=��4:NE��]*�0����whe����M�U;Q�ſ�&xi����E6�ɳ�P���cS�*�G�l��L;���3ZS�W%̖�-���HI�E'�[����$�e@$Dr�0zM?lZ������� �i�ي���P��}�z���:��$�q���2�.��2��.[�T͐.�V|�!5ZE�w;d)&��p���:�Uh�٥��8(~��	�T��X��̲��e�1�F��0��
}r>I�oT�[���n(M�ȶ���<�'���@@�:����t?}?3n��Y��:e��@�B��@��ѱ5tq�΢�e��ۼ�<��Y������%�O^�A�����&�鉰-�ֆB�-����ߢ"`�ᑵ��ɼ/R��,�a��Q+i��m\1��X����.,��t�~���̱�ك��"Y6!��c�n��O�J�H��b��t�c���-�����b\�V!'���'�6u�О�x� m���]�#`�C1�}���,' =g��:��	v�
�j �c\��1X���ˉ�fQ����;.��
�7c�1�+.@�ŗ��k���`1�����_��7��B�|0���� � �Q��ۘ٥�i���(� r�y�\�;U�����ï�o\���� WWN>,G�7h��c�b�F�G,��͉~�H���[��`����lkk/����/�|�X�/b�� �*
iJe>�yT�
yVSK�h\hn�	��7�H�55������f:,�����F2����[wp�x�z��0)�X@}�b<��ikjq?YY�{�%��w��&(2z ��2u+���(>���W���c5ݨ���{�a� c�1�h{f� lT`�Շh� �@;)�~����p���M-�]욕�����Lw�����a�-7XԱ�N�D48�Uk� �ó:e��0��x�E��a~E�q�'l�M��2��#@�Sc�>�}
Fr� /���y��aR΃�!pdQ3��ĺ����0$ ˭�F����5�h�R���������Y����é����W���C/�cʚ{C��I�:���+�A�g&4�O��t�:�r�0V��5x�� ��b���ֱ��Y�fբ|�K���!��^|�?�N��.��<��CE<�	@]|;���"�'h]14L8_T���Z��7W�'5���^�˫>�~5��v]�X.+E�)�x�ro��?���5�g"�����*$Mqjp~��K��-��M��5!�@<�j�5��m��"�H�2iI��Ո�Y��ꬎW�����{�+i9�=��/tj�o;W���4��lP;S��Z������F6n	����0z3vV��W4�W��i�N�&]��D�	�cB�qD�XP'S4���~�Q-2uԲR���Sw��Y�b%�Ÿ��C�sc	S�S���q�F"�\����bS��l}V=��'��q���u8�h���Ɏ�3��]�1��َ�|K�� �����
��/�v��ʽ`@�CR����OQ>�a������It�\�=`nm5B����~3�K	<�(����m�1�]�qpc�0����V�Z%�י�9���A��~wu%��*ǭ�A�}���U�}iO^ED�sKHJ�alY���̃j1; �>�j�����|��w3���d���*.|yV+U��|�cC����0̓�s/���+�/��ieT&cs�j�F2�#��.���L�'��<Vֶ��ޢv+�>F�M�Q��GE7J:t�D �octU ٶ(�_d�Y����H��sIMFZȴ��	r#���O�#FQ1��e�✴�":z_��c��,�e�q+8�t���cQ��ә�1�Y^B%�P@��e��j�6 ��QQv����W�mD�	 _Z�Y��E��A�cZ�[�G2/�:�9�7��"������	 ��!��vn0��΂2���v��-�e� ��G�?�+��t��c�����cy�-<J9v���*�5���81mVv]�Rn�^��nD`|s�݇mz�J�,Ǯ��Ll��EQ��RY�q�.���	�'I0v܅Д�$\~�pW�a�z ���y>M�gl4�>i�Λ>dK�oM�G;M/e�j�������GB$�;��8���Ƚ��Ec��o�tŭ��'�ʰh��6����Y��xL9�-O��4�q�aj�?İ��,�o�d��Y���DW��w�,�����G�2�����1gi~�1MW%�X3w�Ǡ^��W�bш�G3��y�2y�E���,އb|�.�4��]ʅ�/s#@}�/]�L�;� ��3n
l��H|�E���ōԶv֋?ј%�� �=��$�S}_�Q���X��=ɘ����Rxʰ�h��^p�:���]��#܌�oW��qΖ��1捋�{F��&�]�Ƈ�M��Xd�,� >�a��)�@���Z;�P��5�O�I=�$־}�
-��)�4,'������s���?�|n��}}Uw2�t�&��p�5�s.�����87�^T�H8�ȀTf��9�6�jk�f߉e\�"<y�*n�Ԉ e�Զk��O�9@pI���hNΥ����[`s�x$F.`m�P�&�$�wܕi��
�sܔ/���U��X��� �4��Ҝ��
�u��y�������5�u�[gSx�)�g�����o���B�����kه
#�09$��'b��enkĐ?�xr8�.'\����� l��~�<��F���x�F%��J�F��"p4B�a�%QAХ�gM�
A2�S����ۓ����L�� Ia%�)��hk��C�p&Y>M ����H,~ ����ͤ�0���z5Q��f�u�0h@ωo���DAb�P����ݝ`���w�|�$c���M�K�;��پrr'j��@��ֽ:<�_��,n�fC���e�H�pv㣠�Ɲ�w��z��\v��vXFq�j6ǌ��h`1Y�E�����^��uŨg�k�n�T����� Q9&���a����WSj�x~���~x����(� �N��RG�PȔ�-)�dN�� ������E�1�ƅ�Wǁ�+��OQ?�׿)�UC��P�ו��	�M4η��p���k���
��gͲC��B� _�R
>s��h��N�q��3�hl� �]'�������%{�t���<��s�߀~��y������޳$ ���@�o/*ATr���55(O�x�� K�f��3۬���W�6%JZV0��̟�,���
�&M�er��E2P���Y����B�p����$��W�	fܗ|���-IVZƽ1w6��Fԡ>v��-UOg�����Cڲ(T��E'���Gݴ��:��Z�tP��O~�L��.~(ڐ���@޾�Z�A�!M�s�Ջy40�#��^L�'���g%�|e҅��6ғa�c��5�~?�o�g),�@�/؀�M~��� v��$ff`	�	��io�(�����Q�MN�F8�8�;Ce�=��ۑ�j�裙2h�Y,է ��G�p��� �̸������f*���h7��9e@���� �m�V3������M�θ��.�M�5lA�1��?jC����M�-�hM��M���E�Հ�v�ߗ1�A@\K\�敮[�>�i�v��@эtp!�ؼO�W&���}�e���| ~���kM�$��~I�1J��+�dv�f���*�!s���ƈZ��S�����6՚�g��w0�d�294G��qkα���H܃����]��>���!9��a��Nq�mq��-�l���5�p���#A�g(�7˚?��N�P!��*.�r��d�X6':�1K���LW�H돺o;�XXŁl�� �Z�y/s��jEs�Av��Y��2�,��V��C\ �۲���	�l��vOb;��۸���Ynv��h�_�Δ%c�u�&�6�'��K1]�]�>Y�.ɼ��3�`H�Y��O��Q?4�bD�2��y/�';�§![;�"@`�rϏ����(4_����s�'��\�鳈cNtYՁ|ƎE'_.��n� ��&LBq5w_eƽ���CKf����y��Q�dJL��F��ȣ���IaO�J����`D�u
UD/��1����\��,�:HE�`�):�4�͋�#Da5���î+v���ƧRऎ~Y�3c�U���Wk#�p����|�7��_�>	��]n��>��88�iA�[Pj�A$͒`�(s`�6�Vg�=�w�Π(P$�?O�W��Y4,����!<�8B�w��j��vk�����K���:X�ގ����W��5�'J���������إ�q{DnkA�!���k�՞[�=�dH���95�U�?��2Q���ZSG"���r��av6�K͍Zx;�Ğ�������Z�Tj���|.��e�BJ�
�e�Q�+�:�@��3�Ғ�-.�c(VP<�& ������v�A�����+!��!�`�v8���9#�H��t�b>��oU֣�_���ۚ�% ��g�8��&c�~wlO4�iC`����(-IF��F:^w�# ����8��1{ �֔�����'f�	�	ݨ]4�:�]�������:��Uc�ނ>G����1�X���{F]{p4 _-v�N%k|k��Y�e�z*��ȧ�*����W+g
ߎ@�iU�M϶�F��eD�,�"���.��>RMl�Fy�K������<0m`�̌[{b' �]6��-k�֋ƒ����	��~�tƟ�R��X�����olp�8{��_ٟ�nkG7:Ж����ǅ� @�ig^�?��[ނ�W��������]
0S'��or�m0�C��4�ؖ3YCE�C��eK9���i�Ǡ�G:+�Z�1}�u擦f�!��+��R�5dzѬv�sRL�c$t����@��*�L��`$b/g(=°^�GRd��oK��1���
kz<�[��]��:o���b�s����2�g��{��7S��̌�K�/�褑��=��V�@��e����j�������>ȯ\�m�ޭ �P��9�n��d�D����3Vh��c��� ��a���)�B�ndĨO���4�;9������z����ܮ1�n�];�\�t����`�%'�0oO�����:���tA	oH"����5+�`�!���>Z�u7Gd�Y�!3���V(9l��H��፱�>L��>�Dk">\���ሥ�%�}p�
�2���.A\��?I�r��z��wJ@�|�B�o��@X�"�q�\�Tϩ�{�C�ԹW�0�aη�l�1u�}~�5Q��>��\�;�J3�b뚞�Kz�p�iIL)�Գ�;6�G�9m'7�h����UN��i�Q�BT˗?�r���|V��f��_�s�r�a�g!k[w9�<}�::/v������% �٭��Y��\b:|t�\�H�O��;��K(��N��Ae�&,�@}y���t���ytGvg������������.�Or��a
����^� *�Xo���M�o�¼��̷U��m�u0Z�ʮ`�Kd���U],��a}t=��B�`E\>�d~'�(�|�`)�+������]c厬>K���/�-���3$��Yo��#��7!����#|�H�W�Ԍ�>��S����p����XK_�ͧ5��ų��l�kx���i�4�"�5�`��Y�2��'���[���M���"&z�ݣ����l����;��Mw�hIB��ź j�᯸�.O�rP���R@y*���4:���!޽6��k�af��O�.׭�J���)�� 2��g��y���>e�G^ ���C��ʡ�*G��2���]���h�^$�w-�B	{\%�V3[�RJ/��Mg��2��2���oP��P([@��5�;[ј�8E�!��dC��72N�@�i@���30�bs����,Z^��π�w�u����Oh�3qzm��$a'\����o��C~J�g�F,�B/H��딷��� (�7��QOߩ�L�"rz�e��v�`;�߷9�f�<H7��^���Y��4L�5��E���,n�.K�K�aK��(2n)��P]�!%�ku�ʖt.ve��.�B��Z�\qJ�����<4W��&�pc��'Sv���	ۛ�rJ���BA��-ö֬��x� �PP��O�_�ྦྷB�퉐�.ݠ�Α/����#G��t������&�ʟ��"㼒�ؖ�1�W�,C�M��Z=�̯����'3�pTH��eeKO�@��j�48V�Q��^�@��zo�P5hÓt�����m�~`ϒX �:d��m�]>��ETr�R��d�W?[�N�S��p��U��T�Q�2�t�m�S%�_H�F�o�c{�$O"a�A�aC;N������z��\���x�ӏ�|�F)Q+�B^�I�����T*r7E��z��hw�C�^�N��S]1�K�Љ���{��v,���(Z�<�����J��v����b�N;���������ܴ,a&�t�MK.+Q���e�o@ҿ*m_��<���<2�3���s�F(��'������%$b���8
D)���z�'�\N����B�MY��Ndr�?�o��XS$��y��바d'`F���n���-}gc�qu��1���2k���?�ة'anC��Y���z0W\�rʞ �s�J�����SH�6Qk��a�;��C@t<M�y"F��yәB�(���9����B�����NW	�dҮ����Y��,�^�s騈3Pub�D�'V��_:���T�߬�4��s �QHC����t��x�.�}���&������A�J��kh�E��۲�(!t4���T��38��䏌��5��څ����`�GT9Jk�l8�1��~��s��T�\1�@�2b���+灺f��R�M|8`dW����]S�e�N.7��~)*�x2��Ug�ۛ+��(oϋ�R��.�q	��"��#wѭ��mM�ʬ��@�I  f��-�i&�X*���L���'��ʯ��j�mNv�] �I���a���;��@�U$� c����\���&7t�6ߕ��+%�����B��H��\�����b�J@����=���e٤�2�#�6%�*|����&���w��X.��	6�m/��'�9��0Lg�vݚi�<��$���9����FX�(�;����f�z0j$�*�C �mk&)�'��Pp'YV�q��ҩZ2�y�6۬��$�n
O*,z�v\T?̢��rٖL���K�=`:��G>ha�Kh��%	é�WWrM'�.��%N�0�TNq"r�32�TGܖ#a�=�\\�<;��=���z��W�x64�?g���t<2�>G��S��;a*��}�46� ~���&���f�}��C c��0���h�<Cg/�D�׿�2ItL/�䄫����|`�r>�10j�?+�|òV8��_�1B2���]y")�tAJX�%�_��6Hv�p�qV{�r�}m4"�r%�ꆦ��D�m��JrE֏.TX�пm��+������T��n+�����&����͕"�Ay��.���Y��5|�56ݝ�7�In}fG�D�_�$�m�����X�ӟ�`D�4\%�#�s����z��U�!㆗����3YVg�C-~�ȇ�A��a��ȣl��H����/|%zb�m!%�� �T�Q&YE��N���wH�$2!gO�i��մ�d�ָ��n�-W�\�f"���Q�+�|��> \��1p�3��aA���*�B��ʝ؁0wT�U=�lN����lLP�K{4�ٴi�4���}��h��]3�c�����;$�&���Y�n���� 6V0{64��	�
CR�����1T�SͰf��)�?m% ԅ%�`PL�!�k��{ʹ�U�He5~����?XjM�t[�?|*���z��&0�-�[��޽��<�D��&2DsP�(G�|G�!���m��6&ϟ����߼e��*݌('lw��ݯ<d�r����ba�n�謄�u���:jS"���4���a)<0f�������A��:"q6]�~�Ԧ��ܒ������vu3"}������5���ݹ@D��J�Ņ={���xd��^E.�	�3�(�����R=�J�^/K-����I��~(�W�m�/qj0}��
ah%~�Pd+�&Y~2&�z 3{�Q)�����,��ۆiP
.�7�kр�cj�����(F��E@�!�_�MH6�
�;���E;mR��p���xQNW��H�����K�8���-�N��Mtp3H�ߍ(V��%AU)�%�{�Y-,�ᖖ�)o<!\sfj��R���U�+\�䋋-����O�������/�˖H�D׻L�ʴI�m2b]�c[�D�̆~�g��*,����w�e��N���h
���u|-3{"�cz-�����>�	3*����	�~>��r��E��Z8�~:�oU��?�gE��bLE�*�q���"3l��&�v�����{bvu�&�9�[<U�^\w�Is�	�4d�I`l��8�d�őxBח.��ЛB|���Ov��;����n�	����D�4��a��nUin��C���I'��jX��a�~&�%�ω_}�b��/���a2C��r����ȴp�����/��\����{����,U���Q� ��o|
ȷj:�h�)߾k)��۲OT�d�d�y7�;՝�\צ�\[ù�+�SE�t"�;�WH��^+aIdTR��XǤy�* �֖T�v��)�6�Ue�jy�J��#n�9���(Y�|�Z@��ma���ҋ��>�/W����@�w{���f��ko��"��"F��J���$Ⴕ�dO�����K�X��Ց���f�?/��	K��zb���"�!:�W���+��R|&��ʦ���1��BO90n�O�G#4�R(�{�W޴��6M͎�/Ω��E=-5	���܋LOq�]4Y$s�9�[���~���|t���FM�~	E���wP� )�
��fڮ�Z�9}�|�X.㣬��k2J������?]Ay&�?���}��X6���(�_�0�=j�`������6Ѝ1� ��`���f��#�̈́%<�?a�XLr���B�ީ��Lc��Rx�����%�[�;A�L�	����^��1������?�v\��s;��K~��p���P"THw_�E�~j=˿��2�S
8ɘש�oH.C�@#���@-��D�8U�HR �K�[6(2�<�A5i���۸��(V	�h�9r��C��б�w"y�X< ��>,&��hG�i�J!�ckE����eWiv�����_��������`XG�e2��0ވZ��<�Q��Y~1�\3y��QD,�&�g`���aF�� ��k�T36*ũ�]��+�z>���R�e�����#���X��yл�O��B�,�6��Ub�!ަب���v<CB�c�ۦ�*��50�ip;�����l�H�S�ɑ�t6���;���0:��:t����AY�QfGA�<�#x��o0�Ks��gWJ��j�hK��\#��bv�յ"}�|�4��dL:Ņ������j#�h}+�I 3)RQ�3&�{�d�	~����˭dW"��N^�(*n��>|ʰ�Q{<�=����X~�%Fg��R1���s��j2���m�����2e��Zx�!����=Ck�AV�/M�D\TQ�s�,m;x�a��+6QO�ҷ�!X~t�!����HSC��Ǒ_�r� e��]�5�s�C�H\�M9:Ⱥ>��O��-��� D]_Z3[�����ȇu $���8����5&�{��m}�^?�����a�|��װ%��*�tz�,��^�(ݛ�#�Ԍr�ub��
��̆n���a
��i�k��"�B�ەO(Um��?��C���� ���K��B�y+��t�O�����M�_�G��u�cIޝ������~v�E~��|G%�p�ל&�^�m�>MIf����N��4	��k<��4ֻc�en�JBpԣ4H"�٢m�)o����Jo����'9�~�˘�����Y�F����Rշ~�^ԗ<�;�,鋋����_[/�~/t�/��G>�\�:D����Lo_��Zg8���nr�g����#I�Ƞ��:å|!_.�>#z�7�ɝP7�d#�5�1��O�翤FL���I��0�/]�>�a��H&��mSa ��[a�O@�m�b��ҩ��()�Bpۏ`UP�1�|Q�mAD���euj4�Imñ���p"⎨D�N&F�Â2��+��{8��'�R�ŷP��4e+��������n!jM�H�^^��;�r2jL<��=���T`F�9-�g�D�/5���x�z���l�����\�[��Єt��������k}���� mq�^�����Ы�y�i��i�d�O�1hm�-Od'�u��?�\�P�I3c�U�xgz���\���~� t��䚉-p|���{��!�s��=����$q��kZ��_T�Y"rqЗE"̀1OAղ�K+^1�y7�}pD+�kR=�5����[~��F~��[_M�L`�U�"'�]Zܟ� �����,��^�Τ�~m�����F��Vn�E��RR��?����_rK�H��~|c�����-N6�b�]g1��~��\��r6y��lc0(��P�P�"4�F���$Ѷ��UؖaV!\
��kğz��m�W��sR�x]c�.:j���@�~my��V�Ѷ=����P8�{X�i2b���\5`��۵�츶}z� ��2@�2;SAW��a��L�l(�*эb7[��[J��S��
A��(�������\uhص&}���|ԛ�����7��Y\iV�:��*�6~g����jxlO0�K�m�k@!o���CRڻQb��
F�gwP����ّF9���Mz��@g�y��`tw�Տ� ���^�6�0N�Bе��F�ɸgm�����iӸ:1u/��^����I~6&��bs����i@Mn��o-������CW���u7��A�f�~[��f����?�K+��'SKs�?TP��)�����C,�������8/����Nk��q�N�C�4�$�V�ӒTNPA-�*���-�4��{���)�����3hk�|�>���T�̹�$�f(��c�!�zP�Z�\����@_'���l	T��x�S�%)�L�O�"=�G���L�)%a��W���71G��7ސL�K>�n���E7����c5�y�j���`�DL��ukѝ�d�S��C&�����F:v�\{�_���sE]�=2��>pWڧ�_sH$���Rw��Wb�g�k�$4��{�Yހ���w9�$�![����4�;Q^�W`'�v��f���H���!�nX]cO��&*Gj�Z�}4���9��.��:N;��^jr@�DH�k��i� YA(�U_r�-v�����K+���a`8d�͕�l�6|]��+�O�4~1��:� ~{�e�6�4]e)(�c]u�݅n��W���ULP<ɦ0��KTC���QC};���ާ��	Y�r=��c��H�y��&�DF�=K����W9���" ;w�B�D]���ToH�?n����1����T5B֜����9��@��.0e�D߆�.�lQ�;�f%���v��{���*&g��֖��R[�d��^�`k3��UՇ�wC�3	�s2H��s���_�B��-�*�=�ט�-�+�o0�J�DZ<�|��\��7	D�rݭ�������x[�0�(� o�h�x�t�K��%��^L	\�,r�.C;n��2�� �dvEDev��nm<��	s
��ORErM+��?�K���X,ǥMeE3#���Rw�&?�
{�sRhK��s"�G��)����nS&&�Eו.4�i|�s���m��6
^�b��V!]+t�[)<
0�
?j@>V��3`�V O9�>����<�˕� �SX��`���F[�x��� CQ���?�%��5���q��tM}��:�!�y?��|�x7�,K�,=1���/���Wƶ�������i?4Y'r�!zM$}X���P�[0��)�YwK�<�Sf�V+������ۉB`闢/���2�>F��;�=N�u��M1��@�WG�*��;^=��M�r��W2r��x>��6ƙ6�iƹ�h"�p�zu���z:�`��퀨��r��L��-$�oFG_�W���D����՟c�,b�uA��WVj�Z�"H������ٴ��#�Ra�isdM���u&�Ԙ�y��|2v��fjs~ة!"m�B�ɰF>�#;B����Q\�/�k�I��mh��(�p2�ɒ��!�^KW
���1�x=�s�ú֯r��ټF��r;� �I!�[PmOw�Q��H�M�DF�����䓭�$�H���md�H�N-��T4]�Ȱͅ�6��-Q�����P�xb����6;�)��t�~�lli%�Ӳ+=���B�vp��i�Om+lE��\N.�
�����zH� �0�a���u��r\����۷vrLq,�#γ-"�N5�菛��y'�̅���އ>9e��Dzu����� �V��B �N�)�!qS��,������J"7�T^X�{l��跭0l�{�yk�^��b��}��;�L﫬���d��]����~�x�FŒ�C������/�%��I]j���Lb3t{�i?�]�FC��%	߁��9a�LS�˱�:;��h.������R��wk`h_w ��S>~x�f��tbjA�$��'
��=CǺ��;&m/M^E	a�7v�Ҍ��'��$�,`���v58f�u%��#�Gď��u_�@`�Z���:W�Z��oS�����2�}i�70Z �� ��J�7nX m8��D+W��XM(�J��?�c���hs�JM��^����V]y1� ���z��C��}�����=���Ӫ���^�m����rG���b�R�y�C&71��5M-6� (�����(�hy��A�N����C�.;��2��(�'8i�Y�m�4#�'Y��k��)r�����י	�D&����#�-(�FV[� ���p�`�D�������FJEiA�������0��L��'[������)ܪ��pxQws؛V����Z���!���yFP
�0di�5�8����>�v&��(ifRM�z���偑}��*���M��
�>��qD���}��cÖfr�<������X.q: ���I�ŋ�P�:6�����}��-\�E���D|�\q��|������+�4lO
��S�(���1�C ܖi�툊>M��:ܩ��~��c��B\��䙭���5���f��N�J�����q@��)!���靧`��T�SX*B�+�1�-x���!�E_�
��	�|q��N����"v�"K�C���� ��Et��`l��[P�/y2�:~EON!| ��]���`a� h�K�����B�ٗ�% �}����n��b��Ɣ��?-N��2�`��֗�| "z�_������̆�G����;��S헧�Bf���9v�/��s�C�`�MfHPp����6�¤Ȓ�z����u�t��z��l�YV�:g!�9u��<?�.t���?�9n	�h�F������y%�����!�(~C�$T�$E��2��QRN�.��H������̖��3:��!anP ~z�6o�5�(�֨+Z����ع`䓗�a@�:郮VQs
�k�h�l�Sd*[����֑�P�7I���6Ihc?��r��EW�I#��+e{�M��l���t�;���mY���6�����+g�\���-D�Q�tN���q� ���t<h�����pʥŴ�W�z�/n�}bt��К�]z5�&=�d܈�K�pu���r�$zm���讟���e-��"�f@咻��9���{f��B!�W��4��k���摭X�	�(I�U%U0L�B��.L���Er���"�"o�&ۮN��NKɐ_ �3�\w^7Q�P�e+��/wצ\�5�S�ߺ�w���E��y2M�wŀ5�
�8h����t���5��_IeF����o�ꄸ% Y�v�6u��	y�00��Ǉ!_x��� :p\pm�'Z�9^~���N4O��J{�M£�K�S�����4}o�x#�ר�µ�)`5�Q����"YuF������0k,Hd�C�Ζe����N��v�T';B7ʔ�d���\������j�/�Q���ff�0�<�� �H���l��Vi$%fK���A���9>b��X��q�\3[�k��]�[̛�3�S�nA-�9d_ɗ�́[/�W԰�G"���lx�h���I.�Tbt��E7�Q&L���#�~�|ْ�}1���{i�ѯ��p����Pt{PR5GBHA1T$�oS2���6��|���))d�'{{�Cn2��P+~$ܤ�l󪩪w���h���xmX���ɞ-|�CQ�Bx�}������뛃���Y*�r�i�;
�i0�B�ݤ�.\�YXG3�w�T>�W�:u��6��vg���(���s��D�A<���/����y�2B�%9ѽ��"��N$B�f.ߵ0���2�t0��������԰[��s��YC#]�J'R�8D��f��ar��.���C�sr��(�ԯa�\�2����R��xl�}uW��+=��T򋅀�s�d�S'��q����z��hݹDU�9dj��Wo2�x��K�R�=%NC�N�
U9��}_��N��fy�$KS���]6���<�l[���ѡs�̦]���0n'����yĘ�BS��#�DƟ�BL�>����'��誝�6m��E`�Z��?�L�\��_;x�]�*�Ť��Y��IY���ܳ�E�"��鏕<^G\�N�N#n�G[�p��=���a��G�*?Q����~�A��(�6�*:߅�
�F�F���F�f_�47�#:�6��v��=긌�K���gjrݰ)���x؄���m���
2a��dr�����K����}ϻfUAU<1��[ˁ���~�#��9Pa�.Z�O/�ǀb �wԊ=#f���n(�>~�џ� �xa�^-�W�$�p~�e�`3D��xcZN����U����٤3�W,��u�n�;	�,����=��F��i��vm;���@������Uk��Z^Xٶ":#��(+�EܝFA�PjͪQ��Kw�珠u.j��M�,��\��N��>��\�a��u��
���tp��<G6���H��x���?&$+����C/R;70}=D�L��{%��0d ��1mC(�����?��!��(v��1N�S�Rղ)3�ULԱX0h�,���5�ޯLtlb2w2�nwtZ���t�*��O��kH-(n�%Vc�[�1���_L�\�ɞ
��f�F�׏�g�Ù&^�(����>���ww�k��4��>F�t<	����W	���ݓU �������e�~��a�D�nIQ%����2���R}�e���A�y��IH��4z+)��i���=��`�Ȅ#և�w���?�u4�6��T�^f���]���'��0�,"Ȩ��Z�}�idl�|��q�,ޤ�a�֡{q�����zP7p�nõ
���r1��p�����5G�Úz�'ƀ��?��j�I�(�ѿ0|u�sH�nqu�(ZQТ�������?WZi^��W!���!3(Qr������e�0���Q?��\��V�bKdH���6@v��pZ��TݳJ��i�x��#Vku�����gI���\[+p^Y���A�(L��
����RB�ƚ��Jn�����1뗊���Xa�w���qzv?���/�
[JA5rg�h��w���U9۪_R���OQ�5� QK���8��8�60�"�a��|����zfܣ=�?�7�d�g�hMB�1Mp�n��m4�/��i��<�� Ll���,=�+�~��fPr��<H6���d��AN����x�,/s�Ȥ\�DhgMo�$c����BPHq���>�LƝ	�F'��`�n��~l��+��i������j��j�!)�)����R�`���\�B����?�8��5���V�k�㡚�/q�P��ϓ�f!�u����p�
��������6ġw\���o�{�������=��K� �b����3I�;���QBQ>�=��Kb� /��I��Ӧ�5��/J��C�pW�f���3-��[���	+r&´ع���Lv��)g���Y�yWDK���O��]e,�6��F�R��5Ɩ�� }^'��,3�P	�\��"ѣL�;pbTg!>�1�uB~2x���!�
�	��C�������/���u]
�9��-;#%�p�/ō��ر#�j3;��hUpF�����tn����&
�M�3����H�/7�ģa�qb^�=�����4>r9'IVv�O5�!g	��`��,�����)��B��,�YS���I<���$�F�<f(ؚY~��$�D��]���r6m�z�t?T�?�(�Ti6�O�?QT|�م3����=U�  0Ö2����&Ɓ>����N�
N0�s�o]�8��Eݳ�1^�Y�rc@,4:��GѬ��j�W�y�e,<t�
ý��Q��o�j˾�K)�A��}�m��!��-��U������3t��9�X�$m� 8�p���G�WI���0����$fC"o�M|���m4m��ϰ^�,��*����]S��L�9��gr��.Q��-��n�g��Y	�8����c�s��&��y�h�ӫ�޳����6ȶz�ݺ\Wr,eY�J1��NH�#=���Eσ���>�N�(�Dx��M�w)%r��`G��\�S��5���5��K�A<%
By����|�v���k�i��-mF]�gg4�G��Ȗ��3v�`n�j��Wzm��9u��Ċ�V� �f�����yi�yQ"���`�^�~XnC͢�(N�}n.^Nc�X�2%8sH�y{��arV��ٚ !a�Ӡ\�F7UӮ05� r&�����b��bǆV����M�h�����v�~�~	�^��J7�չˎ��޺��ϗK׫���i.��JqB۫V�@�z*�����JϷ������=�`���!�ku _�fi���1�L�U�T�㰾�-���U���i�_:����O�_�.��~Kchn�����W�k9��	t� �+����i@����;�D�����J�Β���!��O��ɴ��yț���G�7v��G >ovR�g�&���G�e�R>�f��]*��n�3�Zu^�׸O*�@�^���/�'|⼎��[�Ԓ�fx�J��᪎Y7��S|���8�3���s�(
����P]܇�g�
}ѣ��1Y�C�C����ٺW��X	T͒�L�$T�n�J�}����Ì�cU��o���^΃b/DE��Cm�"��t~�A�	�x���&��qN��U+G��$"����:H�󳀅���)ӡ���3��-' 8*`<w I�Z�Y��-�ɝ�|���b
����d��C���g�mL������W�[J
��vUwq��@�UX��l�K����64S�TN'���`ħ�D��U��"ҽ�'�)c�>��1jbΌFa%1*J~����k�z�&G�͈�%���~�ԆKş��L,O/��G[6�c�kc��X-?�V�6>1ʞO�HL0�=�< �Οx��jD�ҿ�	��H �Y�a�ɭۅm�R�";ꩽ`�ܻdjrD�@ŶL��]v�6G��[��b�!���.��ע���{",�z㑧&�1=oom��F�j6���m< ��TV�T�8��F'��BBֿB���)�f�z��%�|�4|ӝ@���'���&�hkWYvUd��J@���G\�m�dq��bK��g��!!��#�}�	Y�"�s 1��S���4��J�o<)�ʸ�a��B�ZyD��A�
���C�ފ��(��rSG	g�tIt��x�jj*{k�'
��D�]�\2\�Hkj� ����Ⱥ��v�Q�L�,��Cjw�q�;Y�fn��݇�?�, W�.�#+=�*�c/9��;����p��i��/�4��^��cۻkU�R��7Ŏ�i2�0k�Ul~�u���7��ۺ���k��^��O�[Jۼ=��N�v��q�]���U���i7[�2`l@�1�px��_~l��P��n`X�UCV`�&����,A��x6�0���6�я�S��	��@��o�H��e�&���*�\V�@ߑ���!�Z�DD��͓QÜӰa4�=ҙf�
;��*�B�;E=釳�|��H�h�3���7.���������z�A�"h�����|���.����[D���Z���U(H4Wǎ���X,�}yo7�1�Ժ���e�����\OX��E����ͱ�k�Y���瓑��	Q%b"_�4�(��igEwT��[7�b!�k]��wD����>��������Ǫr�<y 4`~�5p�R/���
cJN>��Za
�q���|��jv2��s_c7v MJ]�e��Bq�Oߘҫ`.���D��y�����7�b)}>���iF�P��&Ŏ���+ai9Tn&��@����>��Fƞ�pQ�O$� 	պ	)g���^L�D\Nm2�J�N�{�t)P$��a(K�'5�>��/�췏V�{a��dY���x�XH>���8&����t�Ot���L��N��b�S8X`<�����n���ψ�ߤ.n�;�t�����1,��$M�^ ]캦�I,]ypj��~��wf��ʡ4Xca6,j%&N�|�i'6���u�k�zB��9��.�m��8�_=&��y�2̍}�E]3p��2A�ᬎmt>"|%�oU[�"u4f�@FN���p`X����J�ʜt�ӧP��h��]+}�TP9j_�
��Fx���O�4�tWkC�'p��Yot&t4퐘�>�L��\َj���y-���p��p���9�("�=I�D
�������v@z=��0u��A�"�V����h9�g��[���pOJ����6A�Qġ)�2u�Z-�F�mr� w�����8.�͂�X�-v��8�^_O3�5�9���S������Eީ`�&��f���	T�R�MP�&<P��b�j_dQ�����3�!�l�1tj��>`0^������&lb70�E`~���x���K��bh���!���#��v?>�j�ƋeZ�]=zp�F<i��'�g�tɏ���bi���!��ٙq�ma�K�p]��
�T�e�
��ȫbZ�%=�R|w�%\�9ު~���	��A��ѹ[rwC�����z�~�onܽ�;�f}�E8��,ԁxE�(LV_�t���I��)+/6��N��6I7[��w��^�0 �:�7����O�{����Y}>��6�L�X=�"�~�FF;qw��?J�7��Ƞ�&,Prc՘�c��".��.�!N�t��T|��
;<o�� �,`r,�#�n�1�1�%NV+]�V���߃����?���P����$��W��Rs	;�tʭ�M�dq�F%�Q�}�82'�l ���@z�.a,�ԶdD�pf�q2���Œ)��7(-/:M���H�	�%���l�R�P����T��Z+�����2��5�`�l�i�ۘ��P�\D�-��>�E+��A�����;k��]��a�l)��(&̺X�T�U�R��8�K������_"~)������p�y�)���](�*�n���_#�B!P���}��Q%���)`��t����sn|�mG�f{?6�lyYr��f0(m���N���r4�Zo�m+���B�'��l�}7o�^(�;��O�Oa�x �����~gq�l�x"�';�����5lx�R��i��&��k��ɕrQ��7�GXE�X0��t�S�4Pr%5��X�Lg�:2&=)+���wB�[/�Z���
ɡ��c��m�EuKІ ���Eڰʹ������mD�>r��Ľ�C�Q!X�wbd��7���[�<t���-��&E���h�0E�h����8�ӌ]��)�o?!Ph,��	X���'��$.P-�/�'S��Yz�JmU�7bʩ����k���Ҧ8g�0�6��NA�.���8���:w�"��9��o��������alW�����uN��bEl�C�o��!?8�ǎ���X�; ָ/�#�����c����߃݆b���f�ο��//���I�;��G/\B-�<>������c��¦���*�s�z_���G<��E�v��D��)�,C"7������4�akc�o���e�g���Z2�δ����EO3a�j(iY�b�֍Y�#K�فT�7ƛ�&�C@k�@^�6�n8q�d��+��;����hύ��Gǐ^
�o�P�݊�ɇ�!����뎧]S�\ s���ܶc�^�	c^r����{7e&A�ة���N�3*�1'�]���T*���h��cX:P�}0|�7���K1�v-,U�6[�Z��g��� ���f��@|A�PBX�Z��z4	�<5C��X�wŤaFPu����T:=H󱀅�ݖQ	�%Sk��jor`��U��~J�g8ǁ6�!��9�3���*�<Č�{��`�.��V�B���F�0
��7l�[�G�	��GMx|C��:�O+�wvڞ^9��ldtqE�`!4����-�����K�If�"j
�?2�f�{}zĪW,a��x�Q��VZ&��!�)�"��> -��\�~��1��`Z
A��a�����AU�I��=p��P���(�(ȴ�̨���A�YN�2u�҂�+�8��dI�t�d��)��Xp}Xi�>��R̙�*!�@Hc/���3%|~m�4b�(�� 1l��w��b�.,�!H�����"���d�r5���(�a�y�5��D�1}E(�o���B1��Lz�LG<M���q��zL�/�*Xq�VBz7"Т�4�	/�]O�Br���HW1�>��M,|:�����S�ǈ�r[(�WƿTw��7}˼�8�Ngs��<e���ʂ�ʛ�����:�D���@L>��u��v�T%�U�V�$��������)�8;�"x���C�ɥ3�G���aEC+�q�uᰊ7�5B��Ѐ��0���Ie͊���c[��VPJR%˖V�h��A+`�W�>0?q2�ε��a�=L�>����	�P���饺��Rjt�C�]��|(��U��k�Krv���ᦾ��0�n.>�u��V}�=jr�2_�N�/٥����Z�u�W>�l ����R���0���F��u&Fs�6-�>u�U��u�Sl�  J�9`9tk��X�a�6��@�W�FX��m����}[Ç�/����5`�_?0�lHU?����~����k�JŒK�L��t���0�TG����bg<�o9�?�9��$eq�}����'<��lV��z85�<� ���{���&���r����z>�I�ɂV�a���-l�b4�|�b�2���CPm����h��̑>��U�Čö0�R.�G��q��k>T�L�I�N���ȋ�S/�!��Hl��B�S���4h`U��ܸ�gkԘ۲d�h[���e����UV��'��
w贜����7��9���GDe�U�ce\�>�)�P�I]�2X�XP�Qu�s��|)�+3{�5�`̌^�t�<Hg�Qs�z;���U��3�s��`�A����7�  E�D�RN�`~@#E
��&���;��x{J���>T;t(dqlLPK (��@�D[�u����%��|(��TX�L��Vz�a���	�פ�'.Ƕ�8CG�h�W���fFTmރ��j���k��5��
���z��d�SC����(d���1w�*�ɿ�8�������{�9)P-�wpۺy�`?X0��!���H���ez�S�+s���"`O�Qᰂ���"�I�k���F��?��(������Bj(W��U3^6e�I����+>DY�"��l�?���� �j�'�I.43�!��L�A�X�E��\V'P�sX=�:���R`/�����SL�Q�n��U�&=�(6ύ�= 8��9�_�.Z<w���.� }��j����롍*��B/��%�x��ϚjJ!�?eR��BG��C��}�4 �=�m�Y]���WWg�$��:Y`�TTe:����&���t	�q�H�sL����O�NAT p*�$�nu΁��OU�8�4%A�Ibn���-�A�[�Z�f/2���i�<��P�ր�@�t�%Z������x�5sz�6�/����jr�LNEu�d��!/׾��	��.���U�'��_IB�^&����J�.%�����^]
�)�N�3�ak7���ҏ���g�[ܹe���(�x�ґ/*���ئ)��w�,\x�1�ub��q�[�=�A�q�����(J�/$���n����)O����:|�i�W���_+H��e�`�&M�t�iSBA�nO�s�<sW]��֕����kc�L�ɤ̠�?�@�IqU���qO�8xl�U�˲��.���feĤ� ��Qc��lm=+00������H��'V�]>Q�e�6�H�}���Ik�H�?4
���.:�\��D#(��i+Q��}:�Qa��ennl�w�QY���(�O.%�}	�H#����νqr�/��RC��v��@q�3�ʅ0��4�H�Zѧ�4�(+��sO
�@�@�J՘����|c�[=O1m��y�bQ���H.t�̧�_m��![���T/�߻���-HJ�e���L0A3�9����I�Hc�mܼW�"Í�'�G?���&\�6�?�{`5�����<1MD������g�GI�tu����D=��#���YPة���w�GΡT4�/�+�2d�
�i�r�ߘ߄g��D��ZX�qTr+ye��O���Q����݂&�7�V�����"% �"���J�̀���sf%��03�7��!7���I;�T�Ћ�k�ڣ�c{X�|���.����%�76 k%�X��4��M��-�5��%}�8Ԫ��IlC�H�!�����x,���D�_�����2y�����="r������SX�*r���}�N�[W�/��1Xڏ�MmT�.`j��� i�E�Q�>.92��L��o�#�z��D�O� � ���!���g��^2�C�َ�w�
T�}o�R��B�(nn<`���6���8��^�m7I�=n�P�N�.���H��ָ� �Y��������	1�ӥ�ߋ���Xazy��:R t~8�e �}<4�[�x�)�<��jŵ2$��Su� rG��]$4,U&g��"P�<+�\R�ޏz�����
��jĲ6ɚ�z�V���6�FC�3z�?��c�d�z�Y��� �8*�yn43�񴀗m�Ǻ���xӆȊV���`�������=�ɤU����ca���p|�`K��&�L��[u���z��4�8��{�6�Y����R��Y����N���vgf�QC�������6fmN�D�ϥ����. � �)����� �0�BUj*}�!P�t����,�O߱"VP*n�++��t*�K��R"��1�ٟ"2h�d�7�;w��G���m:�'�G~�a��7�M=8�+�%��X�y�C[�AbK�_�[�YĲ��]�#w�P���!ݷ�d�B 7���hvcP8���;Pgje��u1�rL��j]А��`��=Z�b0��s���`�L>.xϱ��Ѝd9�n�M'u�F��0���z�z�2HQ.?`�}sL*Ȥ��=�c1���*�ٮet%";?r�"�6�B���m;��a)���f�g�;�#~����A�[�y�%�;6@��Z
���=?�G�~��b.T��@�:�g^�=3���z E�J�!��M���u�zƸ)QFi����s��g�;�0���B(:AgCZY'/!�Bog�f�Ղ�9}������u�wr�H�߭ڸ�ǛM����1�6��_�u�����o�OR؟���]�ּE8mQ�?�Iݲ�x�e-yY0hk=T;�oŮ�y>��fj���D���W�*"�ٚ�T�ۑ���z�;��9���7\'Ǉ��v��J��z(��EO jh��u���4����U��X(��a����5���{G�-�-���F��+�60kOmj�5����1G��dM��=��G�6:�T�^�`N��𛷢����w����zd/�{Qy5�*�r�/XV��y&�dm�9̬���eǍ���i��	iX��ą�hi�tP<�f��҂@�C�p��Z�)�����Ճ+j[��	��~�o��qp��ٙ�G���l�X&�%��n�T>>������� ��U`�d]�& -;T]�UY"=�6f_�N1G�z]>�9�^L�:�~o���'���C��n�ڈ�CZ��ԛlk�;籀z�҇�_���λW��1���Rx�u[cc+ŵD��D��d|�K�cP4`t�!-��Ůs] ztU�x}]#�2 W����y���אt�+����y��Y&m�^���1Md�)z�'�z0�p��s<k�C�|_5������LS�.��Э�S����؁���^��q6훖�6��mܭ>冈����r�,��ל����T�۸��h�tzVtD8NC��I��ZfU�;F�j��Z%�?o.c
�A^G\GT:n"�^9v���R�H�LM%K����\ӧ��j�:8�R4���Q���g�s�U����%}�E��> ��e=;�"}� ��w�z���ԫ�p�K�7^�*dp��&�
��c'��(��@�	ٷG�!��痁��{_����
�����3z�}�j���(�y�LS��\']=_�>���/E�R{�l��������.oY��O�(Tz,#k`�,G�HhPr7.�/\�\#�uG��o��\`��S�qk+�+�]Աq�P\��`f"[޳с�g+�C���ߴ�:�e^���۸s�,�	(k70$�_H�/eu`�	Au�|�M����bp8��!�6J�9u�7Z�Y
�� 80�Ny���|��z<���\'3���7�?��i���gǐy��_�?6Z�t;<+_]���D0�B�$�/�^�\f����j�෇Oo�*/�X���g5���^~��<��I{�5����"z_Us�_�!�jZ�V9��*�s�� I��e����|�s
[~��Kܫl�
��T6���ibqf�`S��v����������^��ݽ�?�$?xf���͟g*"�"�D~�V�#��(�i�y�F����ې����Pf��{�B*�EC���Ն�m�6�<��R�������ߡ��f�?6h��O�k�c�h�)��g�5�ر�)!�$'��E]X��%�����æ)H�����F7T�g�§g�����I�_�:���n�K�^�dY��n� Ê����d�����V���ܕ2��N=�(?3����U�'F<\l�/��(�bh^�H�x�{��k�a�z������Uw��`�w�Y��(NCۻޗ�A�:,H��@~v|��ӃQ�0���WK@�c�E�Y-0�Ƽvv�u>(Uj^�ߟot
K��<O=��k��]����d���%�j4	�b�*E[m����!2���d�0�q(6�����wO��TrD��EI�kN{�uf��N�V;�o���h�~+��n��m����ڸùE]�sd���-�hP�U]���*�v�-m���-����m��mڦ���)�G������bݛċ���@V[��=�R�'�THJ7R�ͺL6�%�E�YZ���_���Bѡ�5���IsLmh]}m�#�{v�FH� &�凅�� ����/��%�i/(<0/&$�A�N�D����^�M����1E�&�\���-=T}h���.��4�����J^F6��	�dO��f��ꠓ��ɃB���4���em~W(�S�dx��+(�y�f���+��q�VļCy���i%�'!:�uO��C��s��X�rM�#�&���|mQ���ğ �rPoC|G��֪bH[Ih�eڝ��v��W�\l��H��9'rib�!�{�I��2i�6�C�,�j�/0y~�5�A����K�vJ$���ɧ���q�pl���Pa�M*�}U�Bw8���Q)��^��I&!B�zĥd�+"�r}ǔ�����e�S‗��>�  	���؎R/��o�Y}3������bI��_4�$��6;�w��0�l�4��,�E�*<���VS��K�a�k70� �Q����1L�� �� �c��VE���8����`�.t��i~��V�"�d��iH����"g�jKF��4)o����1E�q�x��ZѴ�Beq.-¼;/��^�?]�WP�i��g㖥\v[��.���4���(��v��QF�k�b��ɦ]5�c�ѵA �c�J�����qj�]e]"L�0��`,
o�@I7deMoд]],��D2G�m"7�Unn�f^�Oulm���3�Oۿ��-�ow��$epO�ca+$O��-��i&�<d�=��pW��c-�d^�r2%�����[R��Н#��U]l`k�vj�=�#�k�#����n1��S!�
A�M4�.l�ȣn�u#�:�*�Qč\�%���|9^��-�.�drڠ9��,BO��"�9�32A�p�Q���cAvs,_Cs�R�
Ӱ�M���{e��l;��� 8T6��'�~���N��
I�R9jl ��#��_�o<�FbWO,ĩ0���/F�&���ԇ���\>��lȾ�D����J"�Fa���Y�U8?��2�P6S~
�>a���!�7�X\/d	m`��BM������e5N�F�&Փ��-�1��87&e��k/~!�tH���`a*}�Òg=���8p��鯧�n�,t���3 � }��S��T^�÷��k0w���Mk���/��rs�rý�m�~rJ�(1w�	�.��A��3e	5�e����i ��FD���H��Zd��ԓ���w:"`d�ĖW�ކ����'��ɁR�FLިc��x1�
���}��2=ɿ	Gp�Vt����bW1G�ؙ��NXm�r�,�D���9�`���{�w=4`��0 ��F�h`�^L.|�z74��}��Q O���G�'�'�| 
�{�V�!���d'�s4��?�#¹�L�b�u/����ej�ޣԎ�?z0�˴�U���ƙ����<ؤA�CVV�+�`�l"HW����N�dB�m��W~D;&Ho��Ja��Z�$~��#b����p�Bi,͟�.�R��)2�͋�������!rf>�E����*:�'�ft��݅��k�՘��ގ��*@Dx	���C��qd�(Aފ>�k��d/O*�[@�ZOC�h0��<��ʔ]�*�C���Pp�
��9X��j����T�^���^|I�bD
z�y�5��6�fУ���~�aV��CK�MI,|�����oU��=UPyg�U�v�,�*�a�bM�����-�5��G���Ⴗ�m�l��H����۫�� ٧��CbS�P��q�
�y	ڟ4�)t���U@%�������p�����؎�8�b5r;2��F|F�w^6=�.c�����*TL�GF��5疱j�s��Y����0}SF�(o��g�����d��jI뽩"7~��ۿPT�&�%�q��̐|E��z���ꂧi�H�/���[�&
��y�{��6�:R� ����Y�-�����?��$WC5�PS�*K���?���Όd�x��䊹�t)q{uU'����m�w
��hHĆ���֛��I��up#�[��;�=�q9��Ođ�NNH��:���>��o^npN���A�!�����4�vT
��d(˲��y��c�\�R�G`�j�m�;�����[J$Eۗ�r�V��4�Q�����ؾ;X��f�OI)?�U���~/H�K/�͢ '��k^eϡ��H���lwk�y�*$��m%H(!�6)g����ˁCG�&3F��a��e��ٰ�1C{��6^�f� ���~���;3�5CJ�h,��+�T��HѐPFp�
!��5��yy�� �����Z�����b��Y�d� �
�I-E)˷��4U�p͉� ��H.��lL��pЃb��q�{�i�Vp�̒o]��/q���s4:��P*��"�r��	�Y�1䘁�z���?��}����0^lK��^�bǙ>yl/YQ�?��NǛ�Y�'tw�I�F�ʺ�E;)�)�v��~��\��N�@�2�?[��P���1�3�J��	3�%k�m��` �'o?p�Z�Ȝ/E2m*
��3Y*��%9�ohH�>K�è�Y]��`р�����f>#�T�`FQu瘆���c�����>C���r��dQ�����MgS4eQ/����ɟ�z��=as�ă<� ]s ����YB�9��/28T��Ԉ��T�x6$-u'�=��]���]T���ՙY��~���7�%�3���S���?�Xc�EK�-;L�[�0���5+>z.Wq¨<��/iGJJa���c:#9
�߉;}4��&����5��E�1����a�*�0�"�����&)��L���tOZ4V���Ҧ�!rp�(H�XO�?q�����Ue����Ѐl{{�e�5�e�$�S�h*T��y�;76l˂�Ze��i50�G��aq�J�f�Cz���,���X��I@�M$f��;��79�kx�g�+�S�#۱�2^G�r{�
 c�=����H��ϵ%�%:ؼ��S�X���S�QB:�4en:gی/7v����ݕ�E�_`l���͏�2\���;oV�}�E�+df g�R�1֍�=86��@1wG
��{	O2�]�w�E�N��p��U�k�{ �d����1����Þ��Tk� <��|�g���.��	�W�4�����>1m/��Q<ws�ZRS���q�+ٶ��_�F�ߍ3��m���dA7�/�
'�l��W��շ��ԫ4ZL��Vx]F0���0�}c���º>s���kf����`�]ޤ��H�����}�,$�g-ߢh��7**�,'h�`��y��P>v��Y���p���u|ʉF��\LX��8V���q�yH ihGX����aoI��ptWRT_��J$��6򤅅�\�Pny l�tyް��� ���j�V�ՠן��)��֣����@O^|�����#�����i_�$�DQ�.8U�4�L7頫�~��EtG��~�q֤��27JQ�@F\��GTk�77�,�MXt<_��:��+�쬳�C��-����~���xF��Z�=p���U&ʾ���=V� ����
`��<�{���B1y�XS��(�|��fF�F��|\�F+�W�q������ˬN0vy���D���M�8fN��t��AO�	�����q�
2�͆����{	<�8��R�O�d�AƄ`���a��\~�}N9a��t��p'���u�l�\���&�	0-�����?��0�����c�E!<�-B��v,��j��z7=�p'P�����+�#��΁9����3K�%�I���c>��68��ě�MA�)�������"���	����{��U�y�����-�
	�/@����B���#Z�Zt�yO;1kb�GI$ƞ͟Srj�4yTG�W1ѯ}�?S��*:�~����v�:��Gŗ5)>E��\�E>;�髷� �"Ne�]�C�����d�k���^4Ȼї(�l� �{���[eɝ�4c�E�i�Un���������tB���,Gz֕!qYr����xo�ز��&�V�T��X�#ęM��%�u+m-�3�h\]���^���w�[?�W������̤�c~�r�Sk�����#V�uBH�wx��ױ[Q���ț@Gޓ�����˃#�M^�L��� ÀT3ntr����ӑ6�%@jKy�@u���E<Q&o"bl�ʘ�Ҳ
8�#=':�vܱXa=��!K�㸊�]K�{G4M�G�#倒(=�����W�����ͧ�<��jN.l3X�]@��1�i�Z	��[4������H��B�ĔZ�x��H̸�zri����]@j�*��*�p�kYR�0�>������H���s�|�Q+4�G�%}>��I]?�1=M1W�N�}ܥ�Ii�~�K�oя,�y;9y^ ��C��薶����|��&�?���D�?@Ak �լ����1��6p����d�w��yP7B��z�c��;i��1ʸ���3~G)��D-ɦS�� �H��4��{�(j���V���Nz���~pٵ��,��%O�yX�h`�F��8K+(n_��B�Ŀ\
U7�ӳs�,�1t/d�ħW�F�Ƈ����ٺ���m�r�:��Z�F��5P��L��-�9FM��J��Ͻ8�e
��P*������f�S�~t�
첕 Z����!��s#o(C�Z.;�%M'��;���V�7jT�e*��Ә�����;�q�_z����T(ct\�Ҷe��쉨5 �=o�(L%�8dm_�Q�k� �S�`vU_yx���__ �y�6�
�*[�[fQI�(\� �n���5������'���Fũ%�dǂ�ل�P�)寝������p�I���p-u����F�y�A��� ��Z7itpʷL���$ʂ�m፨�E���~08#c�t�h´���mp�D�'"��7����o)���E޼�	�׻W_���n�
��GY��j%$o���g��e�B�1�6��v�v9;����̻W�2V� 5�sO(�Q�=�.�y�$�5�i�l�*��P�u��GX`nV�^��m	F��(����Õ	^B��A% ����A��r�n�0f͡i1;7{�|Z�׎��J=s.ᮂ��fTh�T5�/����"�&S��m���Q�6�;?� Fc��`uu�P�7{B�7	sH%�j��w*�*W��0e�����Wc:5��c<���8�*�=�0�o;m2�Z�%9BP���	����4n�'9��g�>�Z��}��'��Q�h'f�6),	�����\����7������9����]�O�P��Թ�PftV�8� ��F<'����1�����E�ap�3 K0w�s�貚�'�|LJ@�B+T!�Y���]��)b�+� C�Ma��"�o����A�b��hB�6]�cv�zPh�}n���]0�`Q��w,���K��kI�I(7$5N�8��76�N��+8|�|5~O)�O��t��.w��Ƙv�/�q�� 1~��Sh����}.f8��A����j�i��E`�*���T"��\L�@�[:�����v���tߞm�\\�f�{�mR����I��W=��4魋�ۨ��Pc��ѝ�~�D�N�ۢ�2�'��\a���m���d�)F��@�22OD��!�s�"�s��y�>��1h���FEO.��H��J�!�v�\XU��@R�7,:zE(y��BJ�-�ew9���}�ʇ"S�7�):�@���JԨJ���WĮx B`�	�]��S�S���Ct��|�D���K��%�y��%zS��{-Ӑ�F�B9n4峕Ä��9��DL7۴wȠ�NiJ^�ո�g*�Ʋ{G�RqL	���W ��m���$�Y��.j�i���\�JQ\�f���TMOϥ�ض��L����z-6���F�Qs���Y���F��W��qk���N&W?�A���n���5�`�hN�c��`�
���7h����d���N�81��S)�F`������k�`�崗M���cY�|�?|�G7����R&0fn뮋�,A�Æ>����W
�m4��b�A��{�lrg�#��*�2������[�#N�6�ӥ�*�����@����oy���@OhUƓj��w�_�_+��FZ+;�z��p��h�xL��e��r�4?Q��WʹJ��s�Ӆ���PȋЈ����8r���H�qؒrη�Ү�a�̮>��Z>��=���N\���v�ӱ�$��AJ�H%�5�d� �̯S��V��⒩j��P����^Ι��/g�'PiF[㟋 ��B�[�2��uڴt�͊�(�Z�l�8[A��*T��)/W;�_C��B�
,� �*��cWIj��J2��`w���-�Bj7�ڊ�9�#��z=�(�sl�ېWM�e�NNB���p����D����c�^J	r��q�����ˬ�qwn�g�Ns;JoG������,�[����+ V'���@�N���(��}~�p�㦎��=�t�j�c�N�
�_^�v�JJ�mxK
�b�g	B���y�\z��*����<�:"�y3%��s�L��[9�������1�ǚ���li-�ҥj�a��/�yy�ra�#���ֿVl�l�a���.�a���iy�8�b�w˺�/Ĺ����A��ѮV��UI^@�o�����S���&Rn-f�d��'�V��|'�к)iC~@��:PB�r��r��~E���F���K "c���3eG)s|V|��K�ОDJ����h�^� �#;S�����Q�ߓFle��?ƼB�	��6������-1gJ�It�v�@$�ew���F#��o�Mjm�86
�r|�WP�̍��Vs�Hn<7����M�ԁ��;j}�n}�#��.��F����f=����Cl<��{�戤4d'm�a�<6f1ྚ;�����H���^�p��lkF[�Ϟv#�����Ps)~jh3�e���~p���wR٣QN�aш�=>缎ں0��n������]�����U7 vx��^Q��F�st�)2Y`���R�c�X�I�U�<!��`��r�Q�{���v�pX?Gq����X�,g@C��Y��m���0}G�]�e ;rU��ȼT:s�k��zI�����O����]��4��j�Bǟ�qI�H8=Z���}�n������`�sr�\6�p-m�/���z.)�зF�Eo�8���������m?+k=�,�2*�U��r��d/����4Vg���g��U՝Ih�R�T�.�{r����]�
¯zr�;��Y$��D�|D��uq��t���6_�@�4�4I�~�&���%([���{D��=v��{���#��^��#�!�e�Ũd��U��ܷۭ�������yƏ?�܄@�A�_^*������û�AToX��Nô�g�0M@�U˲�SbKmt�A>���(�!T��e}��5���.h'����~Ε�;����/�į�DD������]�j�M-�f~ҚqtT��d}�?�����*��z�2���|M'T�tJ+<t�AL<ѱ�t�U¶r�3��R�hM)p���I8��
�"ٜ3�����Er�)�+�;Y��r�˥l:�Xն�M6_ �c;4W��;�F}]3�f���c�cҷTLu���)�7�����W�pA�ċ?R�X��g��O�=��m'�����(�)��gT5�<���%i��ǟ㜁D��*uݦC�BZ�pD�s��)�kj���_h^/WVyZ6��c�m�N����fb��o]F�-���̀y��=ٿP8��.W5�s�4S�D�_�\J����X����H�ЊT`����������ce�0g��cŉ��y�G�!=x��ө� ������|���v��s���Ή���[�3�	@\��?c\*�
��6b�1�yȉ�&!&v,Q�P��'��$�5������Xf]�F�0-���)ozD�P����0j8�(�c�̳r��D��bl��S3��e���l�q9*?{#X���i��.�7���Jh� hN2LB{�z�F��C�N���ԛi���v����r�z.GcՕxa륬7�FN�x�D�V�u����������"5�P����*�沥���r�^C*�����nU�{���p����Ӹ넹z1�s�v5Յvj��'L�?���Y���Y��Bz"��L`��n����i��5�r}�`ƹ9���GāP���e$�MW ɇ�D�����w_��2�_Q��~�	��/7��#ת|���*�筰sW����>�G��4!��k�^?���u+�I�*��D��n�
B������L�`��\�<.���:R��	/q���d�Mi�7B�ao�_q�L���\G[L��ξY&�y�������Z띕|��4�P���$k�C��$�N>_^z���C�O6�=�V�L��!g�,&3���S���
�^`1��7mL�d���'Y�Qڏ�>l4�;\��{u��j1�'��ƣv�48M&Y�ׂ���l�G+P���{mm(9j�}cW�v~�t���V�KIE�?z��
��h������,��U�'���P�o	1Gd��2�e�0�����C�D7]�}n,�@�yI�:8�_����~~'+���1A���� �az��e#]ޮt'T5K��"�L���������J1g�b�=Q��%8�;����=�w�l����:�R�0�e��q���>Z�����ipU߽t��dQ|��7��9�AM�
����j�rL����#��U�M�P}vD�y��B�P*�s&~����:[��Wį�������,�dMF7O���$������3Y"w�?
U�I<mD���|�(���c=��"�������������2�m47�L�����9��b�����:��B�;����ӝ0w�2�S���~4��{[�ZQ5��]#�]c�Ֆ�2����f���"�8D*�C�5?����v����Lz�X&�N���������2�76�!��avP��_1������:�x4�?��#�K�bl}���(�
L�4��8���*�(}�K8��<��X�U+�;,����Br��9�v&G-\#�G�Dj�޵V}L۴���'��}����1�6ѾH���Ov��@K s�3�C�b ������n��p�^�������	5������e��$��󀘙.��� ]�?)��،�E�zd�`����ʭo�Dʠ�rYx�������N�¢|z갖��?�?w�k�>��@�#��ߢ��ʪZ��B���GE*$s>�v���+�$�	Z��t�St��� ��o8��Z�F0L��i�Gz���́ �<�!?]f���	Jx�n�/�r�,�b�aP��pu�1Ak��ݪ.�����70���*dZ��]�[�=Փc�O�B�Ϛ�$t�@�1'�%�9��a޵�`����R.���UO�������!R��;��-!xTڨ��� Ň@דE��������èKuxg�s|ݽ{��Hwrn��*���]�"�J#q�
�z
���ZJ�NM�{�mf~�)�be���z{w!zblvmf�@Yǎα�Oʤ����.�� $�?�A
�zY+��{z�����cO#��wyhb}gN�uֿ�IW���O���Z��X�P���V��s��.}�6�U/�Џx��S�B�q�����ܗa�;:�����E]�ZG�J���e�Y�,��T0�r��i�ro�!I7����^���f��I��ё���ͤ/)6I�|�}k�6Ὑ+�_��N��g���<�����g?)hHD��΍��!���	������'nłj ��]��WW�K�����������l�VE'��Բ�IZ>�,P�O����ڤ+�l�Prf�t
)�$l�;Pf�|�`Z��Qq���~i�g�|4�3$�����Ma"�$j�)Cؒ�>$i�3M��@�`i���Y��(���.e7r��-�8mU��4-$-j���t!�nX}M.�˗����u@�@8o.�g݁xj�o�7���!?��B��t�C�;�&`~�0��K����>���1�#�0^� q���NCb��� �V'o-�Kw%9V�.4D�����_���~� ��k}\6�"RP�4F@���uX}j��R��#h�saf�x�v�셾�OoBܞ���U�B�Ѡl�Y8Q7�Qw�ti���^�'AE���&�l+Re����:��"I|?s[�)��~.2ߍGuȠ����a�r�x:�������6��r���	���z�K�D5�+v���t������G������p�r��b%GF��r���W]hp��X;�XP��	E��f������D����)Q]����.���s˖+@4����Gt'���eRfȐ8[P��z
b���G��/�kb�c��X堥�A�y(4K+H �'ȫ���t�R�Ѳ&�R���y��Q�;�fL[�}�$��#�W	|������Y�%=>f1����N��v�8�J^��Nn)�~�S��s �irX��^_q���|��9� �6�^�aA��rYh�D�s�6�+h�񴶥��w�	������f[?!���{R�4Cw����)�+���U�ra��&6�	[i�6]3���~ d�E��Yױ*�MF�te9�"�o�;����W�e�ݢ�H��K���`u )清r�RG�9I�yt���"	�/i���ڳ�y�5\f<��Z?b��(�SE���
Jɠ%����u����ԝ��Μe��[�X�^�ͦ������0��6�����~�(U�0M!���x(�^�c-x:��(�L�~�5Tv	#�֥s�d g����y�Iqph��tu�������(Qs˔�&o��c��V��/m�l��A��m�rc,��#����Q�ha�3�`Ɵ��(�cX�{�^�9F^}����P���vS��qZ��*�M�����@���ކ��'F��p|h�Z`K�Xn���з��򑲼�i9�C��ڡ'p��d�r��$��I�]�&����.�J=���k>(��s��ᚫ��L}L�~��$>łUŏX&tƙ�� =Ev[p��w��1��(�R�A���+��
Uե%����2��}i�G�X�x8��
�aթW�6��-�g4Q��� B�(CgD�i��'!b&R��a��Y�C$���M�j�=���u�:`<+!5�͸�KI��`L��_��0�d�v�-#��k��u�^�p6�~�I_���gTtQkd��28�FUm_�q*Ю}K�/!�&�ۇI��T�t�O
P��{ެO�|3 �B||�h5u�A#�^7|�@)����Ԣs`m��!kP ���s8������#@<�i���~��2.�I��k��c�ʙ��=P�Iϼ�'v"l�Cj���pt�aD+覨띠l�cΉc^f݊��! r\�D�_�,±�إB�#H��kmsh|��ɭ�d�}�KW�����yR��EU�Pti����t�Y=�'���B-���U��D�z�ga[�Wlv����"'bv�d<�ҵ��rA#av��7yL>���z��^���0!5!�P5�﹛Yr����]��6�)�^�RaV�;���<�>Ú�8E}B�]3�@��C'9"����ߒ�b�JRTK�֕���*B�{SŁ�/B�����~k��>�:��EG�jw��Z�i?'Y���V7	�F1$�)�����C*����9	��o]��8��B9?�����'��e`��z�����!��Ӵ ..F�V�4�1�%9_J8��I{�,��^�ʚGa���l�����(j��a9p��х��Rŉ0�Wr�%���ڨ�ݿ�0���]�N��lO�
��r�ir�+}&����d�f�������⹪퇈��A�GoAH�����\w�����;�kr��}H��EE�r���@;O��Ku��t�t:r�=Rs����m��+�DLثA�U��b⭄�ٰ�����&qe��	��+i���at�#凿�:�q?[T�bo���X`ّ	&����q��,W�A e�~����KS�1lU��=X���g��[�j�7Ps~��)�����'P`�u�l��x�6=(҅�:xMI�'ߋ -�$+��\�b� �BM~x�[��*q&��N�A�R	�H�}ہ���r�)�/ʳl�NG��QR���?��'5~�b�/���dJ4m#��oG* w���˟���^�Tw��iM_�=���Q�_�ﶃ���9��f�jJ
���-�?��
4����=Q�s�)��Q�'���%?�4�h�ȧ@LT�$YՄپ+٦p6*��{6�Ih�]M�m�v� E�O�I�&��*q���+[����Z��~0Ko�w=�kׂ ���5uA�`c�h�4b�ld�0 ����oi�Ί���To���-�j��ZjC �Eˠ�o�@t]���e�/��>��F��+z���<�;��R�o��|�v2=e���J��FAI#�������E,����'8�IC揥�n�ly�E����Ɉ��'{w�3pVe���Ҵ ڝ�ݽ�円&7G:e^�l�vv��}��"Jʑ��D�߻5z6�3g~k֧��!�#���E3_�jUX�I2}���gtG����>A�r>�ǯ����2���vF��MF��*���\�$�ۀN���p�w�ax��Sߢ5=��A��6J�$�[2قq�6��������_�Ϣ�H�!F#�o Q�w�gӢ��s̄!����K�t?�u��_��v�0���hIm�<+p=��`W�Ԑ5��r��[ϯu��Qt��9��N�e�����P H9yI$���@@fu�ᚠS�B��V�ʰ�/��SΉ��s.R�$�H�}X;�nt�vl��&�G$�ں@c3R��J�,� Y�j�x1�J(��1��Nn����*���ny�Ŭ!����|�7<,}g@�:"���H�x���e�}��iH�
8�*�7�䝅�C'b�|���ׁ����� ��򢙾�s��,��-˓�����L�u��P�w��d9���}r��=��^�9k�N?/�mCv�A��>M���^xP���slu���9UR����-k6��83�-`=�˲h��j(�V9�v�:����������]{fӠ�1h�%�$�+���N-y<%$��.L.R��:(�!pZ/Q�Ү�X���>%5���<8�C���9��cqC�����ܬ��Gj�y�w��5Sk1|���O�srB��l�S�9�-V��.�2pp�^f(^no�ʌ��gǔ�{׋�ci|���ԍRh�vi���E���4A؋��W�<��p�JPT�a�)��7���'YIM�C�:�b g�*��泌����* =�奻�"m�B�F#?j�@�f�9���e�5�[r:ؕ�H%k���?�Dz�7"��|�q��t��Sј���J~g�"8�O1>��E�2j��p�v��.��xK�a��(��5�Q�Er�k��(���g�)���]���D���b���q��3@���NJJ�s������4tx:+��ݗ�+PT-Y�	9�*��i*��I��zs�`Ŷ����|�_[s7}\�/�8�'�)��J�FV�qq3�-G�<(�O��\��5t�*V�����7�4y{eo=1$�kz��
<m3`tg��Ag�r���yV�4���������;�TV7pzN~���<�X�i�4�0ҧ��Ll"�z��sϡAz����NOf��!�M��+�f��$��>v�F����*y,��l2��}�{TH���V.��/#ޛ��R��^�1�(�:N�#̔ ��	���'�0�~N�ԶP�'��h�|�_�Y�3�U:`+�t|5��>jXRߓ��=����"s�҆��gq[E�#̘C��������9B�=�) �h�C$�0�Y�.��3E�[�5h'<n3�Imȸ��77��9?O"���O�� �+\�bEv��v�k 0�T��~2 /Ǣ� `�W�9Fn&1�ʆ��wv��~����}���бגE8�/;%�G�w�Rl��<�ʋF�O音��JnQm&�'`��&��Q��D�W���W���Oq�x��H�P��p��*\�Si���"�qW�Q�y��8��nJ�,���;(0�t4�02�Q�j�Rz��~���I�pBǳ٪�T#1=p�b<$K��P�����6�<�v���@v�����Z�S�0��I�`k�+��@4%�a��-AQ�/����l�>5fs���T����o���XB��W�B^�!�% 6���܉F+�_2@̫��ð�+l9�KE�$%XB0�|PH�_����͠ۓ�t������Ä�M���!���K%:�t0bzFຘ[�T[���t$���E��zP�����>��8V2&d�ͣ��c�P(Yi�rP��m*аdت�C���#n5���ǬSo���{�#���z3����^>�$���4�ujؚ�*KCV��^���9�RV�T2
O��k4�U6��㱩o�����!.hS�	�`Zo�3�/f�u���z�g�5�鶣�&M��/��Ub�U5̞��~I^؟�	����d�/�k�9�#qW��TNՖT+�4����h��t%��y��}��t�C��IIӋ/(X�@�6��;,/�1"PI��4���G(:��ͥ�>��Z;ǪX�kla"@���e:�51��'�u��{��V�:GI|��r�}��F��(�@�F����#bMǅ�+�Y��H^����h�{3�TW��s�
v�{]n�ف9�T{#�pډ�C�c.���i�WV[��@v+ҟ������<���G@/���]�e�CS�`1e:��g����}��UOӝ�_'9춿���>.�G�͠*�&n5������<��=J��>4�a������`C�`�e���*kBu+�&a����P;�������eM��c9r���&�w��M��8/M
f�J����H$�/����lж��;L�zP�X�gxEXr�z�NB%r�UX��-Ws	�EgJ^�`c�s���:�ﶢ핻��w�A������JVS��'HÏ1E)������	y�p��~��=P3�i��Keu��i��c��f/�)���8���qd�a�`�����r���fcw�@��XoB�vƱ��Hŉ3��m����@"�E� C�Xd	,�^�Ż��v�zP�$|?��O�&W��@��%lnI�c�����X����T@���js޽��[�{�y-jfʞ���^����CU*lt����R^����51���;i�&8"$��p�aN��8�e4ʦ(	1Ԉ��8�:g`4��x;��n���V@��@5��<��Y�-���
p��m]�/�i��<�,  {2��m��P�7(����.,��M��.)���e�#��*�p��q��*��W>V� ��8��C�/V��{���.��b���<��'�`c%�aT��dS��f��.��*�!:���.��ߊD٪�]� �˓�"�n�N;��|��#ݹ��]�:֬�N�=^����AB��-4Ru��$�����Oީʐ�{k�S�����1t�Qq�;SXB�X�eͅ�B��)��+P�"@�ѵf+g���myj|���`�z�	U��m3\��~e��������`��:�'�܎쬻3e{�-�_;"VJ�t�n�^">>`�~ Ijb�@����q�bY1u��{��U6ýL��ٳSn7�E�^9��i�~U���#�f�"�()�.�v�6�xOx5�='��Bh�p�@�;���Ƹ��VQ�׻��>��nO!u��*X9�I64M�,��)Q���nގ�:�q���+��\�9���L�F�ƍ�����}��9O3G M��/�OFt�i,`�%K�m2��D�/�.b vw��qJ��Xh�fk����l5��}u2S�$af�,�V'�6�&�@,^��Ƣm��Ie#���n�0	�DQ��L�� A�i����H�Kֆ�����:�?�9�2��k.��b4�o9,�6#{C�|�{���gO�0�xA;u�ʻ��zz�d� An��"���q23��F��������n`�w������c�	��d3M�|�j�F.��q�D�[�:G���|��ݴE���	�T���q_;�G��&y�����߻`K�E{��@ ��2�n�4�9�B�,��0T.W�q;�?Y�+aT�-)k�#�[̍���)]+{W����KD!Gt܇�jh��r��C���k��������Nb$��Cf�������cg���L</_n������z�D���*
<�QK?
��������㲍 �<?+�)�ry�,��	H�΄^���=z�ga�ǋ����0N����@~AU���m�����#\���&��Ö�+U�P� ���ccC���~Am���#	=t ��}�	�87����0m'�|�m�����2��A�i1j��߉WU����6g�J�4�<�>��ڍė�I��O��Ma�E�LA���B8�ʲ`PiN�r����y�))�|&����,n<}D���#�	W����H�(zp���=~�xĸ-��Z!xI�5�Y�ώϛ�r�$rI����J_��!�-�f+C�hߙ:j,��5Q��-�b�HDjvG�H�[񐷫��NB6�l��	ʭ ��B��Jw�AYvw���ed�j�ǻ�7~+
Xso�R���������� `*��C�.�`�Trw�=�<�]e���y�hrloOr�e�A~՗��LA�j唡%R�>A���p8�5�n�y-J��}ݘ�\�S!�0�U�����O0s��-KI1E��C�r"DE��6�#�	J�:����0	Uv���ߡYC���:�2%G�9zδ�@��h^<$���^�\Cf%*�*���JQB�ބH����Yzqu��ngx)��"��w���ť��w�]�Y��˔x���t��$'ʊ�x8L�[#��MGl�_7j�U{K�Hòow-0��
~'у��'�>�x�=�A�8s��"��~�6��]��	��O�M2��
6OŃM����/q�瞫[�>Hd��>;����'�ga�h� ���U\��6߸��U_*�V�)@�O���f@0w��}DNΕ�?�l������>�Ǝ��_N1��v�ʈY;ɕM�H2�c�҆;�i#�8��I���k��쪥�������9sJ�$B�5�e�������Ҧ��RE��^�>M�Tn'])���E��̚���[�#���*��h-tfh��,!��m�G,Tջ���x�E��0Vm��T谆
*�{]?�\(�8`X��Y�&��7�}=��H��T�����Ͻ�<�/TP0U\H��1���v�6-1����IB�o�CL�eDl��N�l��/���8�����X��A���'ʡ��W�a	����YN�*¬ߟ.���:��\�v�R�J�&p���$��s�w��fw`(��L�����(;�]�Q�:�? +Џ߄���O�6S�ٗ*w6�����T;Rx�l�tZC��1��A
׿���w�kz�M�psqT1�!��ݿ�+[��AIa�v9Ԙ ��~�4Z��n@R�6;�������mM��Ky9!B	?���{��%|&>ɹ�}�0���6�h3bA"��;�Ɇ���o���㢯M�0G���NuS��Π5���B���q��!#�Zڲ{"2V��x¬H�������$\�E�����p�_u|+�r<|AxT��k�/	7~ٳK��X���p�@�Y���tt?3����a%�Ɣ�fw���`َ:��K����3���'`K4CB�m��d��@#P��\(ѧ�H�Jx?��#��j��9F�t�SȊ�H�� Y��%Z�y��I�C�$�_��=���w����:�PiŠ.�$��A���pNU7�u�'���9Ӱ�K��o����TGbv1�����g�|��\>�i���	��n)T �5/7��g[2�Q�h��|�հ����;�b�Y�G��z� �>�y����Dٙ���ح
��2v,��f%~L��6�E_�#�u��$�d�����Ti%vjҚp&��u���NT��� �En��8j2Øj;�吱�-`!n<�3� �$xT��~��[E�#Ν�A�<��"�%��&8��N	e킭��hV�VP&l:��8����jJ����Une-l�h��_в���4 �A4q�cv"z�� ��2p]d�G>��N/i��2������Ap�I7��(��'e�^������DU��9u���P�HcU��YPT�O�!��M��U"��RE��"��B�D��Z�4y�0F�7\.��h�v%��üt��iƅ~���{�����k��Q��Hw�� 	��������46TY#Y�
؉�%��/�HҠ^s�x��
|��?�1]��֡��C��u����>�F�)K���$V�"b���(��]v;����m�� �b�����%R A%��2�,L�=΀۞+U����å��-��tL���P��	�O��u-?bbĥ���L�ղA����9s[��{H�%�J�l�!X;֯+�6iU���9Bvɨ���mC�lAX�%�l���$b���@e�~o \�F���o����\�2��d�(ҽT�h!��:1��9�4�����0P҇�h@`}I�ǹ	0,y	�(B�F'�=M�1�?@&�s ����������T�{l��I�h;��v� �=���T��5��Rj��`I�b�QAI`�ˑ�VTW~�b�s��l�Ǌ 
��5��>@�������[��G�֮�)��(ٚ�D��m�)�6����o�&���o�����(sW�I�~�,0Xv��+0���=W	������JyO�d�j($�X�(�8��A)U����_l6j=9ԩ}�������T �͈N�bz��� [�"�֎+_�Ť���4�p7�����>W��`�`ܳ�:�K�z�Y�YV�O��^]A/[��k{�[�@h���|�tk�pKMd2�):� <)2<�&�����}\�6����R���{F���bz4��»�?�Lꙶ�&x�����陘B����\ ��S��I��{Ys�k�>�
o��2�3ך�v�k�"��*���L�$�w	8�
����6k�A��K&���P�]� �G��4�'KY���,UE'�+)b�@$Q����u '��wl?�G�B�xˣ��w¿3R�-vC5x�����d#��ķj-��&�
��8�j���d<ϴ�?W�͜�~:��ad�7��|�_��h� Ɠ��Q���v��]	�/3���%�B�{�`�7��]��\\�f�IV����� ���9L�<��ʁ�m$�%S�띏�L�t�� ����f.�E�8���cI5t���O#�n�>�14��I����Ss��_�)w��V6�S�&�*��Wp�S�D5۳{�mF��Iך�;X/��� i�dn�<m�4�@��_-�M�1&Z%���'��0�:߶���=����1�{%ّ��r�C�o�!�&̄�b���T#�&�6��0"�(�b�[���
�A��􋛠�����ڞ��q�%/�-�*��nI{�U��`�Ù=�a���V�>��?lx]��Xѳ�-C�I�7 �����ث����m\2�lw�l0
G4v��b*�/C�����xh��3�'ix��*r�7{��13Rr��9)4 �z�:)����I[����d-����"�矬�}dE(U�qN}���ͧ�W�@e\8���i����ۃ0�$�{��u6�Y��7���ӎ�sjz��RSJ�ъ]Y�b5΃�n�2�UU��g�dL�z�+�/`K����a����(ۮfQq' a����pY%";2WV)G��1�^�{;�nӆW6���"S#o���� �U��(��&��OѲ4�C�,����gԕ0Ͽ+~�V�I�4����C���2�c���raD��"������&���X�E8j�	mʸ��ߨ�Xko����k����㋊n��o7��_}��Y$����1�ژG�s01D�*i����f���@���ܿ�a�:�&j1��T���B�2/�=,�Y81���\�XA3��C<^���/}�G��Y�&�U��7q�>L�q����C%��ޕf��NO����R���+�(�^߾�'��:>�<L�M+'�X���}���K/ �H�2`c��F�QJh]��R�N��␷p�[=u�	mI��Jh��,�B�r����ֶ]&��@�j�#!�rY��L�5k�ƣ�a�cҫ���-�Y�A7��`_۷�{�� ҹ%#�2VL'$�O����7��'ҝn�^r��V�T8l��3��~��0�q|�үh0���%J϶m��� ��UOY�Z�)�i�P"ƩE9�n��7n|dt#�x���c�Y?���E����)gm��+RH�a3��jc@B=F÷x�=h�؆��c��b1��|@���u&(�#�[��IU6[�� ��n�5�am'F}��;�i1�����)�H�ܪ���ܔ'�r��U!�=���+5��q9�Z.9B�G�ԑ�MY�kg�r5z�����W<&?�,�-S�ΐ"x�֍e�]���]B�Ujm��ȣ����W�Z6��r3��~*�t	D'Ǟv/Xfȓ�)��b�h/�����{"�u�æ<*��v������r���g$�i��)�4��cJ�sƜ�Ұ,m��O/���e �
���?U���͂��fh����*��i�����^hĳwz�
[�]�i�zf���*�ڮ[���]+]�x�B|��:/p��qsUE�!d�n�h�)�N�*"]���Za��Bs�����LBR��>y[�v;��R S�KsfQ����^��h�ƛ�)&�{3'_#cƷ�A�ᬃ���[;�ro�"m����]7��k�IO�`a��3�j}�C�i�Ƀ���rL'P����Py�>��]F�BGY�v��5��6Hk��"|L�|­�!v'B��x�߇��T����l�	�R�s>'��֥��ʺ�]�T*��r��_���Q��W<��2�W�n����@��*T�W%� ��X��`�qq~�;�A�0'�/H�F��~��T�'�sIG@w�'������K�AcE�ݴ��k������1wϷ�*\J	:1��I�L,����Q��/_b����a6���IS�2�Q��Z���7w�f��%�M����� �W)J5�p:E� �e'�3s�*i45�X���Gxbz���J��1KcX76�[y� ='�^8o��H%��x8�(j��B@'tfVS`���s��Y�[����=����y2!l�*E���`��&��N�sF~Mh罢�m���7��$D��َ��j6Z8;r�o>ƎY��#�n��Q�E�Ag������+��Ǒ���;��z��������}�9!��qN\����o{L��h?��N�LUm�����ԊF�(V��ӜAVez��K%)�7��LL��p5f|6���~�����Z�`�"U#6t�m+�R�2����O䮚�\F��:go|H�[\�+y�xqgV,CG��N�H2�p�+�2�y	�v�T�� /���>�n#��*��%/{�ђ)q2�/�U�0��ǋ�c!'������@�QT ��w�jjl�L�)�����F���
�����A^
A�:>,BK��i��Xʺg�U����f��1ʀy�0_���
��Dh��E��(#b�&�#��U�!��l��L��,q���W�ܠ�|��ߜ��R�R��4��Wd�aXV{��0�~���N� �G�����`�����lRڀ�Ӌ�sN�;(��l��-�̴��P����z�U�����t��ʺ��֏^�#�S�v���p�I�J���ţJ�ؕ�$���<�qO{���ׂ��dO��ϤƏ��rN=D1e	�����`+�p'תI����K ���܉��(�r����w�o�I���:8� ��_XU�Ǎ��o������j|���`-���d�a,���_�=����U�L� � y��B���3�`�5U��g��)iSR����0Z{ � ��H鐨�ѕ��DC|w��6�y�2�2^@�z���(v��Ɓǔ `�/�+�dQtL�h�tӰ<*�E�9�|j.�[��r�ɑ��B 7_  *Q+���^����;�`�ҵD�1 Kﰀ�t���;����>��M�XFiD,�5yl�Ġ����"������!;���Qr���-�M��._�*|��c΢uV1�$_���W&/7���a���Yڵ�*:>_�-lR��(9�j��(���i$sS>D�;�0�k�\�������$"p����jZ��.	�t��q=P��l�He�3�:�сf�(/{���%N+%"0 6,]�T��k}�[�}L��2mV��ɰhC���JC���$��.~Ҙ�I��'9D,-��>����ؖ�7����]�����=IM�ZZ�w.���Pj��FM����Zc��~xD�B����RD��D���&�Tf��ޔ��(�F��_<h'�! �G���"`44GJ��s����\��+�'�ƨ59$���Y�x�y7N�t��C4k�������>��xca#�:`7n��vV'_ŲF����� I�w�<mu{A�G)��'�}I���y�4�"/+v��#��nk�d�.�(�4���&�Qp3r�@�֊֦9*�5Ye�HJpRKA��*��l�n�}�+��<c���͝*����c�"e��a�}�8�BN�k�l��%��Uk�zI!�g?e��W�s"F���<�r��$�铔��_��	1�)Q�H�.h���G��8���5]�sس*X�V:)�#�'ɣ�$�7E�{'N"�m���JD�E�}���Y��M��1L�?���z[����4S�t;,{Eb�8����,|�&l��G!U �o(E;DZ�Su�x��ٹ��oXn���]����B>XIo��p��V��WY��Ue)D[��
__6k(�3tr��Mp�M����&�t'[���(�`�����j2��_rÎ�g)�nK(�#k�L��_u��#1��0䭽N-���&���%��,�Bv+s�c�-���#���L�"���B8j��HD�=[�G]`O�#�@�ڜ��)���+|�Xw�D-�R���f���ˋ��w�"��U?�
�.�m���tj��v<��P����{�1�JxP�_�� �mx|*�<�����r��p<Ԅ+>��R���JK����o %Ŷ��~��D�5q�!Zd��㈸��=�vo.��3�4��ȳ�R`�4�Y�UU<����Z�ى���پ�J C��L��6������H��Y�Jy��yׇѶ�k�\��[��'�I��T���3�~�t2������j*�"6$=�
��~� ��I�(N���Y�q�:C:�x����CI]��:7������$��%�d�{o*4���<�bMUJ@���>O�m�_�ȍn�c�m�fRu�� }*F��_�W�o��rvי=o�V��@c��������1sc� �2&�8���=����k]�]jz�qUVj���A�iA�_:{U%W*���� ��k�!N���� ���
)����_�EE�㝇��
yW�(ە�)�^#\�{���\�"�.R^X�+� ��ѥP���Ӯ�˔^z�\֝�`����6�])��wK��J��IQ���wݞ�q'նԓ,<��P�%��f�誜�����=I��|CQK4Ÿ�X�ABqܪfR �{&
��n��( ����w;bY�۞���r����������u�/��!�Y��~��[�!�}HԒX���-}�bK�[�����e���c��s�!@u��
2�{-�� ,���F�|{�A��mBd|�+��IR�1���9=4OIx;dUB*�V]:�$� �E�p�T��P����$�4��ɴX"0�9� b"Qw�ժ�+�v�
<���J��J��T�O�s�����V2[Y��e����h�d�=�Hޒ�ݨ@�]��cj5�b�p���*gi"��zUf�B�wL�̿a��kO��}�-�V$��0C��WA7&
�G��c=�W-{�2 "a=���Whv��xy	�j�3��VK4<���	�������"L|����G!� .����?����(��b1�+E��uvks	Y�WwU�v�@*��O�Evr���*��"f��u�=6� �\N���{��NC"9�p��M���f������8�4Zi%�G���Z��v  ����(��qE��+�k��O\�d	V�l��5+��Շe�z�E{���	Jr�P3ܟAڼ�w����"`3��4�� G:������ߥ��kU�L��h�<!��%���u��i�-���Lx{z��Gͼ�N��o�t���j����7��,�!E��Q�G^U�۵��V;��z�Vu��)T��EZ[3�Oy�4w�Xl�\FS q�BW�؝��>�eCA��f�*?I�m:[o/f>^����	�Zg��t�p�&�����
+�yt�o��|���:�������=�#Qc���x��{��˯�0��>�k��Vg^���n���tT�u��4b���^B:�8,6�6u�=6=���_j�Թ�Ϣ���P�����T�� ��iO��ݷ�\9Mg����F�[M�>���M���]�(��<�2�o^S��Qs�N�zK L��pU��f�A����_��3����d �����.@v���`��fT�:�.��0����������o���N� o\Pf[��C����^��T�}�y�лEp�8$�P���W�<��K�8��uo����a+U?yf\�%j�kɨ���8� ��B8��r�ۤ��Y�QX4膀v�pڑ�1PtS^���f�,
WmV�,R�~���#~�v��!���)�����wU�!nLK'dP��h�����3k��U���C�C|���a��o]����Ф��kI�Λt��u���Y����GB�?�w�S~�-�lo�O�����?Ϊ�
�
�mZ�ԗPx!}��4��
dX�=���%o�i���>b1�M��E�.a-���ǣ�Ҡ{�{�����-ӄg�.��{V[U�hL���y_0���n��<��x�J=��e���n�,b�xԭ��S���<�F��D�l�剆�ݢ6xj�w�9�Az���vئ�\�������+��4%�?_ԃ��P�y@��^�q&���&�L���9(q?:�,���
b;�~�T�]�X�Bp#��~� �Ar�n!�a���$�j��!�?�$9���3l�0��0��ŉL��(7����,�]��+�^1�5�k��L>�{]�5�+��r?6i�u�xR�����&)����h���������@Dn.�Q�bWʽ����v*S��	j���\��aQ��	���\���2��
w ��QF�Ύ�;���n��|���'l��N�K�������{�Ȭ:$  (]�;?;�-�A����b�V������Wt��G�4������V�oe�1Un��)�nH����Q��M-�뢦�����/�Y^:*6`��F:p��\����w��}��"gjsNi++�:�ܧ���;�=��3�ߣ�dU$;��S�u��M�pt�"�D�4
f��.:/16��������f�@һ2����� �i�`
���7�Y�d3��Z+���@/z���dѾq]u{��$��|��!Y�2�KPok�Fc���`����]I����N:F�-�T�vs�`���S�y����k�k^z���^�e���z����V>M%s
��=i��-c4�T1͏�	C�%{_ʶ�L]�SF��0�3��u�,�����}�~��k9�����5���t��[fڻмܹ�6�������e�j�|��F�h�����
y;t����FV<�)=pe�e�w%�(���?x. /5-�k���.����Ȫ��UM�y���}�N{yS�Ɇ"u�v��;^j��\�̎B�M�����;k�6� �?��f��7��a{V���.��Lk=�&���F���!u�z�nv֫^��8vM�F�坉�t�G���r�V��=��uo߫�bÍ<�8;��|i��pǲ}z{ �簅L���x���FK�R���k�]���y=�+�55Aꛤw��x�W��d���=<��!KN�|��G��9�$��h�P��5P�swQ�T���o��З��7X�i��/��s��� _P��5F�SL���2k1�����q�S|��x	�N������zo1	��m-�w[�ߖp���w�2[?剿��$7����f<	��!�/��;��AQ�L�K���oe�|!�YH�w(�D��^�`�U����Ǌ��D��J-
�3���B�6jM�Ս�������p:�N�R�w@����5��Y\�^�,h-�x����\d[P����1�y�N0C@>�=C�:����H4�uT���<��O#����RE�$/~��pTN�l����_�	2�r,īP�χ0�D��˛�*8yv����,�Ï��"H}�moUO�֔�ɌC��)�U���v�%�0��i�U#pZU��x� �G�n�<�"J�>+� ���@
����A��2�B?uHB9 �c�li`��j�Bc�&�4�#�&������(�Q�����Ql�Xr��t��i�( R��@�Q�ǖ�F����kO�j��c"�٧Zk[���ߏ�Ž��Ԥǚ݁)�(w+ ���^������D[�������:��Vvm���;�/AJ_C&��V�%�r���
�l|���I��[B��g���&��X<i�y`<%sj��:q'x�����ۇ{��`���d%|H��Y�5�P_u�؋�`��U�*6��c��@�vY��J)�, �7o�������<�$�������k>���_����?%�%d����&��;���I��jN0��R�r8e��ޓq��xuX�<����Ʊ@|�اD"�/::	nD%��@,�|
]|!sl 7nr֦�<@��&ëdZ��tx�~f�����Y Ph&lO6ۚ��J6IA���ԆD������+�����n��\�ƃzƩ+��wQ�M��ȲC��h�ُ#X�S��iXw�ẇ�����c[1�Ȋ�^T�س_����������Cq3eȒ/�����F��� ]Bi�|�.�@���@�D�-|�ޱ��3�ѰF9�� :�U�B(=n�vp�n���틪o����pj��*���]��B��
�k��{�8 ���M�z	P���ۛog4��aoڟN��[��q�z���VVDeP�&�Qc�n�.���~Q���K��F��Z%7(��m+�ߪ�,>��c��o�7�tV���lS!��d̼6�������t��y�h����@�w����3VPҼ$N���i,�2��4��1�"pߒ�8���	�4����H��˄5K�w�[Y��kW|��
��Q�F�,!�eŕ{s N��cE��-��ّ��0>���~bC誰}/��T����EM,�Y}���1�êҊ��[(.B`ڜ�Y�����A�Ch�s�0�!7��ƨFt�B�(%#t�q��@�V�S�B��#Y]+��ǻ%L(:��@e��@�BD��x��/�K��^Y�^Ě��pt)Ē�ر�s���4���<���&�ð��W�McZ�&;�����ց }x�n[�g���G� �5�B���q
�� ��jAy&������%��fH�.�8���N#l�+�hw�5���9�_6�M��]��;��>�-��Q��Y�^�V����O��aO�jd.�$8��t���1䫌���\7V**�!�D.�4�9x
�gr���� ���,�e��ܩ]�}�Q��Wבd�#��?�h�� ����:�S�}�S6��t3�B�[vHjfmب�tnutj�J��1�si4�@U�S�mv�Ґ��k`s{���E�&�rB<�cfv'S����Yo�3�8�w�ڸ���Dx߱�!�Y�jӷ�u��csI�Y�v���Fz)���*)��\�NjC �������d�"v��9!v�h��y&����ޢ�.SW�н{�9��^���hU�:2ג'�1����2i�_Q��E��EeV�{<�Zbů�#��NEZF�ֿ+ݥ��}<\%c���%dDݱ�J��<������34L䷍?�7��_�i=�J���c&���^(<�[FG=�n@c
q�o�:��i��ǂ��F�<I���y�iM �Y���Gΰ���㿏a�L���T�0��侎�I^9`��$a�KDyA�X�o
o���e�g��! 9��������mD�]J�]���!�/�G�� �K����yIp�~���]�H8�P���=�z,`,x���m���:��PR�<��}��I���WJ��V�7^�_q#�K�L�q����=���S�-i�W����%{�Ӓ�������%�#^\��h��?���@���;�د�ڌ��:��#Ev���W\��wZ?4��]�{ ժ]lHB��dTο��,#oS��q��5� ���e��au]=�Ն��3�E
�+�}�E��3J����fkc;P.L�V��ze��s���;�fUҌ%���0G��B��}I*r���,Fm|~��� ��#�L6wL���-��9Rri�-C�aU�b��,7Pʪ0�H$�=��D�>-b��!��s���7$׮�P�+���a�iz�
S����d����w��K���L_���K�;u)bE�{ϋ�x��R��r`a�T��/��W��y�g�J��������|��1��{/`��w=����M��.u�1���|���x��j�֘�9שMM�b�L
ǜԙ�ȈɄ���{w�c�AǗ�a�Dj�+*������罗�>>���۫�>|� N*H�1�)�ba������rc�1ixT���*�bOV�=G����q=��iL�I)N�OI3�l�ɛ��v�a-qC/K��%��W�B�Λ3��rų��l24}3%��JB�\�޳
����X�>qD~4�r��^DT�XNę���	C���B����'�&Q�tsI��ړ��V�8�O��A�9����b&Щ���y�꺍��9z��^������'@�cZː���tB>r\EWa���K����Ƣ>*/fhݳ�^^+��D!֯�0�g�޻�xǟ༄O>C�$gc%��&�{��ە�0�0�_��9o� ��R�-��W�a_�K�n��s�E�;K���=�4,A����]�8��-%������qzq�sB��J�pW�K,�=Q"z�����٥�TϘ�b)U6�1K�Xĕ{�8O�>'Dt~��|�ʰ�$@٘m�Q�����*u[a@�d�7��E��02���C�.��q�x;���do�.E�G+�u?�2׉)$�7�al�:�,��3�b}k؂e��b���J�&�X��_��EL
ׅ��
�6�+�O"�T7z�X��P#�S9�n'�]u��Fo��PV��y��b邴�Wܕq)m��?{4>��E��;(��vKn�E��VzІa�@1��³�����������byOx���a�3eG]#�&�m�;��\��Xn�L�T���tD_Ң�JSk�|$���{�{L���a�r���Y����dȝ\y���G"���H�r�]�1�ą���b��K��-?:����0�xlI��|>,��-�B�(��M����Α�^�<�Snي#'~� #Ҟ���O�$�dD�,`�'�7%����V�BAy!��?��O��2�º"I��a�;Q�C�rX>�f�I�mst"�����  �Ji�E��,٨���k�-�a���\��)�
��8��}�प�_�p�C_Z~?���K�v�+@�<�z*����P���wA��#Uy�Xj�&��=�q��a���Ol�ʿҿ�_)\,��Nc(O�������X��\&����i�� ��خݠ�ui�KXn���Wq�Șv9���1�c�
�;���B��=�βːo��6�͊u�2��{*ܚ���&�a�^dG�ŽM��n�d!�$�W��z1��B��̽�ϼ�# |q��z~o��RPm�pH|��=�����,�g�G�n�Ϸ���G�W��������
Ұ΄��^r�#+��uõ+������h�S}q�(�KEc��ᣭ�ŧ_'DYH�]_�Y��/�mf�{v<L��s��E�)�U�FJ����}��w�F"�	9�c�N^B�y��:�?�I���(�|�XŇ�uK��4b�~���t0��F<#3�'6
�;�� ���S���j�K��5Y�"[��`�=�HD����a=��������`�T���{�Ö,�*�/��Wz۝���c�=�QA���J�����\��*0��$�P?�x��u�`(�������6Ux9FNu��o��Yx ����������e)P��\�pk�^��F��4�K�4f�{.i����ց�9��pI6k�l��詾߃Ώ�ۺ�('��i�z���5�;Ԗ%�
�^�_��R1��{�䈡J����-��I4���"�צ���Ė�oH̘�̸�2��坦D㌓�ry�P�'�H �������Oo�:��w�6Ͳ�NId8������.�s��X�z�J��ןӡ��U	�[T=���$��dKu����Ai%�I�A�Sn�j���@����z�"Y%Át�|�ުPz�5\��i�^��)�F1���Ѭ��v�É���Ce�t���怨�K
���#��-ގ�,��嗰��a�{���ڭ.u�B���ҍ9T3F���D��L݃)��Z���7�<�`'����66[X�׋���N�#K[�h�,d��4I3�S �*���f���O��j��ҰSj��H����"����s 
bH9���.v�x��ME�f��νm�z:���;XH\l&��r�Nnף6��[�,��J0��&�S�,T�I����j����+GaM����sd�H�Y������e������M��E��XO�c�AR���|b�O��Tv��5�]����K)*C~/>�O��Q�ԑ�E��

�
P�O�G����+���|5����������ޙ�;eU �`BVӹP`���J�0�p�����؝��'w��a))c�w�/�c	[�������S�T��I���E�kn(���J�S�飥46W{^,�T,�x6�/϶_���;7�۸C5G�Z݂�zi�]��|�f�r���O��9gɽFŁ��Ym3[D����q�Ե�s�E�eYHNv����ot�_�H���f���c/�O�_�����oA沸∝��K�r�YueO�Y���B��yј>�[��e�t����B��B��Q��T-WC��H�vn�R��ttz���+���@�/��ȍES�����5��Z�ir�|fe@"����ູR+����\MQ�{9�R[��hz�z�76=Fҋ՘G!�lOD_�&R��]�^'&���$:�4�z��߀4�J�jĳĦ�-�ri�v��%Z�X���j���S�/�G�x΃���%a/Ɔ��K7Dʥ��2P<��
�c��Q��٦�\(�d�P�?�����8T�B6�|�ȑ�8"|��o����p����W��o`�@Eϋ�7��F[2�:�?��W�$2�P�y��5c��}B��GL$�ں.+�
���7ip��k��a�r� �vd[7����m�ġ|sq�	I�15������G��u��;���Ā���C�����	�W8��yЗ�Vn밊|��fCq!�� �;h�^h���6s�xQyb�4ZZr��<�PZ�d��u���2j#��6�΄ �d�����_}頗���mϋ
3�ʔ��S�Vn��0�)I�n��>�e�$�,��Q���B�߳v��!�A�� �B��JWX0�FJۄ�bs�g����
� �����΁!KG�0�GA�Η�B��w]#��{ӱA�
�{C�Ƥ���)�v`��fo���l-�ґ�G�l��.�3*ǻ\�1l�)l�sL"��ȤvB�W��,�$�	��Lc�8�$o���,RC�T/� �{J�}���gz>�l��4�G�/��6l�*1�NDVI~ t��Z���$�(����o�H����{⛒�t�}�p�:c� ��y7��92�CR��N3�(����OJ1������`�v� �6KVJ������]�	��jE���,��8Ȼ~O\�w�7̇�Z�����ȶ�T��*[��LՔʃ:��f��x�����#������G������q���dR�P��=Wn�~ar�C`�}O'�����{Ί�@����/Ə�&~���qn��V�#RUw�(k2��q/�đ;���2ӝ����B�����`�����=L�2�C�<�-Z��-8�c�������rߦ
\��`�좐���2y㚠�b*`��y.�Bm�~�?Jų#����Y�~P��]�j�>c��.iX��ڔ��'�'O�]w=
��t�j�a�������5�VU��G�1�<�m�4A��7�/~W�ˋ��NhN`���ϛ�J�]�2�.@��ʟ�=��Y?������ZR�ǭQ-$�l�2c�Ff*�q8���{�l�fWB�B���N���_<�)���m�s�t�k���F>v�=��T�0�e`,�y����ՙ~�VX0�m����>�O�dA���h����bd1�x59��
|&�z��X�ِ���ȆY����\!�J�w:����$!xQw�G�3iP���/�F�ٳ�5���\��C`�| rַ�������-���S$7���?]ksP��� ^7�z?��q�z`���Ec��Y{.sN�K<P���i���{F�C��Z�\|�!�*�!���$$d��I%�f g30�?�dA��ب�v
6��� ��g�O�6��i8Rn��a�bZ��7��8,��h4>o`���Ȇ�?L��&S�]��eg�i�T�VcM҇A�HՒ � p!�u{��2��p�ݚ�����ɸ���Ѭ�0��2���L�$ǻ���*�/��e�Q���<}7�$}�D�<�'�X\�& ~/a�ұ��P�T�xn9����u��?߅� ��2$���<N�K������p��u��|/�����LR�yŢo"�S��{�HS�w�?���p�?�3w9a�M�4�G���=��.�.�~&�F�&�ْ$�p�[��T�O�6�B���W���Y���K۹�)���:v8	8�{mS�Z�F�N,�Єئ�V���C���#Z��|�~�>{�<�<�X�E���潴R2fI5_��������U�+��~�]�^)$u����U�6���B��1$xB|4K8�sn+���A�ud*����w�W:�קr\�x�o�a�xڕg(���2����q��]ʩ�(�p� ��9��^,�����(A�:���}��� �(�N�S8����bN��^���W��iO'���ñ��'�Wq�i#OnZg�9?7b�
 6�)o�p)�+w�R�C�C�p-��hiH0���h���!y �E"�]�'h�c���əvm�o����@'s��H}�4�Rů��w�3��&PC��d��)�*j�cl9�lM�<�7�@�y����Mw/�<�{�@������S����P��4������Q8[ՆK��&	�b�����/��4z s�_~G~(��70�oV��"��N���R�%��8x��������4�B����!����JozqY���ʴ�/7#�n�F���B���zN_����\l��Iejb�ta*�K��
ը�)US-T��C�U=��,
c�Te�7/a"{�)��k8��e�lQܴ]3ewu�V��زX����v����l�i,�P��Jrx�
�V(�j�n������c�8�L��f1�T4��m����R��)p�5M���^\�f��;�0�ܮXv�m���@�f"	K%�L���SDk��_[�\��XK5(�e����u^��:1����¤���iU]Q��O˵����,,�1$����2�N�Yû�2s��T�i�w�1�:	s}�s4V$�r�g5�Un��T�*8�}���Ir��[�2"���]j���T��z/&B�˼=���x�A�X��|
qL����k#���5�s������-ļ@l7��By�D3��G'e����/�a�R1�!WbaŴ%�L�ZMa�L��َ]��d��%��!�����o�;'�kM��3$ ����pD����  �Ս9�b���:�?a�k��.:@KP�����q[�A��w��tu�Z(�(<+ &{[&�'���U��/ڳ\7\AO��B��Ճ$��9=���Z���d��L���WtEA�,���2�ۑR*r�?f�
��\T��o��}=�d
I��H�meޖ4y� ����^�M_�XuGmP��:��,����* z�|oRkN5�����_`X&�}�BX�,%�����Q�R�<��(</�[���֖ٓ�����������m�HI��Ej�s�E�ir�)�'>���:qL�P��7�	�M���k��N���[�;�k��B!ӯ���t"ӡ��iZ�&Ὀ�b!�W/{�.	~���_|���pm,2����x�fr�Q���%e��9����Ӹ��_iIڮ|��{�X$G;�~?�m��a�Zf�sQ,��ԇ��M�%�b��d4r��)�Dl��a��Bl��M�@�&�f=L��a'Y[Icb2�T�*;j��䛱�y�|��4`J/�)Td'������W����)IT���3^l����{���]�l�rG��;�<썰������<o�FAL{��#�t	�bp r$[ = ��ʩF�5Dp�QJ��q�᧛W��p�@�dqh�}���BN{���s�C�� 溾r�5I��̸E�O�\�r^�,^��c����9�e8=����9� *��;�[adp��>��\N�>~�Г9�,ře=4[��Z����5T�pi v��8?�;��JH]��h�삔$.����t�g%�}�u�\ɶ�����,`�U��$K�?.�X��<��EVO�d
�|�f�e�H�4�k���s{�_Ѿ�
:@�tY�x�`t䟢,�b�A$�\撍���k����CE�*��-�!���s,+�*��b�v�PfҨ�ƅWV��q�r�uMfHE箺�uo�U�t��0���ӎ�A=��Ww�K��F�@�0�]6�*J�1�w��pY���U�aR͸ѝȔC�,-���]��~Wգ�y�S5m�e덦eU��[�e�9˒E�Mg|]1�f�ȅ��Ihҹ��U!1���}�pAj�]@�,� �UŒA�������Y��j�!hq,b��:!/Ы͙Lu��;�<`x��;�V�b��\
0����W�Jn{�J)�W���+V��l�����9�/rJ�����%5�Ќ���6�%�
�RP�h�ʭ�g��O����fny�8��}!�� ��8��B9��
L��[�TÔcU��rzDf �邻 �9��S��U2(鍁��.s��֖�2d�d]���Y[��f4�0N�xߠ�K\6�j��EZ.J-=��5V�r�ܵB��a��'ݥǿ�	�K�]����@�X�*�#��W�}��n�ݗ2[=Ԡ�z�m���<���D��ù��Hy*j!���Mh�|�v-���ہ�o���)��I�|� �Ť���77���E?��<퀋����iB�d����%M��)1*#��$�7Æ�Yk�;ųyf@�
w3j�}�,y��Zc<���O�Cr�Y��&d���q���0
�h@z[��6�b��1��r3fO#&W�	��K	wU�ث�LE�EY���.>���!�(Thy����.�3O ic�+�yƃk��2>B�t�Ȁu�r���o��S--�T�~_�,���5"�͔)��6���м�D�kթ��]�s.a��ϧ���ψ�A5��B�����܆���|����ft����d��^�2�|�e&h��Ҹ���A!b�FsLZ`�b%��ۢ��բOE����w� ����~�?c�H:�N�J�ot.�yD�"�u�'������sʊ��ne��FXM�jh$ks���4����?�8r�۴�Yr�a�0ȶ�F���M��q�=�
�k6g�A��f�3�%�圐����1w6c��z�;H�]0���āOwk�m&�󪭼_+m
����gJ�sb����!����g���9r�Ws,�%�Z��7�#�*����������*ƌ���Bhq�&'��\;��в��c#?=�hjj��:e/�fqG���x�6z�-����m ;V���"���V����S碗��vg_��@XdլP��w�HsލR�r>�0�YN�"��N�;9�������'�c�YC#�!�G��Ԓ�\*J���k��^���9���)�<��N�m�j�@_o0�P6s��۵>p�m�x��#��8�^�-|l�&�8���i,ٌ�ÿ?4�C���H��\9 �d����P�x\~_����Ʃjg�����\�`!�d��!�XP���8~�]Ŕf�~R~)zg+m����uN��R{'��ᴩt�,Qw����4N�ȡ	Ʒ���c�Y'p��2n�6c!5��d����-�A-�B����V��P�n+�Խn�z���g�e���I������3�;�U�N����&奺�_��R��<V���p�<h3P�@8Ƃ����\�|���{���6	X���w��2WQ��l��(�ǖ���t⼉Z��Z��4�H��'����r0���� ����<�+U!���~�������k�ÿ�3,��/j)��a��Hvh���z`[�����5��������t��C��K=����������g�&���1���k�i���i�8���s�ǉ($��I1�Uz���CI�J���vV��$N�l4C9����|�����4�z2/ ��\ ��s�Wx�������A�j7�y���ɦ�"�9h�  �w�n�z�$��X �D�>pz����+��o�D��y+|\�n�H1? ���S���}�\ɹ����P�Α�/�� �mXGvr�}�'���q���K���
�a�YK�B=q�QNrt���g�xYяN<�k[���G.�p���b\P�{u�9gmن_�}r}L�ޑ��<6E-t������3����ѳ�+e���ø=ݘc73"�Ub����?	&��8A��r����F�ZW����H��{�\S�s8�	���o���+�2�\�L�D|�h K
�ɶ�r%��Q������IX���*�,��X~4g�uC
��b�=۠�6۬Hs�_�R�_g+��Y�q�+��,6n?�7ji٫:�,t$f��l���kH���H�� 2Vs�K�y��!K*�.�-$���f�O��͗)�tёʉ%Y��gT�l(�7ڊ���Q-<����'ۂjs�f���d��c,��C�b�H��T,��"=WRE����/C�Pղ�r�*=\�MBq��n��n��r�*8�.co�p���P3����w�h^�F�v�"z��vh��}��3��ӐV*c*w���k��"�?xY3�;��Ѓ�'�U���JN&���*���U[iWF�fǴ �v�O_"��}ڳ���C$�ۏ�\&7Ȉ���7y)�z��8�Ʈ�o���'�r7�2q����<��^7lwh���o1YJck<Z��3"�
��C�|%~4)~{ Jci:��*f=ϡ��������
f�B�fw�_��AIһͥ\���a�m�Ϯ����%:Y����O��uU�� �y~e��a�o�i��8�NeN�,�G�G�|'�9[�:�o��r!��j{�`
Tz`���)�xcG��tc��OC�ǳ4;�2E\F�<��`��A��״#�?&�jW�.UTao8��`�6��q�uka���KN �M��:խC�狼ۥ��b2 nt�ωD-��磃��[:c��>���Y��xi�]�/�y�g�2�d[ ���]�,9'T�+��E˸$F��#����>9�ʾ�&�m��Ps�`��Ɣ�%e�I:�-U~��/�
]vK�mʗ��:��|��>�֐TR�Z+� �rɭ3�|ӄ������YG�|��7�~j�@"
O��D�M���|j"��K�g�4@-�����r*���ﺃ�_� a2�E��E
/Fp��S�|���?٪j,�ZPt��v�,X�G�LPQ@������+fFc˸����n�{@�Lڽۈ�C���Jn{��g��~i�<�F�,�|���4�|�L�t�GP
k,������E�^>���z��U,J�(���J��J� ��#%-�Q��V�FU��QL���~8�Ot���b�a����/����^@�ư¯G����i��ҕ�ԟ���2�o�U�!�y���
�e�`Y暪 ��
ޓ�$~ L,6�nSV5��ǻ�aE�d7_���?�:R�ká�~�}6.���'F<dQ,�D.�BB�6k|}�se0˃yu2e>�\�5Ky�1��O(��[r��K�&3�W\���)��dx�r�h�BH�t:A�����@ ��z{&�����3�x`�j'+�Ȑ}/�6ȭ�|:�;Z7V�4Sg_����𪱸����$)���/Ŵ`�%R�Je�Vs��-]��z����P]��ߩ���b*����
ѻ��t=�-]�:�X�b�����p}W'�A��[�x�L�����c��}W=!+��͒�	s56�O|5ײԬdE�F�{���b�3́�P��q	[�$#����L-�iV< �߃�3i�IUp���Z��e�6
��+��&�'�&�J}���|ֳX��@���B�u��%�1hF;���o��1���NW�+)M��b/uaV��ŕ����������z�D�&���wj3��Q��N�M��Z��P�^t ����PR�j�F�_gz�x�� /"v�+rrZt���S�p0_��/�����*HQ�+s~���b�m^����˕v�;~G
�W����dToC5 �lo�L�۸�~��P������iT�v{����Oպ�S�5�<��{��C�U�sVG�'�����7�d7{�1ìb ����?�^CG��]��c7�G(6;m(-�j�\C�z�ݿs+���ԙ|r1V5ȉBy�'{�ф�R`�7��ZV��(�O�"DBɩ sy;D������~\\)W��2��K
pYj��)=4�خQ���|��4w��*��`;�/mT�K�c��\�h��tJ�^uE�?��Z��2���X�p󲄘�|̋���wGy�Y^:`J�$��~�$KUL�AX���1�YaА�vA��B!ێ�q���n�(
L�!�%�|��ÖW�׫����F��t&(j@V��0!%b���CE�9��w�zs����_�ViFP���M�>�;x��'`4`��Ғ��%Ĝf�)��� ���q�{�Bv!���� g_ȴ��G�M<c��u���i�/�]^_T�si_2�8�c_c{b��r1 �'��&���Pki��T4�Z9�|��i��C�<�j�L19��v��yXYAԠ�%C�Y v:�X\k���E��{6��I���I�=����N��Xr��d�}n���AONY_��N�*Ca�W�g�~���� e߲K)U��Ƭq�ep֌�<-�L��gO{-��\g����V7�	w�-��MK�ƃwb���x죛�}��y�`4�d>������z);/�B��,�_}����%�C����M^cj(���g%X/SK?8�7�_�6��.b��\��)�v���4�+?��2���$�쥉��l�&��!/>�?J�x�U�Th$iñ^ԗs���3���[,� ���g'�@�����ÎN��MY��3�T��韖<�c1P��.�y��HΙ�;=������6)�	9�@��7*/yI�Z�h+*�w�hف2���P�x4��ErX>��D����i"��,��%1�|Nc��c�����B���2̪s���֭$�oe_�Ջ�}����/��Bh�?^�W6�u8�b�3�:�S��]�k�$E�)15����P���RX<\����(!o�\/"0�G�M�������H�t��pG/��� �b�ڴ �������HV_��&¨��+�IʴY�>98�1�67/"W�A�b$�v飔��l[��ˡv)�X�����J��!��������h��٤B�t�s63��T��!W�J�[��n/�g^Vh�f����c�#�l=؉������K�	VzB=�qJ�	oRt�Ͻe2>(LXڭ]k�+�ҫ�ލ�v>'��◝���a�|z�ĭ��BV� �,�wU� 2¯a��3���\T"c,ct1 � �)��z��Bү�l��%wǋ�r{�ۡx?	���6���$cĹ<B��R�
�;zU�$���B�5���Dɢt�`0sl-I܄�ȭ��B ����B��SQ<�n����l@#��5_߮��ʧ�_,1�{���=H�F����3"n@�ct��`/G���_���څ�'��b1B$�u��Wz��q���q6)y���������=�O|��g"��d��h&�|x��}ڠ]E����P����ó<��N���> �d<S�W�c|=�'��g�����M��3c%���ٰ���2�U�9b��tŽt�兎���|P[��Dk:�E=��I���!��:��h��ɶh����r��tC��i]�6��-ErI԰O/Uo�����+/L�C��>�f����n�l��VS)(B#���/S��\��އ��{e1���h�3/�;�0�4**Zg�f��.*`C�fh �϶<��@���pؤ�ԛ��d����+�+G�/6���I	�*�?���c��LM5�����w�� �bl �EL$��O��&�s��j��6ÄU�?�u���h�%����qm(��2�-��Ԛ�v+ir29�])�y��4n�G}��l�3����/�a�hgV��˩�䋖�y���*뻴h��De�E.�t��5_�������7@��>y��qAʡZ!��ZXO�x\ϲ�W����qo\�r�Գ���奘:GW���ۗB��Ʉ����<�u���r����_�Q�}ˆ��I{/-G�ʕ\Ö��s�c}�[���bmj���+b�����o��Xi	����/����+U	��tMD��A��F��f�c"�~�g�|��h�<�����PqR�L�rg��PF`h��J���a$։�:N���@-�RG<��)|�T�N?��l��w a�3~�M'��A�B|гX��@js-���s�S�
�gVi�=P7����?���j�,`��9�]\m1n�	�̤�'|�dϙ]����{�^zc�6�ø^�\ƍŹ�M����mg}�?G���7(�š"�R�YIz�t�O�z�35)8�;�s>�dw9������\O57x.Q���X�����jÀ+�d�C��6��+FpM&R���X�Dc� ��4�o�#�f �x�����"�/��*,�am�j(����tHf��俊
����d��r���!K��A\b�����()@��f�u'Ȕ�_�b&t�(���Q�mʥ��������^��\���`������<ƕ%!�����۔ hΰ��R9�²8싔 (�1n��}S���x�����s@Y>fD�H�=RY�)���B�����\C?�}2yج��J�;� ����e�s=}cX�4���a!pK�x97D6a&̮Ez&2����8����]�(j�q��HL,)���x!�]?�����7�����N��_�9��~|F��D ����*���<pb�&�$vbv�=�jI���i���Rj4F�	O�C�>�[Ă�J�!�=4��S�,'���������ڎ�n[Eu��	�-�֩�����<#h�ZP����!r�D$�$;x��5O��T%�÷�ӊ�!f�*��_^��?���vW/�?�_P��뾵�\�ApZ��֌'*�뫥INX�96ٝ�d���(N,����}���.�*x̻mB�hw�ثk@`w�d�n�����z���=OjM!�<Ԣ�H<�����D�˶j~X�����;6���� G+?��BQ*p~����m�ck9E�n�}N[���@�Y��+�-���7�-n���-�Dn�ц�0�+��n1NW[	����%w��?n�i��/��*4��(2����+'�����͆"���_����V��C1�,a�0£>�BbT���Z@�2b<�l�5����)��~�Xҏn(�Ͳ��h+1qmT={HlxVO�ivwj������F�99�f�B}�/j�� C�&��O��óp׽"�R|��t������Nv���v���o�*k჈�v!�s�@�	���Ϟ����%j�zb�bĸ�%.������r���y��w���y�%@�t2�B!*�5�|eh�e4|�:���	�bq�`�n s>�&��B���a�f���u���$i�b��G�8d�F+�2��wi;�G��^�t��zT��h�%�h�HG����U:�B�M�Ά���S���HZT���נc��DGU("A�)�C��+qx�tW�Uq���SQ'�=2{=&s먯tʊ��[8�X����V�_�~���s �i��$�m*�����/6=e֒�������H�
�yC���J�}M�Z/V}��޵ڃ+��A����+���P��i���X:`H̿9��_,H�1���q���TF#DN�b���f��lH�K7W:e�M-���>���I���ڃ�rP�0n��}�0.2�C�ꝛ5�mA�3\�n��X���*|�$:��*�p��4ݽ�t��;l���&9z�G`�$����e}H)�E���
֙lhj^i^��#�Z �11iƋ�kp����������>���P�r�t-O��G�s��`J�-�k���Y���]b�`�s' Y���+һ;v8l�K]�XE�bܥ讬~����{O��빧B���,�x�v¸ZZ[�M{}{����Dߒ�&-�aZ���_�\8��n�{��Ls���H�"��훇��wOV�9�a̧b��@��#�Wb�Yh%y�<zO��ׂb
)�u��5��*;Yĳ�����n��!�>���il�O�b.24R�Q��1в��e=��h3X�X��:P��@�5��I�6�T�;آ���Ҁ�q Ɠ�5�RVe�"�7���q�.��'����.[�(�u�Ƶ3L���A��44ڻkzfg>J5��MV0<.���O�wh�JA�wWH#��Cɚ�^�=܍#���/��1o�o<}=��i���_<ܥ�\OP-�s�z2C�rZ����l����.')��,��g��+<}�ڴ��-��	&�z�="�|�=8��o���`㭒m{F���̟<��tu7�h����F(A���)�U�i��2��W`WXѲ<�!W���2fPy�Lm6�S��������)]�eR/߬�M�j����j�Cɛ��(��&Ͻ'j�skYkL�]��4HY��_��"U7+[~b����ze����>�S��]:,ͽ��R��$��v�1�$�s��1c�E�W�+����[~���A�Z���b���c�K�Q���Ia]X@�L�s;�MK=�v�@7L��܇�O��m�O���gـq�8�|���*k^�����K�[��ʴqC�������h_"��I_59=�%m�� )��r�OJl���A=`A#Mvޕx�A��q� 9�W�p���"f�bOmb���>�kk���τZ��bd���S^<��&������p���V�p?��y�Y�� {��QA+�aR�د�-�<�A^@�l@ �r�))2<E�J��������˯�1�����=�]�sa�Tp�˿�j�PR}v{c̖l@�p���F�9(�Ù�
3����"B�J9�`eW��Ю*0V�h�R���X��L����XH���| �m��\�_#�q�ZC�I�w;C���>����� �M����V+�_l0TǽA��<3���v��A����/��akNX�j�4j�	X:���<j��R���>[�
o�ښ�B��@G-�b8�Mm&c�YJ�FYGW'���ZE����>����s�:��5'��Ne�B&j��P���vc)�-~4�oO�w�6�B�"?�^sG`c�p�˷W׌��!��:���U��%à��K�}�Z%7�+�}�R�V"���-Mf�nD&iܢDk��( ���Ͱ`AG��8�����O������D�#����*�k�:���g�=�"����c�:��a�es�ӎ�2���b��������v�]��w=#�ކ�:���fȦy�u�Mi:�.Y?b��{�8��l���b�N�-��n�R��H2�0���w�����+l+�,�4E����>�����v�������
�=��h$� @��������,�Q{��y+k¸{��6�W�o���E�6�ˉ�yBK3`ݼ��6!J�v�.�uZ�n��`j˩Σ�+�N�ٌ�H+�X�`�׽�#�7g d�j�q�LpӢ3�$w=&`=�% �fK���D��
p&3�7�k�a����l�W��e���f��]�2�M鿆�O7�&�WdC�A��[�^c+�q�#g��9�6tZt!<�(�A.�����P��4j�љ�b�_�������:�\�?� ;0�쉸���C��3sM���Nׂ҃���L�*�!�V����DMZ��rZp�\&Y�ߢC!���Wb8i�� 8�h��:ѿ<Mr��k2k�x#�����s�c|���iF�a_��/#"}�Ҵ���M��9~
��:j�\[��Rwݹ��Ɯ"��u�ƄE�l>l�l�v��u����ʍ$33��M�`�w�^_���u쿰mN��8�BF�M"��A��Dֵᷯ�p�eh7I�#���v1�R�>�o2��Ԯ%)��m+c��C�	��E�9�����s��(���'J<��pឨWo,]�O.�h��לk�����ݯ,����$���t:����P��tN�!=O ����|�e�^i��r�I�*�Kd�v�W�Т��ڣ�k�P��7���B3"�7����P;�,���ė]��B)U/�-[����a�}�R�cZH܍16�5�/���	S(�W��v_�|�J�,�������'�d��?�8�G	��҉��̦�G����~/�|57�\�� `��S�[�\h8��Y�LI�m��E�)�sb�L���#��u�9���䟡$�l�����^�[0�X�=M2c�f�7o�uʚ:���[���v�K�F�
��nn���`<N�mjP�S��)q�� ��O2"����MQW��j�I��U���%J���	�6�oX�d����~�UN�"Jߏ�`P���SF��Ex,8Ҕ2�o�-�'z���(�D����\adY�J$k�f
��F��sg�J;��"��Y���r�g�83͢Ϋ���aX5�ZBsT_>&i^��,�0���4�{En�V�c:6��h�~_\�4������6�G�Le�L����j=����>�G���9U��Ԃ�[C0uh�>kAG͡���Y$v��������A��q��g����[�¹�Cɳ�^n�9��' N�-���m�̞�c
��]���M���uԐX/�N�k&;�X��f{e������ ���4��z�N�<���ǣi5#�PbY����Q��d��p����r���G\��b����R$�Ѷo�U���8���&W,�3%q�M{�M�y��+g�zr_�V3��>9�}:���>R\�,�*K��s����*��sA�	�,Y��:��a��RrZv�ݿX�����1%��Hm��x!X��&��o螞��t	*WҖ����̣��#No�E�hJ�=P�t`^1�	�[��IB�v o���	_$~�+c���Q�ɥw5a���kAh�Y �1�p �g�̦�m?���-�'��d�����k�o\qJFԄ��1���h�,]
x��-�E>ưw%Iô� %��[,��o�NB���i-��T�\_�j!4C]�P�b��4�x�����7��Anن��׻`��xZj=�Tm�@S��0G����y71U\腝�0�.��Q�KV�� W>�c����fį_~aGn����c����IsX�u��%�o������HV����X����5�O�d��� &���)��b��-ouZk���km��x�s�s�s��&7͆����C��vs%��7�Jil$s������J�_E+՜��V�uB��`�W�8��At����;��=:�Z�-��X�.Oj��ޙ���c��3�h��)�y��f��*P�)D��?��_]�����KKA��L:�,g�N � I��0۩�m���9�UY��;I4I���O*ed�	yFGO��-{�������
�Z�S3�=WozǮ�?�m=��.�T�~�5sI��p�m��0�h2�`����3�uďi�Ê���T'�t{b,
��k��KV-Zӝ$t�>}����T%!�[�`�ν��=��ފ� �ۋ.����~w��y:]j:3*����� H2kj}�W�KДW�|��g먐��i�~��ՙq�t�YbX���P;�	��ɩ���;j]>��V\���Q��h���ҏ5��CE*���5�E�+1��X4��vq=�*}ٸNHk8�,�:(ٷI���1R��Uf���u���_Q#m�;��V4����� 凱����L�.t.�$�G{oM9nj˪����]�Wxd��8��&����+e|��m�4�cm�~NdE
���_[�xZ�4}�췜ǁ�E��F�Ic�Gy(M�L�����1nb�x� ED��EQ%�=D'�G����WT��Ա�����{p'����J�Û~��ض��V	��TPL�e� ��p�*)O�ς��z�a��Tcœ�}dK|��3m��h�]�fGa阩����yI�R�_T���Q�[��6�q������*'��GY�<+���b���D��L�UmȠ�S���iG����!�UfKD��a�hG�Df�Ux�D|�ɹ�O z�{��}�	�I�cם�C�}J_�Du�P�
n�?���N�}B�&�|o�iyS��H���	B�Y�%P�����7M�%�%��od�P��`>��g1������Z��>	�%*b\��>�p%�*��(�i��!ABQXrv-u�nxv�Nxc!A�%�s�t�J�3��1m/w��a��*����!{Ј�G�/ yQnK>'w"FT!�\���ժe!P ~IƁ|lE�����i���9���+\f����Er0��9�ȯ�U=6Wc��Ě�|b�kc��gE��/���9�4��(�!F�L
���ime�sp�HJ* P��f^A�� ^�(Ր��ڽ��a��<wt�m�?���ˤ��o�����i���I6P"��t�����1{m���&�I���}}�mธ��"ٺj��`XI2���Mh�x�Zp�d���@E ׼%��O9	|%Jf9�A�omeG �Y��^&9�/�5�T������\t���а�`���q��Z�U��.P��i��&�����,8�#2���_F�kڪP��$Jb����_�]�tA�Jk�&h��fS6P<�r"�9�M��n�4�tԬ��~��9��dh�F� �C��C<�,G��}1�GI�ɧ�ҺD�{�fxwGT	��H7ws�}�GB�V*�d���*���*STlI�@�il��_`{��V�ú3����e[�ſ����uo7A�&5:�����紑��H�"��Ĕ�`)�x3$�PK���"�2pE2S��d�����E���O^��mAѴ������v����\� y�jR�2��k���D���h!_ت3}H��G�d���險�`���y�M���$��Ub]�2|f��A���U���v�8���xγD1�ȩ-�@_���k�^ H�Z���yd��i�;L&dōo�ֹ�Z�C�,��+2�wB�w�����;��X���ݓ'_�S&�(����\n�:����4��R~1�����*�˾I��d$\1
w����`���ė�'��<�GA@��0��cq��^�cB�Q����<tOG9�G�lsk���bP�oO=tK�3���j(�؞3?>ݼ'-f�
�`\@+�i3�|H�z��#/��Y�q�!i,L��\�%�թ����I�{ZA3*���N¯o�M� �@���)��(�(nB�c$�	�w|ɓ^��7��H6+m&E��Qa1 	s���k���g)���Ur�p�Wa�w�D;�B�<���08�X4$H����I��hhOK�%5��/��I25'�]��)GQ�r|II߼�����5U$̿�O����UA-�\���Ǫ�1�� l{�(#�:�-1z�������HqI��1V�/���Ng������M�����`B��*Kg	�X�����P����z����Vtb����j��P{ð*Z�X ���/�\�ԏvh�7�Ip���P�(0[P<\ڸ�npb�ߊ@̇��Nc�&�a��Y��NM���Vq=�k�d�ul��6B� �B�~HA��0K(OZ�|�taQ�y(�xn�;��`tp�S�b��/�T|��;eQ��Vĳf��I�ޔ��6;X�����v����$i�|���t��O�Q�4V���1�9�r�a �1q�k��}6;�$��'�vjE0~��г�Ϻ��Iډ��[��{�5�N{x4*��դdH��A��6b�H��p4��,�מ3���ó�Wښ7/�3��&|o��)�x���}R�^g�tM��b��62�$��&��v C/x+vL�xh�N�#�~��o���[�{@$PNZu�6��E���S�,c���Sc;C��b_�P�cd�	|�A?���D��?���7l/�y%�(D԰aR-4�YJ�����,YĝΥZ�Z[�FN�e9�V�Z|�amۨ��#[#��y| �p߆z�b��&	&G�wo�Cnr(�Ƨ;@���GdcO��2�ş=$�r�m��
s�J?�ȴ��w>A�If(�!��Q�<��h����R`P�	�V�ń2�7��G�I7�	H����TT&{+/Z�<&��y��#1Yo���Z��	X@_(�=:�-���Q��A��m �G�7qR����{�;���e��Bqڡٚ@�L�>�+��z�U8�.����iLp}�A�ff���;ޔj�]�K�y�2����)�����ѷ��i0��������w���Y�����/LE��1���B1�~�g��{R�c�;9�r9d�X�h¯��Q�,�y0�1-�*�_R\����)�i�r�'�-)��ʘ?��C��̼?MF�.�O弡MȢ�>U%���WK:�X��l�"A�q����h��̧N�� ˳�O�+O`[L�`�W�WZ�4��sU����`M<�Ϊ/�y r��#�k�@}��:M�.S�Y���8��R�x ���F-�y�1)l�,�a�q$P�@gd�t/j�Ax;"���F]ݗ�F<,��Ḹ.�i�H�ނ�q�x�""��*L܇!�U�!�o�}�z��Ǵ�$�:=�L1�*%��䃘R�,��e�T!�,�� F�7�����̄��ӴĹ�C �h�4<�)=�y7/��X��b�w�:5l�?#Yma4{kIl�\���זoT�жۓ}
n��N�TŔ��]�	�ᕞ��G��Bx��ަm�H����I���>Iӭ�Y�)�&珢��`���;�b���J��#�?����߫���i�:����L7������_��	T(ZK��;X���
���~v1W��9߉m������j�&4O2ٜ���4�??�SU�R�n8q8�Ӕ����F���'	T��t�q���!х�Qụ�l�u�lhu��?���ۻ���cM?�/�u�j��a��-�e,h�0ι�w��{#9x޵Vř���VI������F)��E�rc��Љ_�r��l�Վ�Y�2����v0~��s�9�\������Xh7�+I�)����-Ɖ�X�ޗ9���ywê/>����vz=9'l
1��U�ݢ�`~�Ə���6�G�˖�藹������*����*��(�d�F  ��F�m���u�ޖ.7bV�S�;H+׈����#�@@��������ỗ4�$S!�a�dq��]B�		w��z]$H��Ҏ+.�*��|�z�i�|����_�D6�D�X&XB��9�@��p5����sɥcJ�rC�H��]
ܿ�|M!�|Ϫv�0��րc(�QI��Å�$25(��,wb��,�����q�s>H�T�q�T~;���ĭ!!n�M�9O1�	������A�,��WuX�H�E���o��N��!�k!�q��bhrx9}�Z�̀�|�Q��T�J��@��[]~����͗�g��Z@�܈2ḿ���K��	��6-���ڬYyB��#P�P��_$�r���A����bS��0�3]WÀӳRH�0<8��'�v�Pɖ�$TzM�E�1�<	��`�&��X&OE83>�ZW�����6������ED6q���<�:�P����y�8�=��>�۩������̖۠��d��Ȋ׸���DPU�m��I(��n�N띑���7��R����'9R쫚�ҷ��X�.��b���*���X؍��_�7���p����?>¾��R�<�/̥[z��9#���*��C�����*��|q���t�cY��5���lE/n��V�1(�A��E;�(��.'/��������;ڊ���l���㼪}���S�|���I�[�̐Q��.�����S��]P�:��Q�����融�����g�O���_b����ky����K�26a�NY��nZ�+ak7q���?�T�w�$Ra�[^�� +�K�=/um��j���b�.���X�A�L$bA�6}�H���i�H��P-�����W������NE����W���:��u*կ0`��bÍ�@s��цQ},Z~�r+���y��#�0�V��!w�/Q����!��ړn��=ДϪ������ɵJ,�G���r<�U��7)̛�Fc��(�Lg��qh�"Y�1�[=P����e������dC��z��<�s@���U�{��8ҝ��Q-!?�F�q���*/���̣������ȍ{�q���Y1e��ki���a��.&eJ-�X�%Z��B�L�D��W����|�s퉽��Q�n�?��u��џ�+�����T��͇I�c�C��E�
/��v���R��Lk���
<��=5��^�7a ���`���qU���$7�-�v����.��p9�O֛n�;-G�����6��m>	����Q�U������b�W5��)��� h��T@Ɩ�h�B���>�w��'s�3緭E���c��d|��bEW�K�m��wj�su�
G��z�X^�횮K����B$*x��q_���7�ɤ�|]n��H��_U�����a#��9'���/
@e�
�����b�  b�WN#TE�Y����"������]��M�Ҏ%�F���.AW6\-x�C�.=��ǨA��=���mP� ]��ng��NP� P��HܴV�lGIa���O��t��uw�Xք���X$mu�{�-u�_����0*+7*�%�jX�J�=��%O�Fw�.Y�)��Q��L�ܕ:,}�aU+��+_9�֤X}��v�@�tH��)b�z�E~�t��E�]
��^�H³>9�e3��b�<а�-�� �s#]���Q �U�^0�I}��T0��]�����N�ψc`Z�l�eb�2�Z݃�*���&�����;�;���x����:���r�e�'IZںF�o0O�Z�����Q�Ջ���g��^Ce�GCm�l=&���䃣�[2H�����"����2�tB]#a���lFx�ɜg}�i���/��8;�E�^Ǫm���Y/���#5�,)���_�Fj��}���[յXa:"v���6���<^��}��>]]&>�ې���OH�]��0�ICf����|3��9"j�4��S��b���M�Kx�K�`r+o��:HN�?w� �1���$�=ɑ�#]�zw�,fF�L�kp91������5�w.C:��8#x���=��� �����Q<"�J�	���j=��b���ޱ~�V�r(t��_z��YK4�R�_쳟O�ω"�![�v_�Ly�Z����5��9̰�W�伂�4.�3� �S��Bq����K'd����%��FӾX��{E�{3e���d�r"�!.౬0�n?���:<�l��R��p*�Q�͟��P����V.E?/50�ֺ�W�>�u�5,����J^�m#�X�\���Y�����a��E���YX$�K�wE]��U
�7Qt��,yQ����,��R�|D~ӛk��Vhd9��Ј9���zٜm�E��D� O��|���;�BG٪�޽�~�v��>j���(�a-^_S Λ�^h{[�o̑b����=*ߡZv�3i�!������7�dj���a�4kll�����H/���MLu�Ib-)VCH���֔=�c&&�>z~y����+�5���7�ۺʙ��R�{:CO�^U�a�����N;�C��\@}�@���Q���C�΀E͘�
(| ,^��@MӀ�b�e��/��썠�4��3}��ؤ��a�A||UQ�u=v.>�;T����n��c�q��/���~��S������ ;��"iVӂg{�,7�: ʈn��7�o���d�-�I��M������{A���LEFIE�|��:FY�A��5�LWi�P���-<V]�ǖR��[��l=��06��ZϪɼW^�CFh�i1馴{/��aL@��c�������YR�:9�7��Nk�F2];��-�t�gDHʬD�e�4�b��@mJY1-�@7�#ĳl�\t���>P�)R����i~\L0�E|q@�e�h*�ke���~�d�ӝNK�'��ꀁ��7��,d�b��{��y���C*>h�LË�Y�K֝�wU8�A=	9X���������_�,��!�^4k�*��4a,DBrW��#hƌ���T.�%��&����&��oѣ�L����-n ]w�Z �V�S�ܩ���!S�ɂ�����*ج7�����*��{�k�B�2#JnӍ&�ӑl�[�Ŧ�oj ��:����I���_)����@R�5m$�|���"���e��a�=)A�)b����:��[k��N�ɚ�!L�T���)g���'�+"�̛>?��h���f�0Xwҭ[��-C9�bv"�K��c��C*>�eߵ���A�$� `.��;�upk:1��_���,�IfDz2��>Z`�[�5����e�O�����a�NC���*-�t�@�� Q�f%�뿥�_5������#Y��,=�NN�DS.�2��c5j��X
w�z�U�Pڤ���~�#%���MG0MP=2���2*K�-��sm�I�u�,�v
�m���$>Fܬ��*�gl�E!�c0�S���F��$�hZ�85�)T��n2������*/!���k~:��,�-�d�#@�pH�6J��3�z��^�\�n��������
�oh n�����z%d�wB�9��h�+�6 �|ϞB��K��}yu�l�B��z;�h=��Wy�[+��2A��$U��w�X$6��ޑ�������YԼ&Y��\V�6e���S���moO��ky���2e�OV�f7A2|�Q!(כם�ڑR(!`V6��d�S�r�~�Pc��y�(�7���U�n�]r���Jp�������l���0ʅ����|i
��Z���������T&D�-�sy �E[����&
�[J��r&0�	�����jO�K���͜������}��;���P���lg3#���+�����xJs��5�d�	�^|�����@V8�i�X�����7fҶ��~�,7E�ly[��|���N��zM<�Ʃ�H#rw���*<"bz����!��	�8|�\�g�3�$��{�����CZmF� �v����Dy��s����cY�.mر�����#}L�!4� e��q�.L��MK����3JR��&Ȉq��ni����6�����1���ed .�'h���_,�>��.z���أ��[�E��Z4kޒ�Ӌ�Ts'$!W�=ä.�kL�= kJf�ڋ}�3��}k*?a�?�v��RUv�Ћ5��`�t6`�T>R�;5�Ɨ��GS�[V���nv�-:�˚�e1���0�r#+�J!U�X�����F|����2�Bb�>�&Bl�;nK�{}e�x�;����*x�?U+�_���;q�M�_qU!r�;� n�����]�?u�+2��x���h�΁���un�|��FXϸ��H	^,��Z'G4��|��`��p��q=t��Æب!�e��l��Z���������K��6�!D�����\�	�<Szös�`���a��~菭 L��L�����z5��?S2}$�CwC{�x`�@�]�=��4�v�	
�7'Έ�l%s��lDf������ݠ�/~��r�OJ$�c2��|�_g��"��v����4��-5���4�~�W}��}��O�兩A�PW֐���ᑸ���1
��6��ؿ3�89`z�e=H��x6�@n�|�V�LpJ��6�D�ҍx�S��6�|� �s;�뺕��B���؞q5�$��s�����?�:GQh��!x�̌t6t�EB
Q>l�'C�EN&�g?e	��{rJ��4R'WL��M	n/�K��p!��ts ��ԏ���k��@�$��:�b�b�=�KK����'�����ik5y3	��5��h,��i�N�Lw̅*���*}�KIm����xk���R(�i���29����y�����f `�;6w3w�m��o��zmύȍ�^";�:u���vb�}\�N��*6)�~H`�@H޿Y!�q-.B�׳�v��=�{/RRr�,)�攔XW�D��v ���>��	ɫ�-��;�EC�ѿ����]pO]�(�����ika5�mу��P	��8�������0 ̹�Ů�Q�;S_���p�]��KJ�g(1�)� p6Q�o|�&����nv<�y kK�FV�ԗf ��,���I��~k/J.����k}�xT;��<��G{z�Ĉp��nt�=���kP��ί�I#>�e��2|�@�zk�^��?���n�(Q�0u}=嘺Q�N�r��
�)E�3�F����r��+�ha�V:X|��OS^���0��)��K^��T�������O���z#o7��w�MA{��/<{j�'F��fF��%D���o�MC��	�Vd"�,S�ٛǿ����!����N�x�v���RN��t~�1����,#"|��u���}�C����
�tWm�7��SHU�d^xR�r(���WtY�A��Q�op�oΈ�BJ�t�Jm��%J$�T{iQ��)�_1g�̛��'��jE>����J �\X�-R�A�H�j,WPyc$��� <H��4��%:H@[Λ�/N���$�ְ���2	Oϖ��?�)�m�!�4Td���Y$�1�yt�E?�u=n�xl��9��K����T��k�V�]`����Ub�$uo_��|w�K�m��5��ME��!����0��ZF:Ns�#'�Y�-�Mem��`aKu��A�����^,����,����V<����I��R,W�ڮ�S#(�*�b��qO^ߟ����Cef�λ�	.)C��P'�x�&D����A�6���Q�R���E�z��<����{���}�;F�o-����t;����3��<���Z�-�Y�A+�O/�H��;��%�%�e�uc�_�eF��(EN�Y��^��՚2̒�����/��ĺ��.��k�$V�h&��~�V2�ȝ���܂�qI�Ky�*+A��1�7��u��Aƣx���.b�vDxLQ�!`�st�R�+]4yĽ��>G��1���ދh؜��ѣ�ݛ����e�$�#�ܭp/����
��������8]v�<�����C���E\�T=,<L��2��7zX�Ԇ�J���2QP�^�3�$�t�T��P�0(���V!!T�PW��P�k6�D��śӱq#�d��)P��l�ʟh��賹C'̧�-{�c}FX�f�D?�J�ZE�4y
q�@2���|`��c��i�U<�n�_�Ow�b|� ���>��[4���D`�3����_yў�m�4���nV���C�Ȟޓ�%9��j<&��
��7�c�;TQBe��ǭ��X��_��:�����77t���)Y�����f�>���P�h��.L\�a E8��