��/  S����3�c�ub��_NЀP���t�,ï�!U;�P{�g��Oj*�x �*�'|�N�Q]/]�X���,�D��Z�ps�W����H�P��Α���YďOx����C*v0?�t,&O[�'�~���ۓ�qL��Yhf6��i����n��T~��߶�+̄�q�U��F��$?�A�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�PZo��Ե(��殆Ȇ5K�si&�z��eR3��������Z3��5ņ�X-�yC����y��4J��?,%�i��YӤ7�$�۞$7I5)8�h(tZj}�������.Zꊜ�G�g�M��u����!�0��OK]�v�YA�Q�u�0'�w��+�"��(�u�?�o3m������B�j��3Wz���%�R�̤ʹ���~m�J��'��{��>0���O��I���H�q��ń9I�-��E4�˙3s�c�gћ��^�S��>G(�7��L1����P�o&}�T%y�0�٨'�H���<X�*3��|����_4���!f�*�d8��*ai���������䛾����%f��.M�e��^��4t�=�]���ql�w�sdS�^��<���u#tLΨF||�+Zz�}o������'��*��n0�vTXB��^��;4Eh�sfXb�shN���,���T�D�)(��4���pM:�>�������V���(�o�K�r�7=�S+zE��#\�jEtƻ�vh���`M54K
�]Ǡ�-�;���#ܾ��n�`|�:[&S6)`σ)g9Y�o޵�_���F��P
�E�샋P�Lz��<�Bu��J�Vy���+�׾D9�P ?��A�m�"+���aVJ���kɁ���
R	K�3&Ɵ��#��� �	�{�%I銙�jw��ѥcRΦl!��f�+2T��A�IO���.N���^����j��>�����@g�Pu�j��jc\uN����ƥX	Ϥ"F}�l�gنiYkc�Fd�d�c/-��㞪�˙�4�Hi�2���R���{z̚�{���TSg�Y��bDQva�^μD%��Yz�%�uvg�t&R"���lI�(rC��`L����ix�����3� ����=��n��f섮�T�*���*1��"*Ւ��(c�F�^/Py1��S*���!w�/��!�2���8"���y�՛�uyS�#�#;}귰,f ���Xϛ��4m{�J�bt�f6�u5Ѵ*�PO3�����O�*)�VA�B��i�;�������y���k�	�0��%�L�`� ��c���F�*᫯���]��А��!|��k�(ş՝0���lo|���!�H���/�`��7^*:F2n��/�
�˺U6X:��[��s����7�s��f�'����ФV�ʙK�L��՘��.�u��]{X�����k,;���kA������F����߭��g�O��g)�.Ed,Y��l
m��oH
��R�r��1/R%�w�9�x�y�pB4��Vʘ/��!1���ҿ]]�9 ��S�K�D��^�D�r���q�r�x���J��2�Ȯ�+G?�5�cş5��G�;�U��3
W��S� �S����5�����}TX�wV771�jj��4�X[�	]� ]C�v�{b��.���I,*f1�Ҡ�8K��X�	�>^8��^v=�8���� �21�����!]�ָ<82�t�c�\����k��k���}�p�,
_��BgZ	���虚n�!��'`��=��d4�܉NN�o��d'����z�W�@Ǉ2��0���k��D��L����}���[���>�[ǣ���r߆��(^H?�Cѫ�F���낪��t�j�|!�TES���6Ga|�K�a(h���i}�t��?�m<�'ǆ%�5#��9�n�����9A%�������}��k��<��v�с�ڨ/{���鈈�q��)	�B����!$�7>U�5�s�l.2��ߵ
6܀���şJ��;Cm�v��L�5�̈́-�ʛ���-0PS�"Pi^s��"H�v�0��)Q��ۥ�\~@��Oc��!c�a<��
�N�R@���M�	�aSUf���M��jF �9����
�)Խ�l�r\�s�w��R��U\���Sڐ��>ȡ��k�ƓJ�-z������i_���*�לT�c�U�'�=��7���7t ��R3Y���/B,F������*K�r���rc��h"�4���Y���������d"�bu�S-/���Y��
2˓�YWH��{��4b@�J��ja�j���i���{������x����j����0�	�����a��k��t/�	~sY��:��o�<D���ɵ���H6�Y7�<]^3���������F��k���ٱ�i�f�3�p����~&�&��yʦn�"l+��p^�Iߊk0TȊfZQ���7<�qҰ F��Zu��)�L��}X	w� ���i�VmK��B~�Y�2�uc�����c���i� �a�K?ǥ2_�F�btT?�i~뽖kwF�Ԝ3�_?����o�_��I2p`���$�٥;.�i&>�G����s&gdT����Ç2*����>¥�K��i�!N��Md���
=5Rr�=;U��"���q�˪�~J�����_�M*��x������$;pC	VH�9�=�(������
���s���~�V=����y�7��/I+�O�k��S��֟��O	�k�~��]��F��\g`n�O��s���$DVҔ^{��4xA�n(R�2�v{��,�̿,�	�5�<�n����dޒ��x���������p�bs%�rݭ���Q�Lm�!�"�W�F h������|�����������(��?�Z�DW�Pg�U(�@� ��b\�O�gYO�^y_1���������p�RT�ڊF��T7�����gz[�-��,%��v�� 
��u�FLK� �8�Eep��]tr���[m����h�8�8��ΉnB>n8>��@Zc�D<̄--���&^��#��Jٲ1��b�+�0�&T��3��	4���}-9�(��%Ƌ�:�mP�J���h���L�*VUD7�s�YK�[<Իa�{)���*h��&a{
��1��O�v� ���v`����I*����(�wk��ބS9����|��`	�W�\#�Vv��9�?s� ҉��]z���g�3��v
��$,��/�J�w��yT�B����X����W���$��s��y�6H�f��n[���vY���@�'��#��V�W����P0zvGl�aƭO��V?&	���)���K��J��L�j�7�1�]����tq�!K�����Y��gn]��W�&[���v�l���wc:�������*�ĭ�7�ul�'��W�M J��e�����Q_m��I��R3�73qi��ԽjiGC��Z�>��/	�X'�Fi�?B.���V���%K�#�N��Q��^���wdy�eOY5K����dǭryiƀ��a��X|�-�-eww�խ�O6���Ǆ���^^�e�
~?���������m6|�!ǝ�%��.<�\�5 ]�ONP�6)��=���
=�bv���<>.Ux�k�Hy��<2Q�WpPj�]���������B脶����,���j�;v4�ݐ#�>���s����WД��\�57:L&�gy6tɍ���r���}Z���iD	�Cp�ٜ�7����x8K��`$�,lp]�<}�=�Q��SR� $(��`V'2A�GCj����CB����WG&��8�#y��9���h�BD�����faN�.F�,�k
/��4Mش����T-i� ʇ󀃠o��e��o3Kl�@�����@b���Sh��(ʐ�P�!�b�^���My.w%�*��ܵ;D-�7��8�y���I台�vM���<�<��x�e�{�_�4��u��|h�|�x"��t}�9IX{Tʥ?e,�O�^#|�x���]�8�Ď~m��P�G�G]^�}���A��^c,�점O}�F� �Q�D/��L����c�^׸sQ<)��)��?x���HЌ<���;U��� �T����$zS*���:w9�ù8w�Ԟ��̀�J�8߈n&e4*�B'��ZP'廳Ž�"՟d�"ŵ����5�B|rfp��&v	�Ԙ1h�.��lr�v��Z�Q�S�����b�d�E2�����yI̷����2�����c�AfT����c�]ߟ,y63^�V6��MC��#o>�k�<s�J�4��<��f�ܱ���v��˸��@�=��軲Y�&�D�n�9MKX�0a�.��1K��Ξ��_�C�V?%�soɿmqE���)E��5��+f�5�%�U�u 3BԢͨ�>P�'t_ l3�{2�)bRzc�� 7�z�NG�b�_O��n���wԳ�I��Z���~;"��2=�ψ�(iIg�`�&�95m�H�<Fw�F&Q���m
ah�M����b�&����tI�5�}Թ���h�nd�{��Do����P����t}a�����<�&s�`����j���!w6�ݬU"�J�'���&B\���WxmZL_r�G�
.�����2��t���Ӥ-V����=J�&�Pa�����W�Ԣ�5��H����^�2&c�qd<S�����6j~�t�7��n-r��!�Qs��$y�t�H���RM~�N$GF����+U�dN䭑"�}��J��LDY��_]���н�V{�NۚMT��P���F�v���0��m]t;�p")T�"s��#wV�-��(oU������	����ꭱ;�	�N.�ԃ}�YRa��9P�����u=���#����zʑ�D:���Ė;�ڤ��3�0^Aø��֜^f����ˎv��ԑ/0�R�qЩY��� ��D�Y�[�8{���`����`�o�Q�C�j,o&1N{Ԗ�M��B�(qw�fD,�ߟe��K� ��B�c	�i��E#E���A@+� �7g�,��j&iQ����_���FD6wj��E6�>jt��9�5��ZmQCrc��^�4'hOD�p�[���-vb|��E�,��q���dO���N�7j��D?�,(��"�*W������h�~��&h���()6�m�����O���b��<c�J�V�)�[��:Y����o���[[u�Ї���N>�&;����$�ޥ�р��|z!�Z��/� ,�Ad
k�PxS��.�=<y%6�1�1bE=+��R^�;� �}k�"�*��y/����_(K�"w; >@?iS��`דo��<}�~�|�7���(���k�.�<Ѷ#�"b,�� �R��;*�_԰�->z��k^>���c4�^�:�xAu���uoIu�3�B�)�%v("��߶�̎�b	ƾ(�y�K|�x�
1&��m����b��mY���+�G� d[<��]��G����H���'ഏ��[&"8����O1�17�k��3U$����2�U�b��AH�N�U�{i���[��y(ԋ���'� �wX���K	����|j�y����3/ι��-)�Y�ίg�J���E����X��b2�}�}�e4�_F)Q$q���^��yv���"�"zD�B�Dp:}���w6��(B��3¯u�Tu��{�/:��a���b�E;�o��K��隖Su��&�la����f'�;A��\I3{=�f��F��.�WV��,
�S��(��Whm0�p�)���5�"؛f������D ��U�_�z����C�3�A����=F��C��*Yh��'�B�bH������)B�j�����K�O�[5�t��@�z���\ ��9jcq���rf��`���*Lq]0ʑ3Ϧ��L��2�oUН�DȑK���~03��x����dbD���-�Y�.�Jy�j"���' p�=	L�?��uo����-ܱ�M��,J5m�˽�,����`��y�4�,���3B6�I��IŀZ����9��'G�ۿ��%�E>��Qs[>���fź��	�Y<�(����3$Ɇ���:���� b\��0�P�2l�]�ޞ�����rt#ĳ�{��ے�x����˱�H�!�S?)�5[���O&#Kơ�O�PI���!|h�2��7Y�M�k�/Q�Wv��(R��d$��T7zF��_c�kEc���~������a蟔oVY fk(�� *}�b�I%ƭ)��Ԓ���IW	L�&Vi��D�6�0rԓ��*���Q�4�o�;��"��5�0��#B��4xfO�=0e.���绉���j�I
�4�e���6�Zx8Z.j`�Q�k��j%��4lc�ϩQejd)Q4O�
��)lؐ�w��t����c�A&Ks!���ǈj�S}л�eb����s����\9,���W����mx�}�h�i��IB�Do���c"#E_^WPL�:��%�W�lYs�^VE��n��: ��o�Bώ*W�6��BŶJ>��t�7����|�Dy���x�ukY�vM[b��N�$�<t4�&��I>B[����Ǿ'��LJUv�����d�s�V���S�NbS%Y����B���7Y���`��{ɫG��\!Q:~�f�l�aջ�u���I5��o2C���#�L_��R�-G�D�XS�"�l� ��.Dy�-Y,��'�h��EA��\�4��3�KM�y;��-a?J������Դy��_����a'6�VۃL;�v)n��׽`�۰ �vv��4"�0�ӡ,\dl- ?�Y`a�es���*5�t��Q��ڱ����h�yҬ�/xW��Ի�E�yc>�0�c�
�R�k��+��wN@ʶw;ʧxP"�<�8��$A�`[��j���:7����T��m`GXh��.�v�Z��Ǐ�.��ó���r��+�Ⱦv�y/�1d�ɜ�"�n�S�}�fa�Q�������Wlתi��YyE<$Fkv�j���c��sL�4!9O-&Vz���ռ{��b�t,~p���]@����&��yJZ��ț.���Q��Əl埭w	�>G���,,z�vg:X��PdV
n���>S
� 3*������^��p��0�)j���|�#�9MLv���ʃ�:�D����<�N�!�e�rj�1����M�e��?v�>3RܺQm�13T�̙�w�<5�0u�f��~z�0+'gC�����Z�
	-��J �U�� ��Ƀ-�����v0rk�?M�S:��`S�eY ���(��qN�g;y��C��)�e����O%Ao��*��v��������9��#��:/�b��T\]��Sw���GJ�a���xSt�����!~:}���L�O9�@�=�4g|@��'��O�B���8���p:����y�}��->s+/ټg��N�j-�F��	�4~�#��_���ʵ_R�:xg����y�7��A�S���-f�Z�ut]�j\<Τ8�Sä� r�ФT��	<�Bt�QTHy��d0�>�]��:��{�j�E%�'j��I��$+yڙx?bUr�=�������UҘ�����šA�:�B)����[�K���
츽(T���ϑ#&�Y���Pp�A�A/z�~u��Lb�ֻ2B(��uP��h*޸�UpN���d=w�2����s���q�K���)�xֽ���_��`���,�/ݽ*R�@�c�U��Ҽ	�JR��yq^M��b�S�wFe�OR�� ��8��s�������U��4�vS2�9L��YW@jA����.�W��q�vؒ��E:����)B�+ѼK���Ğ���ǋ�Tn��,���xV6��$셩���t�w�k\��¥膳�����[<m����n�MW�=I��{1?E䉆"[ާR �!#J�^(w��Ljt�y�]���3e���������CoV��E���͡���w5�����zcC����ᒭ����Ҹ71�ܛ�ր�xݚX��[DɁeV$WK�7��q�鳣z��g�:�K���xZ"�tt��RE7sF�,�?��|5,�𸠒XB%�MY�]�.�}n]R��B8�1��f	��۰�#�S*d�U';B4���KA���~-��9����t���1ե5q�U�`>�`�� Op,�~�2�![��e �Z���^Y4Y����(d��١�lB!��q�S�л$q�T9ɭ��eUh	���؃g_��� MeǰzC�7��)��B�
�E`lL!p-&s�foeֆؖ�b�.U��a�^(u(�A��z���(��1�m���Yl�L�i
��̥
Z�9q�U�uttT�64��+�cC�9��O��"�,���k�����Q(���:�M�,��j��
FB]�'���M$��c�.�=㎞m��']��VP�����	6��M�1N
�k�X�a7���MC��ODf���ɓ?�6�|Ⱟz/�z	~�
�%2셁4Ֆ�J�$"�9Z���>Ӊ��#��ap�	�f�j��rf��9&h��Y���˃�r���6)�"%��z��N�v�9���r�Ɏt���{̾�[��<b+��>�k{�x��=���HX�h����й�a�S�{��Z��I.7]���I9�J����m�o
�pr�ѥ���`���q���C�呂�:a]���pzO�h�+�H��؇ʁ�8+�_��rdW:�p 5#ާ�o�m�n"�|h�F�]q<�@Ak���G���*]�]d,~0�A��('��ku��Ù/��`-T��0��V�1��C������J���[1U��K�	���!m�ÜE]	���p������5Ơ:�Җ�p�ʘ�L��VRiߠ��/��n�g0�PF���Ď��P�����i��eB�5��T5�e��W���mjè��]�+��J��>U���h���)gd���e�!��ɖ��^��b	�j�t�P����DWM6��"���z0�Z������m� �{��\0�-�|H4�����0&���p����x@y!�a�ا�Q�8ey�;��1�Ԁc�8�JT��á��.�/�d�.n��A�/����;W�TXL.������/��m�l>)١0D�1S���b�9o����x��h�2�!\��kA����YN���v�d��xkv���"��7��9�����iIt�i��H���{�� ���Pw����^ٽ�p���^���o�n-)	�2���U�Az�Kר������<����uF��~��G^S���Uw��$��p��p��n]!|��Xyi,fL���	c���)q�w�1�)���},:ͪ��om���J�%��<��s���&N���}��S����l�篟�yks��tnD����}�I���F�]������.̣�ޝ��o_
\�,SM��К���|�� �j`g�^�&&��V�YoPEu�H{n��1C$4[�NZ���#*Кp����g��å��DZ�x���~/�wC�;�:�P��f��?g���l�3./oߕ�R`�mQ��ʖ�g�3�V���w֡�H���Ct>{�I^Q��xOk����1K�V�ǵ&\��l��nф?��O��ƿ� �12���%�.�{�%���������YPހ,L8�6�S0�-*VX5�p�[4��a0Qۄ@1Ɔ~�ʓ��A�T{�dE>�����X���s2�2?U�:����6�aK��[�|���ǖ�^A�s�R����Sq)��S`#���>�D^����N)H��H���ډR����~��
c�.b��|�F $²M���k��`���6$:�]'��{-��zxL��~���=���˻�Á�}/�����r��gQ����#Q;	�\��Me�[it�
S� ����Ƽ��u����:=��Knw��j��9\/����6,{���u]'y)�6��$|�x�)�$�;���U;P��9?i�1�f�F�:���}(�Lp�������R𹤥�q ַ�-B2�bV�����15�]~3�S���P����M�����mu�`�������\G��w
L��ƜGx�R�=�� �)�fd���ag�z�Em%t8�
٬�P��"�I���+H�M�^K�@<���1��|\%�c�E�s7vurc��5_��ȶ�'܃�#�9�K��;\M"k���*�� �pC�Y��BѪC{�u��4,ކ^��
���������V
z
��i��ڛ��R"	�DmNM�Μ\fK �ҿ�yW���s���&�/񞎖�Y��Ar��d@~?,��X�����CҤv���)o �����zB�ļ�rBWq}�{�K�f�������JE�
�Q���r:�:�J�-�!��Yn�z_l��[ʌA���e;�9&���f�	@��!i���m>TaV�ZlC{f��L?�~�
1�9�ݾ�Hy~�К�0̑l���ыCy�\����������H���\]���;�1�3@ˈTG	w��?���m��a�F�m�V����.�w�C�+����_Y5�$���]{&��[�$��a���7����z5�\�~�z� �R v  4HB���M|�G�K��g����*��ٱ�P�0���R�p��O���Z[&����Ax՗~]֔NQ�O�!�N��}P���~ۗ*��Щ����Y-��=_�K�Y�9g��u�o���/��*;ā�����:Ӥ
~Li��6��i��=�P�������j��2�` `���i7�ο���Ƌ�C=!��v'����������u�F04L�����o��ow
Ib��" �hRM���~��fO.'W��ø�ea��8���>��^��B�\��ܪY;�|P�2ϡv�<�'�����;��*�qE'��*�2חh��А�!]%r�Ei���66�~�XFЯ�e�X�LO�L�8Ӆ)�4����b4���1�;��Y�h�а���#]����t�]��)���,�{�P~4a2���)@F���Y�iN�ڛ��V���(��w2�14�-�
HP6~�ցq	?�p�`a��m�G��PH�gƲ�#�&D00fJ��rF�K?^���5����d�j�C��Ά��y��hԣ/��P}��@0���,Nߟޕ�Qd�l�7&@�b4v�)`"�}���z�,s�iTA��
�j.Q�[	N��8�䉀w�쓭�s'��u��mT�g��;e�s �E�]���_>8�6lJc�td
Kr'����p�CQ�sh3��k��V�N�c���8��Q��lg�f�F��;������Z�V�L��ӞF\�Z�C7���5#N�2I�`�V"@������kp���q[ ���v֊��Hb�	B���x���~<��	���e===�Mʞ'ƀ/�"��&�^��mr9��!v��:�;��r�b�]����~l)�RD�Wk��?{8��J�D�D�ZִNH��\�(o{�y�^��4�x4�7k1�m�ݪ��5�x{�����bzjL��1�[Vy�f�sd�o-�K32�Q�ه������5�;P]9�G�k8���GR��|J�M#�|�+`
��jݭ>��rx���F_�N�E5��9��[�֛%���+ �")���]���f�F���;��e�5��4#y��h�1�RX�H�]�`��x��,_��jQ�D�������\�d�R	�K�/`E#�aE�d��	L��l��΄�i�:�����-v�z���X�.�e���E��)�Ekfm�:#�ê���Tc��l�-��m:�6���'��{�����l�s�VfQ��k�D��ߗH$�f�:����)�:�4x�\�t��s�CGZ%'\�����X�<�h�>�z�8��iqfB��{14�
0�bH{�OI��%H�Z�¦�P���~ ����OBso����l�
[��,{E�ղB���%�&̜.���U����ɟ��G�w��P8 Tj���WsVb��`� �O��4�a?�'n��IPd29�(��}�"BBh�����3�7H�Q�i���C� ���z�r!,iB�~ 7��S���k���8>S����� 7�%?�i$ zk-b��,B.S��k9�6%m��g#3!���G�n%v������1�z�fu�ʗt�Ώ�V�)�)Hcuv�Sy�V��޵��00jh�mQ�ӂ}�	��{�_�0@���7��Һ�c�Bш�-c��[x�yh�DƗ	��i%-3Z��{��N_��H�A�ݹ���P�^>��Y8Ş�Õ~wHSI���m��Oŭ���X���k^y�6F��0�ϲ�w�N[����0��z��ɻ��[f�CP�a�c��dcW?E��+͗| ��*{����7�Z�Veɦ�u�����p�^D�f�5�{c����@�{�aK�hc�̞�L�Y��1���@x,�hh���\<)����,o�l�>��K���'�(@��T��.űmp��`{<�ߥ\��HBy��s�vMHvt�N�$���8o&)���+����ԗ:؅�-�L��5j͡�1�����ya70�.i�i�wW�f)T��g��/�6$8|$�`.����om��_b܏��5���}����.���0E��ٌ!:s���7	t�4�)8ş�^\G��ɢ>�D����5�EYd=��G�\P�ȫ}���������@;i�Jm����Me��e
ܗ ��7�ξݪ��zU	�d��`��_�({ү��$?<�]%�0x�>
������g��7���?�\{��)���Ꟃ�;�*�l;k �s���lLD���HdQi�s�$2Rýc�7�T�Z%ܕ�*�����gf> [ܐ=K���Y��F�j�d)mQ@f#�V��{��h��/#���o�Q
h}T�U��&ąW��aL̍Q�4���n��n1s��+�-�p��7���p`W֡���׼ҝd�c��>7��4��;���dz�����(��ج��G2P�B�+yG�cɥԦ�F�g��m�S�db3G��T.�e�=�7�!����<�n�,�)��}�m)q�+$2�<�����FC�B�����;�%�ʮ*�~��no�L���?�U�>A^�Yoh�߹�����c�`;5w�*��B	ц�\���Q�)j	�O�]�X4��2yβ7a.���W��L��q�O�@���vG���up����O�я��f��c��k�!���L�3��s �Z�wr+�B����v���El��?+�)�]�qU�a��_*� `rJ�c���}�Xl=c�vy�7��
HƂ��7�H�k��B�[*+nc_�T��}E�}=!\F[@*������Il<�BW�t�3�	)Ӈ�c�ݙ�N��UD�6Mu�w��jrn$�{k�Vz��"���,$^�p@��M�yFem};��p�O��0#/A!�]8��ӍE�;	jϦ���@���>���>``���5l$%k��$r����$ȇ�&~P^���3�y(�=V�n����H�3��T(�����-�P\��_r���>��Ng��� ar�6���)̟^�S��#6ƻ��|&�_���-����*�汁������?�2�jIM��J���A	;�P��S�B��4h����a�꿻*��P^� V���j�_�s���H��V9H��c�߱5�'x�{�ÉP &�*֦�E,�KM�`�DM�?`�SO��8\��Η�Q�V��9�T>��~Ɂ�#ʀݙ/g��?���~j�w�`���/Q��2!R^?����dh�D�[$i< �����]6{�N]�:�l�z ��!_d��0p}B_#� �)��ec,X�c�P�ܙ�����wݲ!8X5j6�X�y��#�0�t�$�,��4U�ɴ��D�.K�|Hl7%I���Ǣ>rx��� Tؗ:"��
pY0֞I��:��crT�4��}@YĽ���=��J 8���q���cأ��n`u�ZwKcq= ~^!y:,����{����t���ꔖ��	��V�#]?�+u,kny �͐�l]6TW��j���Hܩ�تc`�{� �_��QU{4�S|�Ɔ$�]��؜���T0u�,q����=Z�ܞS�VN����{bE���!^-��ǘ��Op1�4��� �>9�6���f�s��+�*/�ҵ ң�����/4��a6��I�.���lIT�oG�Y���̽,݁Xt?) ��}�R�Q,z��=���֡j�B�j'���m&�69��(���d�Şu�ڟ��?����D��c}��p��O�f0�R�o�b�ع���9���S'���Ԅ�n�+�Gv/Ѐ�X�R���L���S��x�+Y��.���%���w1�yb	�yI�`���9٤q"SG��k~��^���p�����=�-B`����!��ͨ����t��'{[}��s9P#���r��J�fe,�|F�v�H7|.���|�&E���g���L)7�k��q�&7�f)U��E�����F��K�g1Kh����R����O}��L���ۄ/M��ȿ���-�	�JF������<�lp�H�bTiE_|����M{`�4�ү�)(�}�|T��uzn����KJ��r8ǈ��f����]1����?�v�x��6�`��Uf{�G|��5�cBNQ��7�'�X���������fb��N��֍�hU�.��Q���R���Q`	�A��X�a%��a �p0��/Wa��?X��FeR)TW%���T k�b���~��t�s�����k%C-�XLxDȷY5��Ri�c��B'^��7~(0�B���O<dHP$<�P�� �ŵ�fR��e�h@�+-��Z;��ki�K��i!����abcY)U�Y/���A�-���q���Gqvᯩ��QIxX�+�;+�Z[��W�H�Q�b�ۯ��!?6B��ݜ�HrУa��#�����	A%�I&>������K��
�X�V@���rY	���1M�T�ǝ���
B�p7Ò�e��Na��
��]oM�6'R�
�q,�'�Gg�e��b�E�}:��gk�
�RoF��^���Ok�� ��WRW�n�əY�W�g1m�L�(���=���/�V�e|%L��|�EVZ��H�^O���#I
�����A3К�'>Md�P����E5G�^j))-U�`�Щ��3V��J��H�*G��~"4��#��������d��R�<�L���[�Aj;���5N��Bf������LK�,"�q*������GE�\��l�<µ!~|�����4���|Q�kӰ���OMV��u{�n�^y��E�"�~��?����\�W��R������T��22��N���뎏��Q��;�� (�9�#����+ևk�A��DۂA�w��[,�Gx�gV�uAo�0�Uzc����1$&��3}�4_:G|���m�y�����L/�����I�I8^vȡ����9[}`
���A�ʦ.rghWF�Si�;��A7��\i���^_����"c��q�M�>��l�J&�b����?1>��n��t4>��6���~� ��%��:��
�Ws�
E���h�q�|������ ���~1��3�P�'.[�ɋ&Q\t�`���tRW�c/�Vy�(�	,Ũ�M����إ�# �����Fɝi�0����h(��%T���~����-��� S:CW'Q�i��o��@z�����Jc�R��\ �z� *B|z��� ̧朥��I�M�⑳{%�Đ�	(π�����d���G>0��Z[���b���V�o9`�;���R��b���
v��l,�.+�՘��%�QEr�5��9䆟�iO0�I��3��-x�($�c��i%'���80g���%#�L���U0��QY#I	,�B�5��ۘ2�0�ɎD_�7+xlL��Qy��B5g�>R柚Mt����؋C\�G�7�cӵ��\&h/��k��$�M&��Y����%"��X�L���t��>[��4H���a{�"��Q�Ki�������ϔL�4��_o3�������)`:�&��n���ణ/���:�t'��j�g�y�E�=��.�4vu���R=�i��@-&���/�����������E�C��&RW�M�d��ɾ��XE��%a�y���_U��-�_g��kj�(�E��R��tO=��85���P-��Wxx�v��/.�R,��"O��a��ԛ�K�:������_�xK엎ou�=4��BA׶���l�5�xˠ�Q-?6/�-C)�ۮ4��2#��O�)��*r���d^}��h;b} �ەG"����p��(��_1�-@�W���f�m�莟�K��(~׭~jM0��z2	�}�� ;��b��&Z�_�w9��L"XXX(�@��?5*�x}Q�כ�+1T
U�XWm 8m�u��o�v�W��� 	�<t8�t��&��B���ug`%!Ζ��9�Y�n�F*�f��P��&)^7AF@��2hR� �(����]1js!o���`�f����u�}��������ώ�?N�O������(`&����R��ghw6J��w�&�����vhd��H ���^jT�����D�����5��K��[��XO��PW��F/�+��Đ�+��y�HG \�a&Z�wQIX'�=�Mn�e�ƀ��4�=b<D5�ʒ���C���R�O�p�W`��¡�l�B]��a�x�	 ��w��C�b.um���Dҁ��AFzu|b�>td�PHW�'KWBE���W�ZAԨ��J���q^�ْS�%����u_ɹ��1B��8�D=�n�Y�����:)��`��50�'�|����e�*Ki��0V�"��jC�5���viq�vd��ee���@�.����`��6��m_��<>
�m֞�x<j�Z�4���'�Z춢��֨U�QZ�p��k6[��|�p��ש�2Y�)�i�S�@}��z���Q�pf�����0�{��D���H������~�
?�x��B�n��&Ѩ��X����@iQ�ʉ����2����$0)+�{��v�H�g$p��7��t��q�Ȟ��#��o4�,���?Mn�˕�Ŝd���4G~�m�t�y�T��FP����a�O#�_���Y��L�ˎ����-x�H
%����&�2��oҳ�4Hտz@��`�zt%�*��ѱ�z��әf{����.h��`����/��R���6����Q���w��ڕ� 	|[��G��Z�������`�X�OD\�?��I�H4q���׆���/��[+�7�z��}�'�����s1���.q��w����zT��c[	�Y�	]��<�m^?��MZ�p#�D-$Em��,g)<_M�$Ï�&�v�����>!��Βc;��$�1d�9��E���>��b���8�Q�<��E�Y�z4'w ��-��<�C2�U���M�q6���"�K���P�;�O�._C��յD+,-Q	��vJݔG��G�C��+�.�7�p���މF��w���N��h.�]9�0WJ��&�d�;�pނ4..#;�w��o`�A.9��|q��P�#*��3y��
C�����,�H�d$N*ӊ���L��G�F��Dk4t} �P��a*ğ�V�h3Ns90-���vjGC�\��_CwH�͘���ұ%��"�x+_�/y�f)��b܎�?�aS��j�ڕ�@Ds�5��mm��*��h7��Eu���ȭ��ԃ7���w�Н�0�y�F�r�<�?����JU:�bqȼ!b��5��y�sf��ZX�x!qTUW%I����e�$���1+p���Hc�ØW���rl0�3����S�� �,��6;<���+����|t��yǻ����ZTT������NK����*�� <�j
�O�{
ٕ�NЉEǕ���sU��ػ�/wy����:8Em���%�V��&ot��q,J�+C��q�� ��[���R"ET���7��r�$�a��nc��2���+�0:;�|��v�P����D=�,��S��[�]�����#t}*�����R3pT�h��]Q^W�m�e��L��L���E�����;�o�B�{k\O"U�S��p���.�� >߹�V!m�Cʜ��D%��X���i	�ㅯ��Oĭ���@���h�e0�����CėWj�}��8��T���g�ײG����j!W(kB�8�<�E����!W_���T?�4a]u@ITD�����R"�_�#��_]�Xdx���^!�W�Ql�d��W!���/R]�a����k<X0���F6� <����҉�˻�Ќ�VK����1�B�T$�pL��*㮠-8��������,:��u�Sg��)�ڹc�d���uI��ktv�{u�	�U�5��g���ʝB��]{�^M��bJa����c��tΏŻ&��|�p�"�^ѹB�n�=�����K*h�?�} �8A����E�59�����y1ƉA�x!�9���P�l3S>�n�|�r�&����:l��x����bV 5�G����h�(n�q-�6A��e���g�D�0�n�*t��Xo
Ӄ������F}ٚ?�5��{QAv�F�y�x��Y�fʣ�)}էgg�&����!F��bF~��\���r+C}1;=�y�)l�+�4oY�4m,=��g���E�8����G��G�K0��kR�;�і��|�t�Um���QI�wl�=ߴ��U��ˏ�1��R�ى)϶+o��O]��HD�k��c�`q��uI0�� 0ȋ�`y����i�n��r�w���V��o��7�GE>���<hm��V�T����A�C~f	������
�)�� �8F���� �[����ь����z�[��ps!Iۑi�"5��B}y��
��5�ZBd���7A���y�]=/�X������S%��`�3�#ʽl:��~�
�p��=�����#ŷ�=чNGL��}9S^i��i�e+F���~$��S�=r��Q�5�c�A��"6\l�$Y�TQ�ڟ���p�[�j������ڤ`G�j�_��D�ބ��ֹ΢��1A��yD�@��NL�,�0n�wL(O`D���l(��M�mV����d"7�XMz�����νj���K��h7��,��.������̑{~<C<�=����h������K���BM)L�׈a��z�Q�*��R��6�
ض2�d��j9,�L|��>�@r�w�Jv�`XM�◤�V�BP��j����H
p�����C@����!�ᳬ��bu��*�-xS��+��h�)b(��(N�x;���SPBFef;"섀w}�+�w��J���ߙ9smmTn�J�ۗ~8�%�3�C�F��$g�Ád��If�� Z�7"�ܱ�9K�v��k�!5�Ԯ�3�V�y`~ܩ���D<?�ÿ�ˢ�¶�T{sŀ�Ӑ���|޺,�>3����(T0�YU���G{Q� �>�a��e����7�T����{B(����A�}N��<�3�� ��֏O�.���u�[|�"��ܠ��	�ϔ����~D�����d���k�����]>xI���r�g[b��R����d�M�&DN�Ng;9�N�|���XqO���h�;m'/�SexܸH-L:��󲚸�U��X���-'5)9���h��0կ&�"Gݣ
����@X����Ą�u�F��o�e�p%w�؀�,�;-�=��C�.*^��g���G�Ͷ6?������\<�[bW�3D�.ߘ!�{�I�3*��~3�~>�"�ض���sG�r�iS�|_�N��5����c�d�i��'�`))�='���E��\��+b̋�f���@�uL���]�C&5�bA����~Rb���5^���;�Z?�w%j7_z��H\��g� 	����eeء���a�k����U��;��PA/�V3=ݷ�D%�o_R[n�|��f
T��L�)��71���QD��rsR�wsbP#-q��?��Nӄ9�H@{�g���(��ς���7�E�27�U�!l��7���9����De��f�����#ٛ��*�P���sY��r�D�t��9���G���gb���I�[lkʕZ�gq��53��@�pj�K�\���&�]Y�F2Jȿ�L/��z��׷q���v���q�*";å��\<���OE�@e��_��U�����+N!W���<��s!��::���>��B�e��rD`U5��fh4��gB���ߵ0;@�\E��v�^H���*I�NYZ��0�X���� v����6Y������tf�ԈfJ�H^��� �w.{���J5����h�@f�H7���G���p��c�&���Nz�q/��3"řV���׹���!�԰�\�=2S�l��1+t��lu�1�5ܽ� ���ɢ�w]�y�!EG��[�%xЅ? y�=��*�lܙ��5(2�̀t`�}Ep��Fc�R��W�Z�^���Z_���h���K-&� ��f��x�+Z"f��/~�v��u��j�̊���Qe�p?D�W�G2�|&m�����b���YeA=A����`������x=�RB@�(FK�knQ�����y�8�����	:���\\�&�xۚ�B���$�(oV�89EJ���e�4ަ6�>���:h�p����z��|N'������`v�*"3�E�y���٣��N�1�?R'm����o�5�3#s��Q��;6t?���2[���b���,�_� �l��@O��������H�0Pt���V�n�����#�#w�	}S󎏽��#6*o�N���P������j����u���d�A��0И�&�wҿ���Dݰ�[Va,~A䳩��Wҍ����?����lYO�p1��
�����R��k����-��!����^���e� #:�C��;z� d䮶̮(�Pe�,E�&��RK�o�H�ˬJ!��<��X|�X� �'3q^�,@O�!j�(-��O�pf'N�I�Z�,ҙ�ǄB���?�:�Η������	�8م�kH�zg�Ƨ�C�V�}���H$-z*zk.r�����I��5yq���A��{�U�cDR J���y�*H�N������X�$;K����$.�e�)�xW��Z��F�	����10���iv`����Xj>�&�;s/#��CߟS�>����c�o'����]@�^�_��(��1J/������=C>�;<DsE,/��\��υn�K/��z��g��].}�FO_�Q��g����3"�`G��@��qaɭl]�3Q_=�Z���}xցÛ�Ln��V�U�|9�vI�V"z��tԖ�N����Xd�<�7�Q���)�9��N���"��l������W�a���<Y*�4&��U"�-eS-i�]*��j��[��}l���%�X�+�
�X��є�Չ`6a�i�g\�`����(d݌jj({N��KO$�aC��Ih���p�U�Caǻ������K=���0�s���f�����# ��͌[9Sa����x=G�@~�j&vE3�2���*D��3r&�z��j�Ķ�1��;^��д><��;V�d�Mi�a�oF� ���\l.n��8����-���	�1�Z��K��$�$�v{�kb<$BYB��A)]����ؑ��` ��j����<T�5���Ex����p�7�VG��Ov��-�K�?jf������Ê䍢��x��kT>a��%��G-��%�[��֧j�r���@_�{�(�l4��pC��j|œ&����L�4J���1zw�V��i��������;�n��O�E4��4������-�z�U���/�^�)��bOUF���nk	��Һc������kMq��hbe=�p�d�>hLL��K�0��T��:����3�'�Մ�������m�Mb��B[�2�tmm�>����[`��g�(gUn�G��l�������Y���	�|���%2�2@H�g��?ς��ꅢ">�A�Ǟ��@�|�^��	�`����/�}���g��XR�b�V6�j:"��A�*���M2��t6��]��E9��޲��-���:��G�H��(mͳ�x@���E��3��O���N�*����H.�=�(�Ѻ�!W���~��ΛH��S�T$n@k�.���b���c�UG0����0�h�������͵�5Q7�2����xa�x��Q(�ƛ�k��%�O�LVQ�tq�9rxlrOc�+�-��V��F䟪�G7V�Bβ�,l~�
�V� ����;��ݏ9銨1����a��n 9x���� $!u������U��R�ÒSi1��)�����J s$M��G*Kg��C�F,�X�$tn���=#��8n�"v�Z�`�h�2]M���<dz|��G��c`�(�h��ese���ɳ歂�ӟ�+d��w~~h�� ��`#��i.��L�)!��a8귬�3��W���P<k��;����4���o�#)�td^A���^;o���^�������b/�d���7W/����{I#�
O���MM7e�_-���OIs��W��]W�T�w�r�Jp]��S���Q����N�6����~�̧~5��D�/�!ÞO~��U~
�<��=��4VX��o7��&�q�ؽ�3^� w����M����}���f�&N|����Z��K��G�=���5l�xf�.B!J:���.ľ����"S���F
�0� �sһq=bR�K��+��X&����H ��}M/��J���т��+G�Ȳ߯Y��+6drҝc��Ea�G~R^n��}Ua��sp��X���W�.	Q{�SW�K4Ŭ{�1SW�}��j-C��Su��D5��� ������[6y���E�(��%�
�yH@5�مx�=}��e>#s�Gr�^���7eӯ���a<r����Z_�;���NW��^L�,DZ��c�d�3����2���ȧhO��߶��'Z���{2#$��	�L�3�$�K���������R����(��K������f;�	S�m�6U56K��>D�����q��<�#j�_fJ��VZ�S��m�-�o��j��ǅq�w^��F&�z�� ���0�_ʫ�H�o��(Uu��"}�SW%��[Q��e�b��U�E"Ǚ�ƈ�����m�1¢U�C�3	�i�*����O@/�I��us��Y�u����r��颀؁���&�HJ��(F�_����C����6��b?r�C�b��t��N2��3�R��������.(�?��/���zc���>��:,�W� ��@�<1��36Jf+
u�
E�C���ⲟ�]�	w�Ruˮ�7�ִ��I[��� �ы�`�Hw5�:i��D��UB� ����4���:��Rrf�Gھ����� 1a~���b1X4���,��gq���9*	Gn��������g�v(�5��m+��6I���[��R����B��8��)EW�9
�2w��>�۰��!r�%�Aj���{�(��#23�ځs3����v��(�m-��3{��}C��I��
I�Oz�0�wg��ia��@����Jx�M�'F8g!>�4��]�$��m:�%L�W$��x�?��C_�dȂ�	j��x����"�$i
�MB�}y�/�^A$�F�����.�M�K���	|O��o��]�MU��-/��>���)̅�.�(��?6���nBm<�vP��%j�8̋��l�@`9�ǖX	��iV�􀧬 $n[�D����*��)}<\lu%���� �\*��-�H#K漝r�M-���:��+�u>��w��	���8����;�5-qh�]�$+z?Ȥ��#�&�����D��njk��~˸���Ь�u�O�o�KXPr��(݌2�.��q�[�i1.
M�V +E`���Xq$�2�!��d� TO�K��7��?&��^4B|�Lty7sے���ꄅP����-'\�;�|�w�����If���	x�.����WOR�o�E|7QG��Y7����>���Rl�dKv���X
�K�qu8��#ɽ���=~5j��zHZ>������yP��R�`����i�J�gS0s� �Z`kB���:��k�N0|��p��P�᠏� +5p$E�۟����߽c�	b*��۱�پ���W]�ZW+C��E:�G�2�ޟ75t��E
P**S���#f'�x����O��?�Ĩ��ӖrC���l�Qޫq��(t�xfUPO�v�W<r�$1¶P�k�J�YN7�Tl��C,�0 ��Ó��Ģ&��OP0}g�7�������g��?���PƁf�du[i���T]�eW�V��F�I�P�<ض�_���V�e�㚴���:PI�����sQ/m�On�*+[�»h�5�Gecu/�k��%��x�AO��s0f2w���>,<7ض ��A�?z�sp��ɫ����z/w�RtQ�e�<�BT6i<u�7p��q.+^�r����������&��P,�Q��i�R�'� ��j���ﯣ�Dnq�v�<k�ע7���2mT[�z���P��T�ɴ�2z�YCV��\����Vzt�D=�*�u��GM܃CV�1?�!�|����6g4��|�^�j#�9	�Ӷ�Gy�v��M�x;�@h9" ��([�gǞ6����u��l f��#��]��5H�p�т�t�C̃)���s��IĞ���GY�H���1��o5G��v����3bҌ�(���r���=�I �-��`�0��tV�cf<p�Tl?l����B�\c�-r�՚�0O/k��� ��V��,��%���%� ��;��_�AK\ui$]F�WVuT��X��Y���:Q�u��^�:˷�{�WP��,�#�Aؤ�u��TaΏ�$��8�/60	�&f�%��i�w�T�y��MNk���A��t��~�YR�uuK'�">���F��,kD��c�;�ך��@�l*s3
M3p_�47�e�2h	{��i�#d���h Ӣ�z\�߷��&)
$m��J&�g��͟q�i�D]��_w[>�|���mh����Аp7�'����� !����x�3[���2���yfx��?��b��}$mҗ�˜Դ�f�^MW��^?�����,���8���!�d�bH� ����}�m��u��"t:���"Ҙl1ƼQ&�^o�\%b�di7!�d꺌��	�����6�O��i �A1��Z�ҷ��
�ü��p���5C�/��ν���1� �v0��l��ء�Y~[�eLI*�&�U����)Va�9����l}@��|"{�A�H��5<]p�B�3�g2*�[�M�@���*������i�)�ڀ�AB>���*��O ~_��5w�Ps��Kvn���WiI���%��h
<��'������)W��g�+kT�
�y�ԧ�Wa�uq�Vp�օ޾=b�4�F��,h���c���h?�K�r8<�� d]�tJ��q�M��W����[���:w9^0#\8֦T�x��ݦs@, U�<�bf�ՕϮق�kL��>AW,N�n-6ކ��fn���,�����"P��Z�l��*&���O�����C�����ˡT�u�	õ�(:��a:���׻<4ل*0c���޼�O�Ξ��%ټ��|&�#/�5�t�6�:�� N��(���p���6t�""ڟܯ�9g2��˱�W�'Z�jjw����"&��b_K�P#���wv�c�]|�=
'�N�Z�4I6����vo�#h�c��q��7��"�_7ڧ�4I���V�=>^*,��]��d��q���t�?`R)<�u�3���	]ވ�>V�%�դ$Z;O��@ͯ�Dpqg%�<��xL�r�wk@�0bߩ�	M���M�SeZ���W)O�AEHvB�<|J�����'�i�ӯ �X^��W]L�"�w�lc;߄��5��X�
�޶�w��B�^��������Gp.)-X""���%���ڋ%���jPFj|G0�8B	7z$�UK�7���L��CR()@���?,
4���N#��J��0�mX�_���';8��NH?l��Ûҭ�����E%��3Q�l�N�0��ۼY�]�P�݊�@|Ҁu��:p�,����K�?7N-�|A5���"��6�(x��N2S&��K&��;|�\#֣�4�D��kAt�ݮqH����U�r�b(�3�y�yQ�j*7R���Pg2�~�Π�"�������".h0�Shl���$�H�,��W$'c(c�6�?�#�3'�f�(@��;�1�CF4ZE�F��MSOs����2\y��AP�;�8��37:��- o�#Q/p�-F�ǜ�Wjr��Bw؉)U��UI�e\^�Rps�d�� A�a&��fG%߶F��W�8IO"-P�0��=�P�󸧽���ӗ�	Tlġ"z]�m�m\v&�(���+����1F���Ja��̆g�gP(�8j݋@��}� u��S����1W���2
:o����`�15̱˯A7; �Ar���ʠ���9acS��O�H�j������d�^�t�X�W6�۽Q3JB���Q�;wl�_���ޏ Q�J*���6��K�MM~�����5�W2
�>e��d�>��I���Yھ6�s��[p[><��B �CL9��y�Ѣ�1D�Ү3����D�[4k.�+�d?T��}%;�1���OX�_Y�3ܯ��U�Ulϑ�C�ӹ��/*#���{�E��������yv��M_ǕG�[���%P�����ٴ�����5�	(5�k"��TX#u�8��N�T����g�� Bt���6��ӵ��*Ӣ�e	X��S��}�
�2��ͰR���WM��E�m��Vt�v�x���p-��s4���8=�b{<1�J�^����Bc.�;wU
/iiA
ş�C�-+������V9ŔX��3̕)�y֖&����1|��K�w|i��~�����)�����I�B����[c	�:X�z ��b����N�7zc]�G�>��fQ��XDP$u��5���)����`�f���3�,2�Ê����x��j�'���%�;}eJ'�e��)�;��b`e�G��*�wMjn'q��QE�S�RoJ��P�8��_��L�[2H�Ł讞��|�����c㘎�����j�K��L�!Ȋ��%G!�����{y�2�Ҷ/ҕn!�Rz	�~V�߳�#�-�Exv�r;�4���9ö�Qja)5��V��ԹȢ�	�8 _8����2��s��{[�0��!u^���f�f2�%��n"���a�25�nD��	P'/x!2v��d��l�Iގ�g��Մ���UT�mj��T��!j v��y���j�T�����,�?D"�fj����Ɛ�hi�͵�Ɓ�yU�,[N$#ã
��6��88"j��_����M6��Ӑ�FIu��[M+�m�C9�8 ��Kr,�դe�8� 
�������eX�13u4ՃAf�T�i]O~V��_��H�D6j�j(j��n.��YM?Fky#|L�����[����Ј#P(�Y�e�V�4]�i^��^+�}0��R[P�ϡ�̗WP#>,n�	� �L}!�(���� d��H�
���x����A<����Bl�����I�P���dw�4� ��T�Ay�� �����^9CۢN�q(9��k�����t�ᆴ��e��W����8o�@���~L�l��:�f�XP�<9��{ D�I�����%��k��%�F 2���yI��][�i��/W郜�~����d�@��Ո3}�:�qgzMG��N[w���8N��e���S��.5Z�a(Y"�_��?3QNV���dg���X.ر>���ȑO	G��f'�=��>A��A2@�k74u�Ir0e�N����������d��^��tsH��*?��A�s��C-���YӃJ!ڌ��;򣺓H��c������Ei�����@s��t;�{�7yv���O�D���NH�S;�����Rj�*}4����ӣ�yH��U��>w�����dp��nh��]�������|�@y�WB�����z�����<�Mk�uT��܂��m����~}Et/V�@+Cc̉F�X��O=�"y*�qV-Q�� *�09��ש�Y�?	�X��O�iӶ/-ؾ;|��!�!�7��Wؿb^s�w���C&�z2[�������`���+�,�4h�=�t�A��C���;��qd�C�����81�a"�
j}|@[y~g��iq��yr��'��j@o���e�F92�L�;q�I�������=�۬�/���+��������)1=^����fI4߉E��X5l�׏��[k��� j`������>�d/xC�e��O��ibIQ��hX��"-�WK�V���^82v����ٵ+�gSx���`���HrH��
�X�"�.�g�6���.c-�F��/[mK��mws~�W�S�v�g��2^��5�?[�L:��XW���h4��K]<��I�H���{�|���nm8S�����z"ka�Y���q|���$��Z�ձV:`���MƵgPhB�[��ZLW����,�hة�@P�R7E�V履�����a8�c��^��sR�.TOV�P�Z+*H�R����������7	W��'�o}�o��Y���~͈�{��]b&�L����d�J�ey�,#Q�)U��J�Q�� Wtˡ�eX��BDO��Y-�An��� |Ӏ��q���'�Jrߔ?�0'���޴#l&2���XR�����Y���M�.��8W__:��3���<Zр r��4a�}�M,���09��F�B�=��"B���%������S�j��-���/��%���R�7[�|���1��NI�ϚE|14�[�������:�,K�"�ش��ܫ��1�Y�#�x���d�+ɶy$���$~��U��X��� ���dgzw��w��e���b������'��j-��k�=x���:�ׄ�g��<J�x (ɼ%�s|��e���ר~C��±�'�>�����/en��)s?�~9�`���GUR&ƃ3�?���Iʸ`M�rYq���h�2����xz[�J�1�Lru�t �h�J�����QK���"H�������`b�=�LC���� j��qw;|�t�PKY�!�/��{)'� y.����:�4yZ�`)��U�������$���$�Lb@�9����Ӡ�rW����#��O�ԯ�]:B�͞�`vt���0�?2^�gŦ[��@s��"���G�?(Vk4�~��PXϚ��vW�MS��a�����+.��ZhoE6�>+��R��âPF)��,���)����Ӵxui�C1�\eǺ�|�亵� �y�7��6�������\=�47��HSM|5�&G4z�9��H���$�_��r*A�*MC�S�B{�ϵ�c�O��V�1�l2�zH�F^��uM^��ǫ�P�-�_��P�^�i"ҞY=�����9��֛rF(�s����q�F��������R��N|�r�5��t:�ͦ��8H9�A�U����]����5�Oq_�#=V�����j��2�i��xm�$\&�R�=�y���bTa� �Fe�P�����\��ʎF�yL;-�D1u�CҶ|���iU�	Cg��b�O��d����`ɚ�tq��c�'�
�88�'f�o���>�(c�*;M60���sLb���]�ؼ��$�=HTy�A�b싩�vж��j@w%/ح@���6���@���D��T���C�#b�<p�O>.�����s�T,���� ��u�n4��g���)^N��a}��-ma��}����,>���U*?��	lC���0�F++�ZB��NG�pĬ�@�� Qj���
�x�X��w��o�Y;���΍������1��\h�/\o���{�~�-9��!G$Vp/���^�Ld�9H�C��P�<x�7�ÜT�lM4`�h�[�#h���`��=7+<b�OU���7�$���0�<r@f����T-��s����~p��e$|k��yT�����:�80N�" *ZG
�p������s�Ǿ��Ї�rW�&!�1#@5��f��|�^�]!��^�.�'vRh��'�8*�+@�g�M3����)t/�>��۰�;�)ƮЏOd=�	�Y��kp>6ek���ٹ�f��Q�f���� ���<��~��	��5�����x�IF�1�w~R��O�+�H�s��u�eB�c�Slf�5淧�r>46�w*Ws��P���-�{ntJ*���y<���W���$[��W�zCG)�1DkH��U��3��*=VD�	�|D��YARZ.+˸|ޭ\��mF3永�w��R��A6�Ā�	:8'n�����+Gv����Q�#^��J����+�i�X�@�E7P���_�����-t����(��ې8WhʀZ��~���5��o�OȄ��s�f�p ���KQ^�u�ZR4{(�l�%�TV	�Ê�i&e��#0��N%�K��4�XlkzC�u¥�D���~�Ӑ(].*%B�[�D��89C���d �.�e�{�����U�f�Z3�\��3�X�8ƾC�£���
&$))(���!^*ތ�[���@�2�RM�bp�,���]y e���$�ܢ��Q�\� �-Kp��[���[���G�UP��� ����\NDdC���:ƗPq��0���X�&:���-����'�y:T@�o��m�}A����\����%��RQl��w�;O'gݵ�J1*�fv��]���l)���p�U�X�2!)���SCDfr�5ߧ�	Αܻ'�G��eK��b�z�Ѥ �G�>�J̈ p�;�[��42*�G
}�G6���Sܟwυ{&�J�p�1Ъ�!W�:��7c)W@���[[�%T��ܬ�~ʯ��E�h�)���r:�&�62�H��l� Oy���C����Mg�2q����o�;�z���]H��g�-)���#��@x��Y��ںm���٭@�_{KYgx���]�
Q�o�+A���KQ3��A>t=� Bc��\n�������~��=*&�Ebd��5^�_׉�E!/�o@��� `��Cc[q�&K�%��5b&U0��bU��Ƽ(��^V{��������^�ڻ���$F�b�9z*J%�B��ߗcs&;l�~S+s���<�\x0��M�n���_��V�b;��nđ�(0��<��,�t�9��3}UcU�4����Rm7u��o��C�Pc��o�e�R��v�]�ӿN� s�����xb��i �����*���}�ٱ�Y�0Z.e����-=�h��]Ib�=�U��$!�p[!��o>[<�l��t,���r��~�C��8��Ź�p'W&��]�:=�s�5�V�.�#2��r���f�.��Yg�:��!��C\V!����������������o� )\��w� O:�X zw aǿ��	|!"+R�95uC{g�i,����d���;������f�i���SUg �s ��$��^baŖ>��_���o�m{(8p0M�u�K�-�^��\̠�Q53)�v��N�[���?����^~�}wA�^�t�M���v���6v�5�QR�(��,����Ÿ���D(.���-�%�K�x��Җ�0�2k��y�w��E��nn�2���3���m6X�rQ>_�S���	Y�m�s�Y����X����q�>	������X���hs=�v�<4�;������[�MSV�v(�K����<Ay��q{Rs�k8�#%	Z%p�& �3f��U�<��v�l�}���X^1�1�J�%�_Q�r���_���7�%I�����&�>@h�\�#{;wC���#t�&��{7�$^4��� M>TvD-e�؆W�?��|���(%(�,]����uS��߿_O;�d��l[����[�{Je�Ϲ�R�d-�h���v,ǐj�ۆn��BQU`� �1E�2�"*��q��D�1�5C%�И����2�D���˴���_N�,�؂L/Z�ӱ�5�W+(�L��lF+#��5_�NS��=�m�@��M^57^_rc���$D|G�Tb5�K���+*�o���=���Nl���^
�7_��?v�W�_�a��q�2�Kf�{�Nށő�M}�8�$�ߦJR��ޖέU;�Ņ��P%Cj�1-]s6��v`�PF��O� uV7�ƱR�K/�5�;�͂�p�'t�c6���N�%v�;ҚZ��*�Fyd3e�A�b��tJN7�N\���y̓����d�e�B�E��+M�2�ǅ�E�g'�Q��n�}v*a�s��,P/FqD����J����MP���~�|e	Vb�WYk`sX��,�-�aN/�&�;IikD�h����$�jx��=����E�6��^�A¢.Y�쎽_�&��ֶ1��36e$�$J�r6W�j�$�ױ��z�E���d�?+n,5���7i�ȒN��5p��`iY~j�C�<*����~&hB����n{_U�V��:�d�WQ&�7��p���qW��B{E�'�m�%����O�M��F�.��	S	��ij`�a$|8�$�|>p�X�Gm��;��ن���	u�2!\YX�R3���#�8���J���(�=����gL�`�me
����	�Q��2y%�I[��;$��:�a�phg\j���{���%S�O�g��������56�� ^tͻ��g'�X�;	}�x�҉߸l�@ze��@�E���2�@���_�n�W���o�8�Q�_����u,��L����q�uGx�br%5�����������=/t��.�-O��p�����]�=�����9���t�Y<�a,i\Q���1�������9�cl����Π���w�ɫ�H�+@�#�Y��FPy�[�Gk�gZ�����������j��T�ς�P��@^���8�m�5�5R�&2_$�Ր*���A�YB�! �n��$��>�5!�N�a�s��ޛp�,�P��'����H�J`���*^�q/Dd�x:F7��ӢQ4N4`%�&������Ľ߀���^6�׉N���9_?78m���ݪ�P��M >�fh�Xȴ^&Ol,�%2F�1���i2�h�T�6��5Q�u)~�ĕ�9
<q�k@����e�2���)�ޯ8�l����_�����}�^T7w����5�os�^�oM���������	�v�D�K�4/�����!g�DD�l�>��ѵ�~96ԲuuHMڴyW�l�L� ,�	���Ϋ�c�G��f��}��g��8�4�$���|�^.�>_a��?���4������-O`;��<��$��J�$��s)<0s��zS����Z�m�l�,�3�.R�r=2ڰ�T������dO<5�D#�c�9`P��tS����%��PC+Z���KR��n]�S8��%�|���>6��>��������٧!�s����)?nSs_��S�{x��AƸN�z���o�'��V��q#Ǭ5/�P�{�B�� =3^�*�u{t����a����p���L"YYqG��k�{�(M2
fX&aT<N����/�O��X�>k�ǻ�}�f����*�Za��"�/*�S2�<2�B�%yʍZ�5syp��0�<�6t��M;\��nD��=�IYf��tّ.\��7�5fD-��?b�nD�1Z�Zҟ�H���{/�|jPG6���~�5�n9% ��̱��]4�����)����lf�L\�KEW��G�D���h���!�� X�3Rk�vȩՀG\>iNx4R�N��jK&x��
/~�,������)�0���5���;�孑Rk�x����(�6@cQ��tX�
M3;q��+8=QǍ^( 9�yt�55.�1]"tG;X)^�8�V4OZL ���p]U�;T�&|�/�g�V*�o���~���#��"�M/s�m|�f�����r@�D1�eD0x�� 5�p�][�mHNz`��U�We��9%�Lp����Jk��n�,�1�Z4YYC�T���hQ��j���w,����_�=/��,1qG�	d�����e�k~�f�I����6rO���bw(OR��T�q�b��Q�l�<#�qI4�}���\�����3ݪ^�2���֑xfB"u�$���#��4���Jmfv�7F;�&�a�Fb��}�fSG/�ݠSX�+��.f�H6�2yN�S���ΐ<�n�1�v���P��<�Q�`�Zi��E�rRP�甓a<��r��O�Ф,@�}� ��q���$�xS�5$�\xhT]TW���)m���2��0l�6:gI�IG���vtw�n���@9&Bpp,��f���OP1|�LW�V���Bf�����������U�d��2����Tr���[]~�gp�X �o0у��\(�C�,?�
D�/� _+�9����XQ��k�A'jyi���鲎�s�A�P� �j�e��
�IKA��L(#��%�̏�l�{D���X���˼�(�4\�� �p�}��\�e�~(��,��$�Z�&�`�.(H�t�%@���!�~j����wq!�RZG����[��i`�U�� ��s'A���&x��g�$�5[J[DŅq�A����Z���Q��}��{R
�`�NUI+���C���u*���N~�f0TJ�i�J�e2�K��_9,kh��Q׷G�ٲp�D+B�aI�����o��I���ihp�R��r�h�K�ٍCqV�=�x��wr��YZ�{`�+��4��R_��逌��RF*�<�F
�c�e�Ͳ$����ⵡ}�(����.�y��]j��o���MaQ�B�ł�c;Kf���k�tR��mD��+�� )d��yJ 2����w���ĩ�Ἳ�n��c��R	uf���g��XV'��I~	��߶���z=��V�|E���9��D�@0��J�'�c8A�⯈ƈ�U� ԻQ5ܫV�uɫ_�έl�үx)`qoI�.�}W��4����y%{�
j����F�t���
��*e")c{+���?M].�G{_Z�e��J�h�����	�y���v(��r��୭�Z������s�><��:�.1e��~`��(9.Y�^��J�?�D�Z>݃�\�]��c{�#�U��bq��2��m-P����2�ǲm��~���TW��L/�ы�ӗd�Rf�Ai�Fֻ�kڪ1�?�z�ax�#�2.=z��ד��'8�� ���Y1�����e\\��2jN�]�6G"�7��Z�����rN����k c�N4��UHbyf�+u���R)�jIZ�	��?��X�g�"]��fm^J���3Iޛ�g �}������"�r!V'>u$/R9�!&����SCH�q�����$������'xi?$>�O�K�"����!dMk<�Yb�ՕE�������=���n��)�\�¹��&������m��kC�zS�7�ɲ�:�I�"pc�\,~��J���c�l�k����m��k�˰�}O�����:Zg9w��f]�hL�SI0"v�b�?��[vmA$����e��m˶���·9������s����!�mϛ��4`�z���>"&�#�\��y�E���`�~�@���������,��h���_�����g���{�o'gN(�����4�>@)g�e�; Hh�k�.z�rK����yͫ��m���C�b5������nX�G��5 ����{S87�8^'6�[���G���#v�_��m�Pp�2˾��@�ȿs\xI�m�q.�n��%;9̓�������{zU]9C����8��|)�B�_}���bw��e#��x-]9�D��2}���5���& S���3m�<��װ��E�U���C�H�%k|�7pm'�H�H?�J���@�k@
a�I���eC|Yz����<�O�x5(Cf��h_�f���_��B�9D��2���)��ƙ�b4h �cO�=���˲#*mP���_���F3�� h����c��ȸm����\�D4����9d\�:�8د��>����f��g���`ފȁ��4ՈR�4$h��wY����1˓��L�#�B�#o��IB���o*}�y�}����
�V4T�Q���N�`$�K{�_�*�e�\��1}&��%��煘�=gN퐭Hi����π.R�]��(	C$�$h߄3f��8���icA�Ҹ�r�"�3��-b��ϸ;�rڪv��!5�l��@7��/�:�YNg�)X���t�3�z�(g����	�N�9y���/v<��ȡ �r'�Cy�c�� ���@C1��TY�3^�Μ�t�APG��oVJW^2��A�w��ѡl3j�"�T�$j�p�܁e���U(>C͸�Ց
�u��7x[*���PA*]���Ӌ���}�+w��x���|���: TJ�2u�8l�%$�+H%
�;i����ͽ��IT�(�����w[�!./[u�iO�"Z(�-d����ߧI�!��|@N�N���;��U�X���v(�-�#��
�f��B���zW�'2ؓ\b��92���*�t~�牾�Ur���qb�ơ���@3P���҃tn���q�
��ia�.R�u=�$��scp*v��p��%4n�'�RH�egb��vY7��rhu�z�e?���W9ܤ�l�U�az����ƪ�Ǆ���y��<�Zl��+͍8��=2�?;|Zز�H�4� ���52�>a�t�d���k����@��ֻ���*��6�.o����bF�w��[F&9�j�?�(T��u�\%�����ߣtm^�䓒��@*l9JMG����_&A�Ɋ�:L`?�O����8^��I�r<fG�]�VfwS���saG/����Ot�{���8Y*S{��Ď~� Ǻ��"�.��48��m��i�ҬT��ˊ�^d���юVtq��D��޼��8�,ϖ'����vG�Y]���n�km�~Ъ6�;P����Ǥ��4�yfHۢ���C[1Yw������7h:x�ae�b���?�`Z�^���:��P�LD�E�����lއ�S��,p��{����E�풎�i9���AX�t#�!L�������o�j��P&[��@K޾��z����L�sP��4��3��������_�Y��<��Q'����FxQU���=0`MD��jdiP-��ֹZ�qs �uȴ�X����^�V���F���� ���ޢD�Qӟh#�j�8����ɀ�@���!WL��
T�T���!�%�5����ț����j��G۟���� ����pk���!��5�w��^��V��FƢ�yv�z<��WΣ��WE�D��Gu���H"�5��ch�2���v��k�kϡ�Kߺ�s|�"��ޓ	C�h�k��A�I�s\����Af�O��2���Rߎ�;x�!U1,h��,sA^Sg��d�����8F��+��I��Y�Ww��Li��a8a�C={���i��:{3XV�����C������r���#Ě�3vj����1�����Tx%_�{F=,���mK�0D�*���8 C߆7�C#(}ǁ����&	�N����r�}�U"�8����4�I&,��5���8���QB���iop4�*���q�
�Ļ'�(��;R�� ASC�y���� ���.��b^��+o�F:[CV��x��G�,�&��L�9��M6r���x���虡B��UD���V�g��s��o cg�x"��x�0{�>sQÀL���H�^�OQ�5H���n��Y���r�b6
�H�*h���ݜ4�"�&�je�V+��$�/ߌ$(�΍�(Ð�Ꝡz��﷔ۤ�Æ������`��}e�:)�Q�TEgx�� ="�G{�c�����C0;�K.|s�}��rɳb�zE�w4Z�����2yx�����U Hّi��.�F>[%��Ҏ}=C����e*�tƅK�:��[''gG�S�����ҥ7i��_V��������}��������WP�;:���P��gů-LG*�7�<��X�/_,yf?3�.Nlqf�LuQ-�lf�M��c<P�ަ�"���h�=�|QM�<���`a]L+�WM':=DҬ��|�!�T$�I��\���;�iv*�Ʋ��_�l�c`� K���m|�<s��-X�;_�˞t ��"g�+��m����V���C���VxVk�z�Җ����kL���?6�G\`�W��RN9C�-n��k �]�V��`�E^�M�Y4sY5\�p��H%%!� LN7$ũo���R�PIKe�e�8�Ý����W�hK�&��Ǭn���q�k�+	�$�E��	�Aɲ�c�f��i�r�>�7����Ҳ(���b�Rm�0�'�+4�Ddb�ڵ:�]���C��H���&����x�=���������[Fx'0��d��h]����,ƶ����نR:��_����A��lgy����ɶ`&�N�rw��:M}�(+�����\:�R�ߢ�Cz�i\�`��}�S��3qdL���oq��/�+J2��A�-�^��^x�2K6}<�f�P��I&8,���s$i����%�������5�L8��jC]��I��9��d,���E�aZ�u�(���.L��+n�>I���@p�ri8^\4��i:��e�x[	��^�U�U���k��%�ܧS�PZ�l;ԯ��,��}��oK�$nei���Ejcc6�)G����E����l^�01n$���~u��5¸Xq�����'wקc�����#F~z�u�|�UT�vʉ?F�<��zK��P`�
�7��$_���^�W;?���0B[�!v�yJ�#��h*0��u��@��U�y7���#�_��;/�L���}NJ��zc6�H�d�UW�B��u��ӻ��Ɓl��b�w刷��X�z�v���C6<��?t�ky�]�XhâR��YGE���t:�jT��5���do�
Ԛ����u&�VW��,��?�6�U��+��~R��%�=�`7sc	��c�PN�:�=-q��m����s�	N� �n�I���|5�:�/L-K��:�ŕ=Q��!yY���V���e���̉ρP��+$$��,\X���`h{�p�xe��#F6�)��"zL��� �X������rQ^4����I��`-{�Ѓh��� >�s�P8��:��p<Ѣ]���@�rM�07�R�G�Y�*���e�3�ū+(Y�q�]�l�����y�F�M�ؼ��{�:Ew� Z�I�����[R~�_���k���zo��&� @G���%���"�7�AJ���c�����6{���D��� �+���2j�5�w�N��Z�/q���N��}DF�<��7V4�ѧFw���_�)����M�FZ�s$(8�e�\ �ﯩt��h��R�0�GJsL��1�8��'�}�M�x���ES��*�LOr�����`D�J��ʁ���=�����>B�r�ԬWD���c���[Rc�Uy��M.(�T3[����-5��pȁ^v���X��]w>�����e
�u�, ����-n����]��M�`�-��~�%+u�)��(�ߤ���D5�A�fs�&)�
'��<�)�S^��ݠ*+�`�Ъ�Ec��M܁G#��*�I'N��M�lm��S�n∨ܹo�#��I�.�4����g}1 ��ŉ'�(�mt�+��QyQ�q�Ì��g����[�b���/@�'f�^���[ 9����RW�5*Yq<���F��8]�H�j�I�郸��I�XzTK�X`R���d��	�(�5 g�M�OC�������"��9z��4	���T����UBeS��?p7F���k\}�D�I�V2/¦�ˮX��m?�kO �aѕDbǷ]�F��e�m(N*���o��,r�y�ڳ��=��? 9��x�����<@�$��:`H����1_�q��!�z̈�!��]��M��DKp�Mj����EV\MBI��E�͗�4��[ IU{��"��;}��=fN�{P�>�R^U �!oS�:+��m��q�j�A�i(���p�#����:2��)v.�R�r!�g���`<L#�3��R���~����7�)M �9C�I#l�Kr��2]ט��#�e��`Ѫ~d+�1Ʊ�&�Z��K���>�Ъ,��R�@�!�1�-#�v{D�|�+�HI,�Rv'm=E���Ċ�Cz d��m>��8Ū�)�lZp�O������C	$Ĳ���HY���왧��I�sSO��V4�J���sP��QSO̱�c���fl��}��K�Z��ep5�iɳ�Kz,�pþ��m�_$?�t�B2��j�"�
�ރ�8��9� Jx;u�םn��Q�c(���������N��FocN�pY�$���!%7r���$W$[.��$���_ ���V�\Ye�-�����RD�(�}�$�px��C2�#�cɄ�ʖ
�2)���)�CO����/��.�A��H�����ȗv���Y-�s��N�: ��Ʌٗ29���3SiwP�8��:e_т�7L�Di��}��BC�V��y�Nސ+�:�p�����H��G`�kK<�!KF��b��F�E��j��D?.��+iAu���+ٝ��M}���UeӾ�t�W�wF��89��� �C�P�0"��f��Fi/@���@fO7axEW	o-졍��~��#�?P2�i� ���k�A4\@Ԭ"nd����%���8iiH@�{ŗ��ޝ����jUI��-����Z��>�FGwe��YZ9�;��.pb0�m�-�O�u����:봻��<h���� /�娠XO���w�-�F;ya�.�xg�3����C�"o�Kڡ�6�9.�h�ɓҹH���M�dr�-����ZO8=~/���9s����k�I}�V�Mρ�l<j,�����7��f�,�-[V�@a�1�(ʪ�C
8Va���@چ��}�d�x@���q
	r���%�16�z#�>���<� !^(^Bx��U��������]`�C��B#�a��b}��1����K��#��͟Y^9Fi�������3Y)Z0Hۜ���Bl[f,)��`�6u*$���d|wN^i�@C��:�����sd�bHX�G�<�.��2_���)��:���-�Z�u�  !�2��K���a�l�֣� �:�{����#{�|����j�Fmsg6M�J�Nt��A�<���*}g��nh-y��h�U1���N��;������\���\c�H�Y$5��EUy�P8�g��t�n��X�	m�9�2�k"�<�6nظ���Ey���'ڂޞ4�P� Xb��Ru�V<ux��V��F5AA�WY�V��xx�eB�a�2N:<g�q���:����,��g�_�8VP8�������恀/��FW�n�@	���s�+JR��S���9���NJ��9�3a6x���P��{���J3�ce�����|��I�h����kNN-�Ëen�~�+��
.~�6GK�3�r���5�#
�9��m��m��D��A�L�-�=���X���E��P	E_g>7�!��[O��N��.�y9�_?�\<��ĝ@ĩI�I��L���O��{�bE��HKqm��l��6���}�#:�t����GӇV���B�x����U<k�x�%�t��c�sp6G���t��io2�-��O��2a &��}Sx����U�45��:cۧ�"� 6Y���J73rj�} ٟ���A�t��� �w��
	'6K�ɨ@~�������`��p@���"�uT�8�Vߎ���]�?�X����c{�������Î#p���le�`3�������l@y���&z=R��y����Bgˎ{��ͺI6��Y�Ds_����*K.,w�E�U�9�aF��Ly�oc��\����]~��/w4�[e4"eA��n)�ۏ�8��|�k3;�����en3��Ѿh�<ӇRb�B��'��i��n����g���:�Cء���c+,�1������i���`��u��	�A2�����}�f�֮�����EM�:)�Nq�֮o=���
��%�l*�pbVH	�.����kH�������"zJtr�εQ��]��(jC��S�#�+�x���\KƦ�,�Y��7�0KDOM��=b	���\��$!���N�]�.���vNօH��T��x��.�	O}�I�%�De�+��r�j����r{��LS\-��2�r���?�rUE�ء��75��WKo��wy��jα0�T݀y�����?G��X[k�ډ~
~�;(�D�6��2�Q+���K?��#�b�����/hD �.����D�lz��&��J%%�c	����E��&�p���oQf6���R�dv|�j��Z�2
����+!�J1�O�Y����N�+[�}膡�CYkqR�R����_� ��u���	����s�F�7�T*K�0JV'E$>�.8\��u��;�S��@�ϭ����`�n�_�l��j�Z�8З_d�$쮲�������>��-w��T�M��.-[lF�����U�Ɋ)ko��8�h!��
D��޽16�;�6Eͼ�U_���f% �y�y:�=p���(Co������W�Ⴉ��;8�e(l��*�$�x$x�ӆ���p��<p����-[@h��0��i%u�~&9 \�=�
��:
H�w{����1!�v��7����&`S�t1���mp��hԅ�n��ύm�����fE����Er,<
�`s`	�,���\�~hp�?�A��?Ah ��)W��Jé�( @��U;%J���T�W�N�"�hiv�.K,y�~��%�{�A�?{���;<�����wQ���pT�<�֧�{5K���YtTڡ���D�~�9	�7k�锌�Z�}�d��أ4����p�y8lZ�IF�O���8a.E����Q����v�<jCɄ�A�~5C�ݍ_���;�/�����r W�3g
L��j%LA���}��C�2[�ާ*�W�r!ZE	��.���Q��JA;Z�h�jvh;.| 6\��_ƍ���`�����O"Y�K���E�sJ��u��9�D���H��_oR�)�/,���+rF�F��sNXo��я�i��>�w�p��-��A�z|�!�0�٦A$��w)�6�7���"�9h>�l4��\�b��	���r�"�z�/.�!�z���	��_�UB/���l����Qm��Iy12f,��a�c��Ynb����I-�u^f�V�g���^�2_�q���̥ccm��t�L�$ɖ�ɓ���{H��{�@�<�����f�L��n�pB��k�Ϡ��
$��q�S_��o�}���TY�I|$m���^`1O�W�S�V���W���n��-B��MG5���L�Tg�:D�a�^��
2UxگAi.%R�̢T6�&���_��O�GZ��|GZ,fŎ�z=���K%�JV���k����a�9 ��X�_\�f0�_�Զ�i͟��,d��ܠ�w����.��{h�y	��{/��5��fLf���;)�Ӯ@u�e�ԷP씃�'��M��vi����� �7�ˢ]�}߼�C԰jE�/U�3�R%I�՞"ջ�(^��q��� ���r�^4�RЍ£�4ž��Mɩ�3��3�vAc���扻��#ꫛZ�������mr��e,t"]�R�e�8㋙OBȊG<����0�_��N<��e��lPe6��Y�!��"C�e^ ��͌f�����*Js[B��s���c�T�h��[�tD����_Y��E?&ln����x�!��W�*$)����$���w�d3�����p����zHcV�	�ǣ����U �[}
��p^��փ��'P�u��'�S�]�E=�	��G|⍜��ׇM�_I�QȘ��g��q�R��tW�O��`\��2{t�[O7\XqE2�72�ˋ��)�\w��-/��5�ƴz"�(�6?���D-6=�H�ibW�_���r�����N�����@dr�DI���	�F�|�^"$eЎm�������H�)T+Ǟ_��7��L?��p"�_�<NlD	��=h���I���!P�]X>��W���Ⱦ�w��-P�
����pOY��,d)q-�Z�`]QE6�c�HևYS�֣�IY2R]��nM�B@�`5,3ݛ:�\@��w;��5�vX�a���"���p/_���ǻ(L84#�&Q���c�b����Єm�_X��r���KQ<�2G�]�]������B�i�Pv�_pT3(E�D��P�y�=���̞�i�/]_��v|ye��V�җR~L��s��0�~20��������QoP)B�K�ͻ�F3�C�4��6V�sY"ɵŝ��s`��WY�U�
^p�畊<U��9#T�i=���_ߧ�(���l�~�#�Bhx-�c�%�e��Z�������eLl��V�5������4���ݖ�C������@q��W(�'`)�ڛL�6#���u�M�H�T^�/�b�K�Ħ�F�|���a؀��X��x�ԍ����<1�|z�k!Wi��65��-kg�o��A�@V�"�u�#v�i
�~@n>�pԴ���G�"�$�Ād9��}U��o�|����m��èf���-��B���bo��@����4��� I�% �]/�%�ێ<�M����j���	�+1dt��7r����<�tܯJ��2��`b�6(��蛱�$hJ%h4�Yo mK�D�+�c��.�[Ad��xB�Ἐ�Ŝ�E�LY��f��6�#�e����_��|X��ilŻ�p�4
](��n�Kh��`�}�~��jv�*\~4I���և�\��8���Vf�b�fc��1%�t ��bp�fS��#z��k�Z��B��OQ�e���n~�m�	=G����-�G�X�������\ЯD��y;T|����t�n���蟸�`�`��m�3zVA�g��Q%�Sy~�a.9!-!�
)V#p�<�<��ƍ���L�2<�x�^|< ��sC�=��ڲ=��N�u������;�$ؖ��j����+��a����\�	��;�j;�f����q�S$rf7��l���v6t��rSa�����PL��s �!히x��;M��U�98��9au��2����q�����?%z���S���H�-�x<J��A�u�퍏�Z})�p�h��b�'��^}��{a��On�߱��L�۳q\�-Q���@ ]�T�S��\��ń'��O��i���w�$�<�����u��w ��롺P��uX�3��T���b��k�#�F3��d���F��1�WNpa�%���'
Ay�cC�b1̆Zx%�(l�����lD�}l�����8[�F�܃j��iKhõ�뉦�gV��ԇ��rF�u�_ף����?Gf���D�~ܕЂ4JUl�uON*��FD>�*<�D�i>�L�40=�a�w�o�@��
������o+�����ϼE��Q.n��٧
B����F�mJ��7�>y
�)�ks/��O��2�^'�h��y�c�U˙�>~��b��4�� �i(��+N� P��'c$u�F��f�2���4VG�ȴ�[K#���
ݪ�J�������X�5N:G�Cn�2;UW�N�FN;��aԠ�FWVJￒ��&[���~4;`-�/�x�&�e
P��=_.6ɑ�|2�9�z��^�R�N�������<��*f��O�쇢�y$�M���ʵ�;�ް,ch��0lx��X�!��ڛ���RN�1H7�v�"�bN��WX�8ʜxW �E���^���.Qu-·��E��x��� &)?�������¹���B�e���u��ׂxK���4���UI[�����٭_���@�7������`�PQ�do�x�G��֤Ӳc��w1K݂Ëɕ�;�b��M;����f���P'����1�:�{���D�}�Zc�b����گ�W�a�׃��j2��Q�ٲ���r�Х����d�t4�n ���������<�9��h�lT�ؙ��	�#	���*��� X�c%[���l!����8�l�H��?*~z�h�&�m"����b��a]�)�{�-@�I"ݮ=��m�����D�YT��D '���nh��!�u}���)��.����6
�Z"��FC�ټM�Y��f�� �؆`6�p`W봋�;Z��X�>�����F�ry�c����
�n��t�h{Я�qa��z�4���GK�*<.s�k��pm% �Z;]�z��Dvl]�wv*cpqQX�	�z�N�kγ�X�[�^�&�*�%-�S�>
"RfK��7CCt f��{�c>T��!'�_��e���^��R�ҡmK�D�������� �ҙ�z��X�X-ZQ>�/���B�E&o:��ͣ(B.�䅥ݯ�f�(�INQ�gOl��o��2���C�l �+G�"��p։sz�:�~�H��4�8��JG�V��>f-!ό㋘��v�2��o�]�A��� n%��6��KЫ�"�k$D?�G�n�W�
;��"\v(��l��s���NR����:�Z�>1���BG�dQee�%��=n��m �|�#	<pQ 5�N��sP6�@}�bg���)*�����7G]�i+����:�(hx4̈́��d,�u�2dn1-O���s�YDw\��z!���r�ա��Ģ%�GfQ����S:��Jw�N]k^��M��n*��:1 (.��C� K�@�U3	�`��u藫N8�3g ���.��2D�ݮR��������`(����o�?�^Ԋ��G�W����E�[�d`��`\]{��ڊq03�i�-wm�������|�	l	��/أ`J�)�[��ر�f�!��Ӱ7��M���ba	��=����0�%Cc5��
���і3DQ*��K��ѿ���IG=T��'{(ᦌCH#��Kx�6ڼ~��������=����{��=�f�F]ܽ �S#��������%����eiF_�[�K�G�����Hwx	��)Y��1}ٖ�ً�]�%���XЏ��@q�����[����DYܭ�Vp�'���>�O�CCM}���(kT�DSF��w��ۃ��*>����'�f�΢{�_���OzdR�&����f^��� �>`�u�U�*}o�p�J����0L}�a�2��o�%�ҥ�s�i�H�'R���-�,7"
u3��F,�m{#Ȍi%��퍪�dt۫V>E9!;C�N���:��:{y�re���w��nc�Z��	�\a�;� ��^۵UF�}d�	�_��"m��K����ԗtZ&��D~L �W c��Jȸ(�ƌ
�)���]��7x�R&m�, 1��;*�?e6L��yrX��/�)��,��ȜAT�Ԁ��z�Jײ��_KV����0��f�j��|#?���>BNkb T,��i�&NM�#��9��[SF��RK�n/;����&0��z�]v�J���tg���M�u^T���|Zu���2H�T���ō�.�!q
��4����� ���N��Udd;/�0�Ū�03��ȅ@��M��ɏY��H6�S�/��<_����u�h+���smE�M0!�䨬/6G��9aS>�3z��\�-()H������y3�G�����c8ț�X�J6JA�'��B�h��'JH�O��Mz�)\�G��6��+/Ї8*���	�����4��
��|k�H�fKx�O�;���݌ ��l���`~;��hj�n�Ci����F�d;1�R��39WR���Hg��al֗�/(@�q�Ὗ�����Ё����r�q��h'�� q�%�����<�P4Yҟ����nG�wӻt~5􉕤� ZYOCϢ�A���|��>��!+����O��/Cr#no�Ij��/��h����u�?��~4 ��O���S"����O/�&�t>3~����%IFX�1��i�>U%a�'�vH��c�r�߂3m9�\By�K8*x5*SC��v6�J��/�[�&olI�D������a~8F��A���+��VH�TtM����+-i\U�yd�h�u'��"��#�btM��z�.����P�J�ߜ�kf2�놕���������)}A��_�� =�E��gRRH�ϑ��-����?��M��R���<�(ΜUrn�"W��#nu(4�ͽ���1��ޯ@#�Tqu�)(���[ ��&v�����ށt�F����ճ��	��X@̰`2
D|VQ���~1���� ��~pPd���*���E��*����X�:�o�G��ݖ�+�,�+�k����J	憜 �;'Nj���X~��� �V3Kl�K��RP��w'=���'��VZ,�	�aAb�"�\O����A�5~�:-I�I��=-w��r�x����0D�D��=m(��p�,�~��Ю�3+��DD�n�q��=�v؈��a�P��=�����8{���>P�,������°�v����Qm|�>N���Ex]燭�3S�{� ���I�$|*�nP&�k㖔�M]S[�7�a}w��7#<����@U*�zC�������cdۛ;X��L�R��a4 �ɕ!Idl�|����EཎR�|��t������`�_*@�t����{��U%f��"qf&�g��ѓ/UI>*qP��8����:��5��}���KU�d�v��j�$@$��nW�Z-Y3S<��T���<�=h��Jk#_���2:��Ai\6�d<.��M ]���a�F�B}n���ɦ#����Ҩ��������$��V��Z^���z> K��\��:`���~@�a`˾�3��(ҕ{-fL_]!L��.�/Ql������'�U���H"����ͯ�is93-*�����Pؼ�hğ�s��y๼b��i�-����+t�N�zX((qt_���C�pf���o��+U~�[R�(����>\<)T_h/�':��.�}KL�(��*�"aD�4�#�*�L~����-�����1��x���9�	9�ȯ�Ye�h�6����������弊tKul�d(���q�����Hm9�<%����9��؉*��?��i���i(���	&4��0}�<~����2Qn���@6x��>�.<�/� �k�a3<�i�Rh9N�:�%q�����N��2�%o��w9����$G����7���(I��(ݔ_n��y��x�2p]:��8m�	"��:��N�r���!��*�#�DݨX�$AX;���^�gWC���x�f7�o����������dB ޚ(%�UK��1�b$�\��H�Tݪi�mK�%�;z%vS��h�dIJ�x�eH	�%�|��	��;M�xVsCl�£�x�kl�d��O��v���vI�M���%��JHëhqi���Ū��YG���3�pL�����L�aK��3�����e��DS-~���RP�~�+z��P�k�LY �Y��;��M&����{�jT���.��i�d@�V�@��Ԅ��[U���=����1�ʦ3.�!;���?�X�y�	���	�9�[����uU��ChP��q":D��{��/��<��*8	O���u�h��d��f�f6��)OUi `<�ښ�OM����Ð4�5�����u�����n��@o��Sr��C%��ӈ�i��r�>H>�Peh�Փ=���t�=r�D��߱(ݬ���~I�4(����Q���ٵ��s4ϭJ��$�45�}#�9I��Cp����E��/���O���
�^Q���z�=���3�HR�G��/p�G��H���R/6���B��C�j\��g�Ħ=0KӷB��]�je��(�huH�r쵡��b D9�����}��B��c�o<��E~��'�#�H�w�g��8��zSמ#43&�W��{�������I���@��	)�c$ީ�0��Q�,ݑ�D����"�2p$Y^��>��|���E����D�Q��,g �Cb��fe�3t�`��ת�ћ4�(��#�12����EW�f�}��a�(B��*d�ՋM����J�m��lŗ���׵���a���y��|W�V�
�{��Ԍ�c��X�j�/-4��}��b��Y�}�-��)W�Ҋ��F�K��U�N3�V{�X���Me8͹y�fE�g����~[�
�rWU%y��P�~ԑY;=7:L�Q)H�m�G,���U�Ò��>���l�#.�����Z��;�Y�"�?>w�e��c��-�c�`N�3G��0PT��.k�nm����׭�Ɯ����)O5�ӞO��w�0�:Yݰu�KI��,�*z�r�8�4Ă³�J��ͨ�q�!Y�����s���2`Z=��]�1�}�������6΁�<�e��|'�f���^P���foַD:���A�+�vv���E�(�\	����O��SZN��𖌀�.�;�e�ǚ7��I�U��&�%�L�U]���y�'�O?8/��LA8=?8���ke���?S7^#a18��X]�'��Jm���A��|B}�v����SB��G��������}T�j����vɾ�7��bj\[���h.��S��3=��#�ә7Α"Ε�Hcb�:��>5X��D��D,3}�6p����>�`����(J��E�������.\����:�S#�P�F:Ol�%��d�E��0��_���!��5:��j0�R
P���������:�A���V���=8n�=����)����c��"E�p��T��]���Ba�Mi"s���}�[b�F���jC�b�⻲�Ԋ�H��ڛ�0@��s7�5����(1Q{a랢`s��zi%M��5sj��*W�f��_�ʮ��B��Z|}D��-S�e.~S���FW��q���O�|^�%an��֮��3浼��%�N�dJ���c'�Vg\굎*�P��d�=��Qߗ$V�>:�iʥN�hx�PW�o�Д^-�m��&�M�+�%��2 w�i�4ց�����[�`���$��i���� ��נ.	?U+l	�8��D;��v��8b�VEa�b�&W�,%}�I�SBS:2O�qM��ś;��f�Xqb��}��FU����}s)�odO����H�L�?]p�y�B�.�E��z#8x�W�R�ٳ?����CXli��ͺ��r�B��-�C�?u�mc�E��.w�Xo�tG�p^H`��U!C��S�7==r:�M������N)�ؙ�:9^j_�tde��r��|>Rm1���>$\D����1ʍ�W5�g�a�M�>�^c��A�=�u��P��g,���`zJ�0��	3��<��A����`�ż>E��l���2�(�	��@��J�0��ϫ�{�e!�(���gv�$t&��J�K0�Z�2,�*[�/�x�W�N�=�Ϧ$8�A�\R����⪺AտD�����L)2��<��K�$���so�v�_�l�W�\�|v�n�[�U]oIa��Q�4_�}x�z���i�v�_�i���I1��a�u����P$�I��9�gᡝkn�,���X+�?u��_��3=���p�:�; ���'��<�M��h�����M!�F��'p�)�"Z�{ H��ޏ��[5���K�ڕT�!B&�}��/�<S���g�e�w)�˸>�al}��SZ_)5"��a62���?�"�w�V�yvT�Q��J=8Bf�,����^^� ���=������I��g*q���V�	��e���*u��`�ͳ 5����}(�|p?�9��� �fH ��2o�c�pJݺa"gLsUV�|��C������u�m�yk�~8�sV���T�pR�ۆ����,�Ąh�����@,z�$Q@�T�rC=Q�.�^�[N�6�>�b������&�s^ϓ�`��˚=�Z���7�S|��j��f?�Za,�<������M�|���`�C���Uz���gz��r j^���P�ԯ��L�2s���H{׵��Kp�=d)b+T��
��� �ƭ�S"���y,��	��]"��W'�;�ռ��_-D\��I�W�1� n�R�D�[>�ֶ�mrA�85�Ak�C��H�˓NǮP��YP(���D�L��@��{�?��Z���mC凵2��!�3Y��`4;V��֬r{䙧`t���J�ZgZ�,w,��Z����v}6\�'�i��]�V�R\�<�\Gx�#�����&At�ְ����I�9:��y�P��?:�iJ�JP�p�T��h%�y�T!H���zb�q]d��i�ln|499��'I�rA�"�8uE�l3F��Ij�-� $3�fp����ُ��"�7^�А�Q�Cَ��n�d������ha�k���CMHXʇ�p*��#�3�X�:Z�@iӨ��vPAo6G��W��&���>�8�p�/wN1��L�~W^��~x�T���r4`���ĺq `v��B�t�B����(��+#����4�+�{�^�|��o��5���<v:�C	qL|�E�ܗ�n�L���Mi�ۑ������=����Aa��v�V}����R�Y��[��ڌ}�M�y Z�2�#�wk�A�9��%&��FFG���@=�"S��S�"���|�9a�y�t9߈�a�ꩄD��8(�W��
'��u|����p����R�U��
y\&X}�;�0�~�M�E}���H7������;+��TL�����R
�^�2b�+���?�����pk2ϓO����)��
lgIp��G���/��Y�����b�~���_�%��(��w�;j��� ߕ��b{�f�Q��mZ�q�I5� r��g�ʐ�8>/˄b]��l
S��C�����uϻ��S
H�9�}�U"�p�0�a;���,�*"�&-C�r��������^���]�F�K��7}Bl?N0��W��p��5����f�P�)�o��A�b�0�ߟ��@��!�Ӈ)q������i�kH\�t��{�:n������Gծ}d4 �%�9	9���rq:樂y�R�����M�����ZL&P1l�����آ3��5�*A�_41���TŶjA�W���`��T�X�G�؄����)��|߹ncX�i�&3EruWsϐ�~JO�'�+6{ ���a������b�f����LL�(V��5��B��j~���`�v�F�ͅ�(������q��ռT�Z���%&E�����4s�F�	�n	lP-�F|ٞcE&5j>��y��&N^�{���g���y8y�}I/*��n p�|C�V|��f��%�[a��-�(0hޟ{xf�_V^h�H??����p�Z�8s��?��{e^u�K�~�m3�0P&���ѶV;�K��g����J��p.��>��Fh����J���ܱ��N���d���%���'��>�G �g�i��E~w��l<�5�;�0�2��k�%S�E<G$��O��A�A��{}aut��*i��Tz{T�C*���������56?�Qv��*����C��C�,��yx����;��t�P
��#��q�"b<6������0�����0\�!�����LܮBC�a�\�p8�{��>#��{�*@��"�S"��h�Ȩ��ԓ���5.	��j�'⛺�����v���6�4�>�Z�zS'�m�@[��x�@�Dm�?^��o�\_yz�I[�^s�x�ՂQ��/iS��CG�$J<-:���I�WV�ZS�yɊ�O���!ww��x��X��J������Ǯ4*�8��|w���5�A�	��D����l�<�J��ȑpسjR����6�	�2�X#��͢��qЛ��"���d�����x��"P�mD����t�����p��K�alŭ�A[1؄16,î뇌�`���?읚�7/�����F%��^���û��D{c��@пt�����~Ըܴ�plJ�l�]zk��l��ٓ�{X[s��o��
�F��tymy?v��4p���L@�D���� ��TJ��׮��L�;m]����4�������S������l�}��f����W�d��Q�Z��r��lj��a:q�9�g�j��v� 1_fv��C���ځ@�%<>��p�$$7��rC]ض��S�YG�U��pJ��CP�ڂ�/Q��6��o��Xc��?��m;v�K>8B�Z���ʀGm��,G�s��e��C|rA�\$Z�v������>�V3-Wu��*g�F�5�.t��2];�j��A60��s>w��_�0��/�｛�W.��G�]��ĎD��f�}��J���ry�u�sR`)�n���ɠ�H:�'��4joD�w���ܕN�-�����# R�x68W��n>_�ه�u��E�@�-�P�1n���j�T$���Cq5ġpxY ����ܓ<�E�V�7Y�+Yރ+Qk�k9�����-,���"x�%��O��u�\ZtI��`[߯�,H��|� �G��}ȶU;[s!V���P��&�x�<���a��?ڃ\�s��MC��������r�)���+�6���Ӂ,���tY���]R�2s�S�
�+�0	��0ݥqKx	U�z��|���%!�|� ���̙$D�=�bc�+����6����OO�<��ȫ硁�y4\K5�X��6�ܑ�s#Tކ+S��`[^������?u�5���#�(�c$hT+sw�L%���C�B���u��H��>,)�^�@��|�+'�_3���JA���x�8}�n��RG�Xp������U^w�lrM�O�
�`�W��n�hԲ�o�advFѮ>�oQ����-*�DB�i�F��Zι���p��u�T�%��UO�=񪿙R�lb�ᒔ�b'�rQ��Y�d @�QH��c��M�IK�2�&ju��,�
J��Zy�l޶��M�-ɥB�;�i���ի�О+Eů^�A��&��:�E��c_�Q����z�����7e�&����B�"2���K]iaa�}���Dlw̧��{�&����?A�5��90g������9e�W8����Ã�T���L���qO�/��=1����{L1NFՈ��wM_���>���������]؝�C��"8s�Β	�@2��KX��C5xk���i������S�ʑ;������2|���/U��߳|��ƇK��1C?��^�o# )'Ҹ���k�f>�q��JC�ļ=9�c~���<\�	/����o)	{�Z�>��v������C�"�l�ԚKxU}ئD�?���H�� �l��e���Z�s@�7����L�j���輁�Ȥ�X�h���(-�؅�$.�#��:���Ar���1�"���� t:��R�W�>ȨF��e����"�e+���xj��)#��=n��#�����}ě�6�4�\��g�!���KmZG���-D#�I�k��-_���\��&o$��O��S!`�(�2v�f���is����[Qc�p�#�vG��,l��;�|�D��j�$X���ə���E �X4��#A����:�L�6{�N�+B泃%s
��n��{yiu��g�3?����0;Й;�J�[�Y!����NԨ]�^p_u��X���.�m��Y����Da$C�Q*��x��C)����2/�_�%�
T��K���Q6~g��W�R���}�io�Z2�댮�~G&r�9�n�yp(ghm�Z���y�)��4��,dw1ZnyS���g��R�r��L�jS>#��������^�T.��y �_)��3��~�|\%�t�_�y$��C;��zWBz��x:�I�C����W\m��<t����4ʥ��x��=�H�H�YӼ#2���נ�Hڿ]�Fm	��-���W��^��g�8'/�)�ԩ#��0[8�&�Vr��!��kmx�;�H_��8��5��.��Hè�s���9攘���[�=�̯Z+���̫�^�f	����E�nv�w�rxD��D� 2K��bz��g��F�D>�F��
C q�[��e��e2"�SG���{�e��G�6E9�a})@.�~N�3Uz�f�D|][p����ˁkt�Msd�q��m׽Ֆ,��;ͱ#��e|�R �X�*�.5���`7�oƊ<�~'����Vc
�Ƙ���a�o�k{%�3�{O는\:y(��mB������W��d�~��
Աk!��J7���w7��:�K{~Q�}y��!ntZ�m��,�c�����ݟwi��G�Ǒ-��;�\H���6��Jș��敁!�%��@�!�?���+�t[�D�P橰>��	�+#�b7�$�!��%+լ��� ̠��MY�")(ig�,�ª��/�Y�1����.�o�iG���@�_������$�/q��9�v\�x
J����U�hI=��r��C;���T�t�$��\�̐{:��9O����%*V�̼��N�}�8&�9ÁX�OJ�g��tr��vz	uc��|]�����n��V��:o��}���د�(��E+��б��v�aH��g<<GU_xE7<���_�شL���1�
�>_q�g{�r�=����e?�b�p����L	<cW�x���aN������_mE�^�gJ����l���	�D��E˔���:p'����b��Lb���um��+�rw�Y���e�����������i�h�t�#�ެR�a�EI��@Z���@�_
Lk���]���}&���UD!q�Q0�-������CZl�0��֖���}����Q�D�B�g�,:��.�]˛�Ngv"�p�zA
��%�U��}@Հ����x#�n�#�ks-�w�t�n��;x�Oi+�,��&�up��q�p9�.���`��
>��-zv���o~ڼG]�B-2=fk�������X��0�P�8��a��\ù��?��t+h�S�&$��x�Zgn���")o>i��z���jq��19C!�4���Ad��o���~��أ/�di�,c,���5����L0W:�+�)hd����p6�Ƽ�~F��2�?��@��/;Ժ2���̓��q퍐w�!b�4]YhC���Lw�����Y�&�싽ٶo�o`��LNg�'���?�I�v��^P�{��E���W��O3�Y9��D-ϒv��5�:���mH�!�wey�W��z��!�[��.}p��Ӡ4I������O�Q��ܴ���D2��R�㜭`	_/�eM��yjk��8+�'T�dT��+\���D�Q%��L䆰;���ւR��(N{��bJ,��J
�[˺� #���ދ�Ơh���Š1;z|6/6L�k
4Ӻ@R�kRt%��o�K��Vέf�D��$yw�4�m�H˙�i]_��=��g��Y/ҤWW��#Aڄ4\�d6�2��g���*��UR��7q~�k�+,/,���"��VK�����z�TZ�mB�Z���`�ZsD' �$ڻ��럒ʹ�Y���ZQo��c����c84��6���u�5�d�"a^Ǣ&d#���¸4l�{�9�tKIh��Bz�Tـr�d�%��X!�� }�	5ۆ�O��K�]b��0����Ve����m�����!b���D�LE1������?4;�������$�F'q0$�K(LЊ�[&IE\eK��=�tc�?ͭ$��H�7����"ǟ;�P��>+ѵ=�5��Z_JԢ#�J�����$��6C5��&GxDU���26Eisl[���X�1�C�ߘ�i��J�c����q�9�
�|��<�s��nwv��T|]�	��N?���/�i&����
���r�k����Nx�I��u-�4�%=E�<��<���{\��\Ge���H�Ts#�$
���C�Zp�*ԟe�i����o5��LV�b��{i�_���
����q��~�;��+ȍ�S��p�ޛ*�z,n�R*���燮����>�'w��F�0�@�!YyC����t��7�[d�k����W����R�T>��ֲƛu��0֭��і
��9�a����妣j�D>;j���9*�Tb����/���o|��9��Z�Ԕ�k��bDQ�9Kbm|J�Q�|�ڸq����y��SN��Fz'5���<%���(JE���N4`�Ķ2���dKs��3u֬=��(��|���ԣ����6b��q��|>�j��J�)�����x!a��9hr��$CHY')ec뢩�Er�بF"���H���1�:y���ɏ��cW~V����
+���*�>��P~�I.�n'� ً��x�_�R`�{
�+��9�w�,&�s�cJ�A=��ؓ�eL������i(>!���qf �G�>�$%d����� 5�������q5�曝�����:��(a�8�;l�s&���O���BϺK�����aζq��{L�"!�Fނ��9��b�%�����g+�{�
T�6����:p�\�!w>e��e��KG���{��;$����L�B��e90�>߲��[�S1����7��6���R�� �!Ȥ�:��Z��>�=p��<"*����7m�~q[~�}7.��KhL���[���*���!�"J�`��Q��F���Um�����y�҉���θ����I��u��xj���_&[���#�[dpA�.�>�� ��V��p�ar\�/o�J^}�*�
Ȭ�4�R��q���I�c1�|��\?������d��(��N��7���@K�R�L��q�`U,p�_��C:;*TԚm�9��`���v�Y�0��f�x�:}/g��n�[��,#qq�k��RI��xC|���='�.�:Y/��k����>T��Zgd�(P�Ņ�߃�A�Dو���ʹ!HU9@X���i@M�N�T�#*�� �C�&�cK������ߍ
�t�<��7;#.��Xt����R'm��,�?��Q[�ᨽ�B�����Ӌ6x��e�؛^�IjWgMɬw��ԼP'�!��g��1�a�p�H`/�Z��׏zF��%�]�H_~��b�!�$(�v"N���R3�j1z \�:�r�1��;1����	�-�)��^�d�/'K���^(�8�@P�6? (C��n:-���s�\<E�GP։.��i|�R�N�6:�)�5/��D�/N�VŁ���6�sz��\r����<(�w�S�W�,q."M9{�=^z�C
�����>�b#*_���y��f,,)zvB2-��>�Ɨ�4��8�F�AǷ�dth�vlq]9���ViT^ʸ�)M��ʂ���i��v�RD�l���X�*�jP&��h''�+��=m�D�##�����qˁ����}X-'jn�ى�tf<k&��Q��E��k;�g�8���L~�z(L��-ʤ>z����q\ZW�W˼��OdŇx\p�ʺ�͋�6��'��4�`�a���Z,t |���m�Y7Ȗ��'�K²B&[�H"a8�h�{n����pn#�+��fK���h�A��Hp^K9�RO�a������]�h�����(�.h>>;l0�/�a
����
%�W�G��O���~��_�=�:���;M�X�
��^�Y?C~5^���J���篣��
�^�����d������V��p\c���p�e�2��ǯW9�-���"���y߆#c/G�(ΫtJ���Į�=��9*�L^�'��8G�"���7"<x�߶�W�/�Q���A��
Q�
��~���2�W*���5%~<C�K!�
`�5,�#�b��򢀙ɩ��w��ϟ��y��)���w��]��|ng�;�,�z�ݱ�>�۪$I6�M5��Iu߹c��c��<n�w�X���	��Ĩ�r��p2c���Rj�o�V~�ʊ�#pj!p3B^傯f�W̲&������\�b�����$@=w٤�!A� �x�&����}�<�6��b?U,ŝ֖�Pi���\ڀ޼|:��3�G���':2���
�/��"XWj�A.���-���ho4i�b�@��%|�k��xPQ�tno�)~����)��??T�#�UQ�v��ܿ�4���Qv��Ԥ�5<������g��#O?�s}�)�dl�}Œy|��FI���[��b��p��:#2��N��Y
�������܄�Cv=n雲 �0ԍ	�H�T�5�Pr}�b�0*;y�_�lu*�Nb\���:R�=W�r9x��ʰD�N��t�֡v�&�]�H�+����i��ˈc^��Qf!邰�"����L��vT*�4۪bs7�!���X��&����nF�:rT�''���şs#�z�w���h��m��4'��Ζ*���7y�zU"�i�	j����xZ��2�[T���?��� ��!�F�	�{`�3��{��g�>�^��h�S���|A�OI0�u�p�+ �^�3 ���,��nf&<':6�:Z��8-f�C5�ղ��>����^qe3?IRm�Bq������A�t�s�O���N7v�?��kʭ�m���g���D�TA���Y���O�Y�A�F��2w7?}3�oT�3m�f)��R:��p�1����f���b�c�4/]��-ny�����7�^�
���b,Ro�9�Lv~v�SȔٔ�}���D��D�Aa���!P3xI"ϊ�u�مQ$���("u}S?��9��.�h?�lu�ۺ���  0����gB�S����E�"3�񔉘�b�v�3x�d��p]��6�Ş�j��B��5���X��]d�����'�d��;nnj��z?� �e_�<lI�o����-�3=���՟W�K]��uc܎�[ �.:%� ��R��r`B����
����F��4��8��͢zn�-�I	f���!]`�Q�uo����Q��q6�t}���M �%�v�0������8B�P1��y>@$J/�-'�O}64O��a\�MkX#�(Vb%�:W5�I0��Xz� b�<���R����=��ֲ�-�75-K.�ʲ��[��8�@�O[���d��w×l`7%{Bs��:��<�����2��>�yhSSs�%��RB8�~й;�(_�(�a��CpީT뗎�@Ĥe������b����%lgxv�]�]�-7>��!t��T2@���[ʊƲF�'���qr~ن���LZ"$LhJ��'�6�)�<�#�X��ѷE�s>�"��g
S������(Η�.Yԟ��Oj�姂� [�������8M.�^�$�\8S���>�RpڝF�����ܣ=1zW��cNN�J�1[��u+_�'����n%�N3���+�G�N�k�>��~e���ѩ��q���S��;���Cj�VƂ�����\-�c���qy��$ l%,�/I�}�xs
��]��՞U��s֭��:��2u��A�3�c9��)լw`ee��6^*LB�<�����fә?2�9s������Y"q��!؝D#���ѱX2��I������Xws2*L�3 {3!�!݉�.v�6Q�*:�:��V� 	�ns|6"��|}t	#Jj,;
�1�.��}��k<��M-[����s{��)X/�J������k�1�Nv�Eⶂ��,2�St�j�	?�=�nkG��g�C�U���-�+A���S=�6�If�6��c�&�s�%\�մ6��%|�B���4'CvE�H�"}���)R���2�]����M
n���X��#������@4w�đ�$�a�1�՜{y�Dn˭w#)�;��)p�w��sl ��#�N����˝���I#��UC��������/>�^��[��ru�])���hy�X�~��MW@8��|":@�ďR���m������輰�����|I�<�xFO/6#cQ�@<Iz3�tuh�]�n=�u%����[yv�q�� j���yS,�e��	E6�&,�=�"Sw��5�$�H�-�DW|�0%kt
M��$���e�,,i�,�5��-bS�AKT2!�=�[qk�Tv����6��?�� Ի�r|���;]��`R����tW��\ ���#B�N����I.;�R�M�H��@�t�=�~}`�����m�0�>�Qm`^=�J˒�_���1.7=>o�z��\���I�K ���do�a�'�%;��%�q�|�H<�� ��j^��X�3���ȍ�BuӼx���澤��@F,�sn�hE�W��``HDt5�FF3!��92�+V�Qw伞\X�����$�m���G�q�P'��(�����d�T��+C���5@ ���>��:~��\��a��XsSQ���=P��=�����!F���~�������Tx	>t8���n�E�-�@�0�c�% U�\��%��}���=�L��r�?وзh��+8Y��Mf��o8��ڍ���!���\�����L��R�z���&����ԩ]��l�M�.�}�L�s$��]f!sM3�X[x�7�[9�F�r���bz�ƫ���/i�$��ws�-yS"ƏS0|&bY�
g���o���h���o�%��.���n�垉����]g��k���d���R��+���$��-�����^p�8�څ�)N�X-�1[
���A���V�,2�:̣E��[�����aUT ��:��KO�:�S:������ѧR��"��Z�\P�A[��R��K$�6�В�b>Q���(�Ņ���G��8:f��0�U᳈��)�)n]N�=�v�7,������7B�S��VJ�q�qȬ����X��W�SW��{�:���ZW�<���o�@���?�1m�F��*0<t������?l�g���6��`��>�%k��N��9O71�����+�N�I<p��$��ɯ�ټ4�S�?��E2"$Y� t,I�0��g��8Ɇ��6�4�����P�ɦ�-$@K��O���H���"Gywq�96s	��;�O=�e��憏�8mF�!�8� �"K��@�L�:?jLv��NH����J8�� �S;F_T?�]]:�	�j`�4���입c�ax9�$�~����ʭ`Ԏ��<$B>!��M��>�P	��D�o@A��.#�%��Tib�h]ssj�ώLT��h�S�yZ���>B�At-��gAD]�;K�ʃ	T��p2'_}���Q�x��
�+5ع'5��DIr�.p�<"�[�F�F�J�z��2d�*�CE�Φ��"��w���I{R�*���9�Z�Ͻ$�T�&_�ߔ.B�)尩GS
r�<&�\NA����� m��X��~@/��+:�� �`�	��y���Ee�:کh_:�>I�b;�:�a$@�ħE����8nJcR%zn��/./z�����<�o�?|���I ��uط�g��\-b��4,ԍ��Pv��|�}:eۖb������-E�~��K9
"fa
�Q)*��˯s�h��8a�Z~!\�o���c���w@ІaU�P�u�oALU�`�P��'B!���2���a�·�K/�_���I�2]S�./�� C��>�U�*bY���2��|`Z�<机8Z��q3\�\��Ŵ�`�A%*�x�0n|~�^&�fi�%��(�|3N6HLp���}�-|�p���$�'lJ(d��NQ��1��aSE�ɹ���zN䧕��q(0�óYfO5�+���]�3�p	g��x��}y�bKe�_ӈ)e!'gV���PZ�ҙbHM�zX���v�N(�i3��dS$���'�+�猾��q�Bc��/ց.�����V)���ٯ@g�[�]�CX.�3��|6X�J��¯{�d��uS�I�Ap�ޫK��*m�d��֘a����ly�Q]zX�10h\�"6\V�X�7s��ܕ,F�,|���NZ�f=h�p^�8�/_�q�[k]�j@zP��P(i��z��*��^Ѥ�8�Ղ?g��۩�>�Qp�$�_P	��$ѣq9M����W���"+�1 �j�@~���Ixm�-��VU�,�p�-���,���m� 0Pbf��&뗘S�Ւ*P0-��y�x�����;[mǚ��N�SN��]t�~�; C�@'*����qb<0�J�.��lє�F����6k�φ�;��f6�u)��2aN봞�A�P ��:@�gJe_�a7��4%8��Y�Dո�эN�v���b���G/��%�: �U��Tj�^BoPt�pT9�!�WI��{��Oȩ�E�na��A��?qJS�ƪ�����Z�Zʍ=�#M��%@��@~�K���0T7G�5��_̞�7�hymT����"�0�_���9��ő9v�u��о]�c]c�`O_����wSr�jrW1�B1;��8��������k�},p+%os�x#Óv�̒+���NVr�����n�V���[�`�d��̋(	�kxu7pcүx��$\���P�n���YMKtW���&]��}���h�`LÍEi�k
�)��9>�pXY��	�{o �1=�Xqث&�ŵ���":q���3������*��@����˺�i�Z�fD�k�uSe�t�,�7�f�*�
lla�
w��D�C�ٖ6�`i&r�P28���w;:֧�_��`^Ȫ�C�>�%<ɲ�� �"7<�����>K���;x�q�����?�J�.*b�F,��E���Z0
H�b��2"�ő��Ox^>�C4�-.�)�Q�Yb�:=�Ն��*n�CC
�ҹ+� L
��MA�tͺq���FP���l��߲�=2ş�Z���YDC;PY�^��`q�sq���X5P����5�0�0��ڢj�M�l��s������B��e����Z �N�?�R�U#wǬ��E���L�aܦ0�s�8s3&�V����ݠ�l#gx�br,x�MRئY`����@�vRg"0Uye�A��"?���	�)l:��}@�ȣ�vo����V��!��`rx.<j�1�-���Fhx^>*q=T���+���(�+�(_k�5��p�fi�"G0���9.b-(}�}�'�uQ[��(�g�m�X����b��̫���l6�>f>�G�Gh�y�$㎣�T��?V�=�Fy�`A�(�W=Y'δ��*��e��;D�τ�R�GM_ P���1���sH��5�@C��?����?��QK�P�a����kJ(y%�33�F�;Q9XOuډ��	\!s�*�מӄ��L�Qnfs�$���mE��Q����ݷ`Ckbt+��;~c�O:Y"�g�He�6�0���l,?��4qи�$��+�AFhѪ�
�g:���s�Mz>?!B�o�A��k��8xYv4/�DS�����
rzU�?�]/N(�C�k1��[��P8N��B-��;�n��i��������g��c/Rs�����d��7I�WfU�O:3+��E��O|.�u�~An���m9fԭYO�v��ױ�8�A��G��|���qsu?`�^�4J�X�)��XQ�D�����!%�^�C�Lx�ҧ�(��O��&���GB悡�X���v�a�a�^Զ֪_&�h�8E�Cx7-�*�a��8H�ΠL�A!VH�B+��'�k�U�8��B'�}OM$qݧ*��C����)�QW O�|��?R�iҎP�ax�Ǐ�)�m�R������;�K�v����m�^}�E ���������*�~��x9�����δ\�m>���Sk@���V��xPc�/�F(F�7���κT����B�q��w�_����	\�,�ք��?�uF��o$X��-u2H�V o��Zƒ����/�c6��U���k}>�Φ�F窕���I']���ܾ�5��OwP�ua��_j�Өo~q,�p�t�_�L)o�w�;y9�	�2��`�����;��%�w��;mf���e{3Ś}�7rfW��I^U(���U�T"��~���Zq�'㥷��~�C�tR�RIxN�b"�CH.rF�>�k=��o�8� �MY����p{d߉>&�078_����L���P��j, |㸋����	 ���1��Q����Q������ȸ�Z9׀G�Wt�d�-�����q8d���~At	ǔ��Ω�Qa�?��!�%�B�b��P�L�3�EQ1��
��S���ǯ�C�(=%���I|���X��@%�}��瑨�:Y;_���F����:o��E(�@n�^N)Gy�Q���C�U���s$Af�ar����<WG�_
Z���mhj>�� ��S�����g+Gz���IZ|D�c�Em�{��ۣ:�i%c��%�Wo,�O��'�2l&����	$��k̍�r��첈�`�-����	��"���[+����:u�y�?ܣ�����2:�eo��si#�w�'३/@
�����f����ɈU��¦	��h9p�Yk�(E�(�n�o�C��J�A;U2��Ԗچ������.������Y�a��.W1�58Oa-���m�J�[��d{��.�#&������hN�]c�O�B
���S��]�|�S���\C����{�J�����o�\�f�� �~��,���L;<P,րdءFH��R�Rj*}�(�C���k�i745�щ{���o<)$��=��}�X�gb��@ �H�����*���h�K{4�%���y QǞb�}��ɣ^�B"�$^$}�Y"�Ѽ�c[���gtHx+J���V~сh�*%i_�m���y�"Z1|������YS}v"��0k�:����p���Ֆ�Ql��ƽ43N짺�	.��	�����Z���`QW�J�rcR`9�<�Fs���R�Nr�Rr��A���k[���&�*H s.�O8mV%��F�ߟ�%�I8u��L�T��Lj8y&_��}��,q�T����ܹ_�`��A�~�1	Ӝ!�i~!�����ɶ;�4�DD����gb����P̷92h��Wہ�OJ���E���;C��	��qm��A
��e��WnWC��q��5�f�I�Ҿ��g�3|D��Wz��Z۰�lu캽4=YKiy.��>kA�g���Yn�3��`�P��_a�K�uÀWu��J`��7��d�g���)
"�/n���k�h�ᒦ��zM�i��5��Yn	������������䴘�W�����=������&�yX'B�99U�Z�68�����'�4��Y'�i]�}^4��s"�fs�x�=��Ig<7�#��a�9$:�c�����j:�����_Z��[!W�ݩd��o�3flܧ"����H�.��e�h�O��hV��lk�)�M����S6Xcm΢��!6�Ňܪ_�h_CжA�N/j�v�P` ���e�7���DB�9+�y�����X��A{~9 ()G����!+}�?Қ;��(�%��U3�����~���ynB��u���R'�.+��ހ���w���Jt�+p��a�=�Z;��C��~lQ;�=֫N��u'�����GّYU))Fk�9OI]DD�W�'�n}�B�k�E������٥�$�Wqh�biF�W]�p��R]�4#�R���#,�D���b����2>r4�@�}n2��w�����f8\�pSI���Y�)o�D� V�d��{V�$_H �ʆ��j���lZN��l� ������*tB+g���e_�h�"2�A�Z|����>��,��T��s�l9��M��GO8����'����jx/(��4����F&V�ϗ� Ɇ�������]c�q�����L{�˱��,Q�_�ѳr���ǽ7Cr��vk]ոڻ�t������')Z�77�h�8h���XQ ���}yr���
��� �i0Lf�o�=�Yls��N�G�'�aD Kv�q*t�ݳ���=��[��=z��q��eW5o/���r\d]Wy���EZ�c[p��[��逭���I�3R-�M�i�I�&Bu��*��֙�7�>��9�J���1�����}�u=0>�J�['�i7��q�B�Ά��f�%�����˴rO��#)��q�є�mnO�J���Aզʹ�8T���r����
 @+��Z�%��]�͓�1r_ �VmO��0�P~g�$�q<����^z]$��ʣ���	�T�h�!+<xԚ����	��A=��t|�w�m��vO>I���2r��/!�bO�C�*D��A��&Y3��oo^]�u��}�':�ΜjgN��.y���6����3��ȡ�w��3�js��l66���9�y��^AR �G6*zϣ���riQ2�$�b�+��9�6�����A�Z���2�7g��K�>�
��e�iL�4��O�C4�o�S���'���K��u���=g1/#��m��m/���D�.-R�M����H�LO���c�p=��K����m�of�ya�J�����H.Jls�Gٺ�P*���9��$�Q n)�������9FD*׽�<���!���Z��ǚ[J�8Ų��J���J�L�r hSr���'j1�@Q#�"e9E ��d�ѝ������|�#��s4׽������6��@c�.��ae�w�,��bA����j�iq��q�_�I�|�[��R����S���O5�E��O^��كZ�Mo���Z郻����.X��4q�Ejl�Mx�7tg쨇��(�-,��bࢃ���A��f�������(�}�6�E�w�Z�E.C��E�ʍ�HY�N�*�vzǙ�K��J~��fd������cԌ�E/.25�C�m��Oh�R �~m��V���ce���_�zJOy��ك�p�d��<g���??fS�P��н�KϣFe-�TQ[��_m��M
�Q
��fq5k�U"�(}�5�/�uO��L2�*N �z�" p/�Yv����	8a~}��� �}ϋ�d���HO[4B���h!�vI��E{�3�7�țl<5w�\��[Rd�_��0LR�����JVY_`�+�c��v��� ��$iV�C8J� @@YFS����ڹ�	�U�S�ʒE,f�b�"Q�\5��łR%K�Эc�bc�G.;)�v�Flή}I ���v�L���;+M�6�0Z�J���J�V�p���ga�@��@\�^ܶ�z�M۫�X�F���X��[�y��m�l�^H.$e����6,"70�B�+��K	���^5z��9a�F�q�@Y��TQh.�N�����R�X2���4V��y�Á�}��l��:���5��	R�p�)Tm���XT�`	�ݗ��΄
3��5��Y6�h�%Lk��S־�}�.�y"�XZ�
��������:-����jw��z)m�k��v�a�6��UIOW��[��a���xzZ@C�\�쭰�VX���B����*���9��S�G��HN	�jY~��io��^@���UwXc2�*�F�/��{��ּ�j��$^�>7)�s|�꽆cC�ܬ�@AԱǰ1x�G��M�~��]��c�胚��ߌ)���o�OygNO��܅�"Fq)����k�d�!b���D�>��+�f�5
�nN��i>-Ld�������Nڄ���MKVQi!���^��>����s��1�IqQ����F��9�[yҍ�>{��~�V�� [R�Ձ$����&瘆j��b�߈�	ݖ�7WH���E9 $f��?�m�e�唘��;�d��1�N�%�c�2�U^�P��2!F+$dT��~�qR`m�mO�|�_�Ja��a�B�:���`չȥB����o�C�0��c,��@����� �!>�P�6,�W�j�r�} u�W��/�[����0zSUp��w\i'�[���@��Mf(�3��Fs�_g<����_�G;�m���*Э�!R�/���r�7�U�
�eF�/9%m��h#���13�v�t����
r�x"%7����ć��2��x��K�*�����1�Ճ�[���R��k��Ԏ���?Ħu���5���Q��u�ʐ��X+�&��<� �L�|�I��L��$(�����c�q�׈dSg���0��:xb��QM�F<�����!5&��%��H��T��!>����AԇTi)I"d�+:���^��I���\�.��λ�a��u�|���4���z $�u5�Q��[E�%L�\x =�N��u}f�R5Π�=6\�����xn*�^���M�
�hN��ь��z��N�f{b��Y�Aȫ�+iM�{R��AQ UEZ��H��:vy��g�M��5sGoy~�`Tj�3���%���jG��D8�7��=�ׯ�x�-܎:cD�2�Z�Q���/
�Q��8�_>Q��>�d'?��6�(��h��t���-�t��A܊��t�4&�E ӮN'8�f^e�F�J�G�0EH%����Óg�]�M@�i�u��Q�%?i���@�p�YS��y��K:�lR���u$2��V"T���3,��=���O�$Π�]���䊢��uņ�'W�8��B���IRZ~7g��8�f���� �Ӭ���ޭ�˨FGKϮT�[��b�n �V��k��4y�m+WE�z�.I=]1�z,��6
"ж�� ��3���JF�y��c I^���b����m�1C\/����M	�p�;Z���O�U�G�ʧ�uP�6&���cD���{<K�g��`|�5�QKU����;�H�2kJ���@��^]R��J͂Ћ��j'���	)���V2���C?9%�| Q�ޟ=0��KH�~�u��P'3	�DC} �QD���\�o���ǔ7D��,[�C�Ja�X1=ZI��<��J��
24e�%�L�!\�e�׀e%�:�r��ke6��p�]ڝ�,�\Bu0��V0u��T�z���͎h�1�3��X Ȑ��h�=��wZ��R]r���-؍^�X��$s/)�ޟ]ݩ:*��/_��H�Fh�.ڗ�5�������A\M��1�T=�D����򴿭��Ia���"��G
�_ \_�1�*�_��#j���D�+��+�o|��VN���7��"��[��.A�� ��=0�k4�k�y�8�,Ar}�����=���v�2�!F0�����������c"�.jQ���7+@AIX�b;�<�K��Ź���r�v���d����NB��f�� 2��1;Ϝ)-e��d�e]۷��?�70-��)t�<ɾ*Q�~��^ϩgNv9�Jl�ZCȤ�8$����!�f՚/IY�Y5)���&Yk��S��LJ��$��#���l%=���ob]�Q����z9�[.(��Lm��R�y���'��G ��as����1�HX�<(|�H����O�PuDp�9�>�X��\"ؽ�C�L�R�e�ӽ`����N�b��#�h��Ӭ����*(��5z���!�H�R�,HK<	2F_��~�&�J�y�%r��2����cQ|� ��l�\��r��=�<�P�9�.t=��v�����_i@r[�W�S����L��"�hE�4,7��G߬E�0G���^�Z��-W����N�F�s��y��L f��S�8��3i�D������\^�����k������n)����:����{#�]��C����R�#>a�yln���ڶ�S�,0��!p��5���V춝o����m ��'�=Q��ԇ�ؤ�C���^��u�]v���}��U��x����3�OPKN/l[�(���p�ӉY���2����L����+�$8J�Ϳ���,��㹧�Uk�G�fcH���6}�p�Clp^H���br������+��߽�
�c�H.��^�:sw���`S�T��Q�ܚw�f����G�yA�wul��Xq��T�6���b����������S�;��W���K�z���ܔ=!0�}�@}��Bu^��µziL�U���ɒ���([	��/�����G-a�%Bݕ<�8�D��]%��9���j������?e����[�r#E�3���/����}���9�\w��d�V�*���Ep�"��6S���� ����X<7b�7��ǽCZ��6����`�&�{�#�a]{&�Y	&Ì�6��1��-�}g�O�؀H�� *�F��/�4��ʋY�^D�Ǎ�D���@Y#ˎ�Z*�a��`C*�����6.��S,�u�=*t��k�[�C��d
��2�!�GZ~���`r�]�t�f��.@zvk�K7 ��E
sW�|�
c�W��۷l�cںH��d�B��1ǚ|-P���!4yD��	1IB�zm>=1���.����9�B�"���7��u�܄��Fbo�ꊎ�'�g=����1�w��wY�Y��_z��-	�����<����gWQ`[�1N�[@\�o�C��s��,Wo�K빙�~ˣ�-�,�Gd��gܠ[�H� �T}��&5�z���NM"����V��_�.��OBI�>H
w��!�J��v���vJU��+p2%�m5pa
�K�ݰ�L�L���A�lu�j����B��������Pbt�<`�b�Q���9���"�ڮ�n0%������|�ݤ�im����-�&�^�3�V'®��nB�v�����a��f��:Ԅ5�T0�č�oבA���t|}���70֒�X?��?"��
�G��F7��۳�3a0�/�=���	zD��Km��&G�>N��8�Jd�a|����iP6�U|����R�ÕM�suhj�x�n*^a_�?�/��-�`P�M8�{���q����S+�
W`4�,�Ƚ�p��姲{,b���D�?<t���hV�x�a.�C	}uR�����4�}"�B���Ҫ�lr(9�ޥ�g;p��.��(��@������yE!S��v���끏�@H�Pr��/�-��r_o����K'd��� t@�>�$�'����V���w�syӫ��5s4y��vY��Yئ�gASV2,�8�^;o�1{���4q��N*�
�������O�Z�<{�~c�䙇�����P9��o�-��o�����O{э�M�A��t(>��$�+|I�kϺ�����"��@8<l�H�y\��E��w�%�3n;5S����*��&��#�{rP�}0��M�r��/�Щ4��Ƞ?��f�v{�/��#�_ԝ=N��a��#�2`��-CTD�+g��,Y �*��]�#s��oz��L�2���˄���0"	��]�X��|��Dy����D��X�L�P�^]�&v�8�!,0d�+�(�J�A)7�y9�~A$�M����{�����_I�gʡ���܎�K�(Kk 2G��yɨ����U5f�)�r:�~��m�����!�������M��u�z�?�5Hz���Y��M5Z�.~�s>�
���ѝ���������B'r1�g�	G9��;S��!x����.��;��r�[d�TNp�(3wE?Ҷ�ַL��8���Nd��L"�9 3a�I�� H�� �WOD�N��b���M�̒$�i�C�@	C%/춯s��������<p�1%�u8�\�˞q�kk�)��"N�`�lk�N^Gd0e`��YQ��A���	V�<]j �Ȃp�s���nW��)c���������k�f�ɧ�碚�삼�/�EI�i�D����9��?MvoU^њ0��n���`��;�{	F����HS쉯����i��G��I���<��Ѱ&�P��E�x�r��������G(�U��wb9��� L�JҽҌH^��n�VĮ�iB�d�& �>�x�����0� ���-�f��ú����h�[+����%�
d���G� ��!�����_2lG��K'�ne����ݱzH2/T;p�=��4������P��$�Bc>Q���':�p��=��z�1���&�����o�\K�?�A�qw|Z���a��* DM��%JS=:pN7˦ڊ�Eb�q��(��J�ۂv��{F��ر��@�%���`ro�j��1�ŵ������;�x�d���2���t<�[��g���1ij+.��:���ŰL���
��H��<��KBJ�H�N�H���٘�BO��dZUꇘ^m��/�Ҷn���,�T���_m�G����$ݴ�%��kÈ;�Ｙ^%��t���B�y'"Hm��[ʝ�R�)���|lXp�;����S��sh�P�+?(�ƸR��AM�����O�H��Xp�p���E\1����v��&$7O�4�*��# �E��{�4�R.��Gs�c0�w9oe$�Q���$P��Ȗli���xXV��>Fv54R ��XkA�⇖�F�J��6��nf��ՕQ[C���$���gWGV�'�^��=t^oP#�>��!7v#-:t�QC��<�M��D�xŚ����n7)ni{�Y�֮rM�!�D(�?�8�ҋ�%�cn�@�߷����;P��WΪ	!vg���{�Bb��[��&�i�<wz�2�</����<��[����=���Vc_}��hli�p����~��Օ�r-e�+����.�=�PRgi�?���+ëS�y��z��ʇ^&c|�g��/����[�����^%�u�H�� �-	��6d@VX�L�B�ŗ}�A��N�uĕ��L�8Nòs��\���_y����T�iB�,[�$����ە��m�zi��1O\��_D��ω$q"�9�)�v��i�a ˼��5�����[������|d��Vt^�g�p�ː<b?$�A���Au�S��b�	��	`����#���#:��W��Zq��&���{V�t��jĻ��i�w�(D��k�.�o� ��}y���
�Ŗ��E��Tꛄp���B�r������.�֕4�dh*i|��Ҷb��G�L=��%���o��עȬ��gN��c5��.��ސq��Z xCX��=`jU��1�B��t��cwP��XjGR0�F�r��jN'�cPB��2-憗K����h���m�LAk��i��^�����vW�'�P�(+���`|D?�{���G^ƃ�c��U�_� �K���<�r�VR���B�%�����5��SP�o�֭w׽ӽ�nad��ӗK������־��`W�C>Z�,��W���^�{���Oꠔ%����vb{l���G鸌�G;tv��m�{� ״>u/d�y�`�X��8������d��0U�[=#3d���%p��m�g=�c�eʩmO�������<�䈶�s�A-]����!u�0��ف�O2���h]�c����2�jf�G2A��
�dD��@g�t���ʽ�$��?6J��>����i烪�%�.9Fx�^I��Q=�Z�g<�V^7bơ@=�z
�ԁ�K�fD>|3n�9b������d-�<����ָ���%��([.��Cy�{ Ǜl���%_O�ݻ�ŸD��~����V� �����s���	�tby;v�(I�w�M�����thJ���֧!\xR��x�;6�g�)jb]�2T�t�$)g���2�P��C	-�S��-N�W�u�vC�?lo��-��� ��a��5U�@`%� ����q��:#��)e���M��R��ƙ��p�xL�g$u׏K�`��g�>+�f'ǁ7*�,	M�U��҄F���D���(�.�q�j��a`��-��r�I�dw2ۤ/���9�?׽��	��6� �'��':�&ة��R�]!T��&�qw����,��a�QV�AßBt��k��dв�z������刴r�mD�`"���Rߚ?�ɡ���͝���p�Y�Z��t�Ơ\��4�-���M��b��+�n���nR�⹅}�P,��Ga��ŸL �!�\g �w�㝱V��s	ˠ�b�N���ƥ�������#�?e��;�d0�)��!-���xjKfP����vJ��]�^C]�Pmv�t�QO>1��e{�_&�9]�$k� ��DЍ�8��)�f�k��_��ɓ>����q~�0J7xύ��_	`ۺ��b�1 ��:e��[(��U!3�ݰ:m�h�k�aB��ߋEt9s��-؆��e��1�zl	���YM�$��C�4�Q����`����eL��]R&�E��1��8�I��v�4dxl=C�T�� �a�0f}<E.f���v��Y�,��[fKL�O		�Iy�bӟ�4~h�{#2m��Ш��o@<�L�j��uKW��s]�=���z����Z �pV���Q+٣��<B���kn�cɣVE����+'�J�t���m��Β�]�a{��%-��Z�r����`Qt�Q��(�����?Uɝ�����E��G�Y$��0N$�,�� Y�o�D���1�߲C���wɡ�����kH<d<	�zz�&ʉV�mY?YJm��A�����7��? �	\Vή�0�����h%���'0 4-Q����7�R��<'�g�3��sWc��5Q�C���Q�@�U������ k����(mi������q���S,n)x�O��rmi���_��x�'߂�}s�0�J�IQ�UqZp7�b1�;�Y��ȹ���
��i��?�Jc�-��OȦ��t0bKR.�-��tc�j�}oN0���~�\�ݣK�Nr�A� ���W�HGG3���(	�0�h1{�Z��4�!P�B�z�E[SPt��(x�O��Z͉2M�K�n'gaO->������,��@��� X�����}w�-�/Q�{�d=����G��4���jGY���!k�5ÜT��ڟ�����ی}F��7}�0��+d/�8��C-a����.V����N�e,P�����!�.¦w���M�Gl�ŗyċ�2�%��=�P����v��-j���n���ͽI�𓃹
,�_�t��4-������0M�0q�������)��P7�(��5D�S���`�.G��^L�!�{�AR��U(	İZ����P��x���[����XWQՋ�G�P>X�M?�wnp�S�H�F��{�y�)$89�L�v�����1�&������kX*j��etA8�qxS琯��\�I�pd��0n�f�K�j&�4����!���b�(X�q&�Txd��\D�|߁��\|;5G�jg�8�߄��#���+77�Of	Y��ѐ�e�
Z	8Q��$`��J0�~/�T;h��+���3T�k��9c�R��� &i���3��L�iw_B�1��. �u�I�xD+�����e�=�x��S/��d�@ܬ�g�D`�u�0���i��=t��T������M9�fdP�'�.K\��~M<��x�P}^"�]�"<(����)ة}]t��-��1�%
d'��I�{�����a!ϰc�/�-��0���Gr\��B�]�1Ғ�|�ItGY�U��7�e,��7��*�!-�*���eP�����@r�S���R�
[U���9������@����}���$����Q�^�pK����[���ܪ<a��y!��L\��|`��;�����]H\r�!T�+_TH'2/��$�����'8�i�*J"��e�Y	׮Z5_$�b�Q��1\_(�
��K�H/kC��}d�-�ML�3���>���#�,zS�w�V_2:�kZ�H��3��"B9J���p־�[�����V�S�(�=�q��c�{��x!)�PE�����K�����g�A~]��a�&�#�ҟ��>�{ M�jʹ���N�M@;���:1- ~�U;ȣ ��6�	Ζ������<;&Ѐ��.uC 2s�����`w�����5�2�!h�w�$�n�|m�Z��:^�ƦU&jg.Z�?D���bac�zm䛁bS�2���:��:5���b[�����v�� N������VX������ǉr6�]��緂i��袵E>�67X^���q�Y_m���y��Et�T� 刧E�g4�e��aЯ6�
�z�-��.������7�ϗ��2����HOy��m ]��}�T��!�Z�S�o�����3�2B��?�}}�&� �ڥI�:���T�KzA�{K��rD��{� ػ��17r�� �ތ��t�KP[�F{�d�j�R���.��	W���/Qfb|�a������(\޾>����SuՐ�O�-�:M�����|@�p@�;k�"�t�c�]j20�-`�����K(fi�Р� ��0ّ�(���P����#���)�vqe"�������I���-��H�R����x��-7O> O��9C:.}�е��O(W����L,3�����(�dō`,�j�̭�ֶ�e�@ܿ?��7������p���F�3I�@R��m'��+ B8��b#���4�:�d.���4A�d�,�*I�}W��2��Z��%�)
<�.(ps~�g��O�(�<�� �:��qa�P7���#�94B��~(���ܛ�c$zƫ��9P��}��Ip�a�,��2Bj���p�c�h���֭F�ё�n�<ڡI��O�YIWEn{�G�Gps�|^O��ǎ�P�=�{\U���}}A�% I���\'ǜ��9t�A�I�����1 ����Cpn���Ԩ���_���{���ի��ۧO�������KF<���wD�Q��r��i�쨃-�ĝ�Hې��˓��: \p�sO�i���L	Ԕ�WD�#~���o[B<!�-�=m�F��ψ���a����IU;Nޏ>�~r�H$I8��c]l����R*~���m�3%}NY^X�s�g� )��A�Z��V{z1�H���īn no?���kơ�~
�O��"ژe�5v�Y]:��yx*fMe|'5t���;�r@JA7P��cIR=�}��� ��[�N�
`�ո��G�K&lOCB�*�F� UZ�s�����U4�=$���ڧA2�,�"��-�'�����i�Ao����M�����@\jAM|[$>UW�������]��U��7�sV�h�ʌ��.�����<C�pL}��"��c�Z������Kq9��(�⮳+r�&:3dME�4�Ǒ���_�l�����	T�]��(f�R���b���,��]G������f5ڂC�A���:'?@���2�]�R�R�ݙRx�;ܜ����[tC�54e���|�q�nOKG?v;s�R�����Z�}���l3t_��fI\0����܄�H&�q9�*�IM������<%~,/�� 8��9BC\�y\�`�q�E���'�kp��\�L�_c�j\;�1R�3��#����,(�-�8c4�mLceo:�?vo�y`f��vT�ԂQ֙^&��זt��ݛ�{Dk<�h�B\������/~��nH��-w����I�a	�[Hu��<��?�8���t�b!LrOWb9d����� ��%�4Q|��`��K��(;�`F�Ȩk��:�[A��TI��'E�`Ĥ�	�M�ml4�@�����݂�*o[�j�ђ��AB��o[W���Ħ8��
m�p�������nOl�+GP`���;6��	�.��`ক�;�������Y=����NXa��!t�h��]��ԉ�<v2�v����b��%�ܘ����/|��W0�+_N���XNeE�5���X�$�[��/~� T"|����q�Moo��|B���\�8��Ԑgl�<���m��> Ln8p/[����ڬ#A�Շ���
�3OՋx�
�L����+*��oh���
|�����"�;F�_Ng������-i�Й3)d�f�۴�!�4q��a�E�#��oK=%ڧ5��8���N��.L�᤼&�{$��E\ޘ#H�HԤ�T<;�C��Fw ����Ҭs�@�:��i�0P��-ϪGn�蘐ݒ�Tg�Қj��u���
�YL��&A�t��s3�g�bg��>��^����p�g��j�O[I���V���J�.<�9dhrkHP�s������ú�7BÇ��晭���ת�@�n�
�B`h�#+?���5tu����:�³��$:�w�<%&��9v[ĵ�4���H�e����H�P$Y[2s��t'gJ�O6��KA��_�<P	�y9�e���r���6w@.��r8M>��(o ����p��r����m�q]�*+~��j&uE�s_��&�������=�M�~� �B��/���/��j�''�Ru�2[N3�MMr�~��b��Ό�ܧP��6�� /{pY:�ȥ��^AJ�p�k��~BG)Y�A��s��s������@ i,�Q�IH�V�	�j���k$q�`�bu����"���O��;�{��T
-�X1`��!����}�y=}��d�n�D_�㷘�O��t~Ӛ\Ϩ��5%�\-d ��a���72��d��藰�т�a	c�B�t�v�NcIs�(a0����,��^�#��ЌQ�{�vvp)@���/}�#�[ؕh�E��-^g]]��k�y5S�NDJ/��.�@nM�|�dl$S�Wi2�b�d��J�6t���'�-b̞�pE䨻L�D��c#�{aEz�{{�/��;c��&�R�< L� �#��"�2��A��Zb&�*N{Y��DIe`�M�%K'���i��yɪ�������K�u\�P��L�VĵɆ��HJ�RCn�$��5�^����a]X�t��cI�!�}�JH�k�,�v俣���:��U�ʺ���s��Ni�y��5d�fZ���* �hn/�Ŷ�ɮդp�,Z�Ш��-�����lV�MᒌCK�)���Y�vy�a~]���-%Ф?���(�ő3�)��lQ�Q%��b�X[�#[c9��#X&���C�5�=a�r6�͜$H? ˼c`9��q�j�G�����%t%i�Pl�NDPY��WǬ=zP��Z�b��T�=�b�]�]t�G�m��7�t(����-L�(W@c�x�Xۤ�r4���
r��-��ga��W�Ө<
ڛS.w�1JN�*�|�B�n`5��q���"�Lo�
���;5�)��C!��U��cٚV;EP�Zhƺ�C?mL��+3g��Y/��	-詔��9�Ҡ*�v��U��ӈ$>�I�e�����A5��\��h+YF�Կ}8.<�[TV�J�AD1���xS�kV�}�*@�}"{�gh���´G=�N1I�	&��S"y�܃e�x=(������H��p!l�_"����x�P4?�g���e �Z�8�ڝo�Zf��81H��0�����i!ט�I?��o�Z}�Ew�Fe}@����˙ ���gHtt3җk�>|V��D����v���$���Ҍ���:��Z+Q�OŴEfA^����t��>RE9��2�9����+d�z̈́ڃ<gn�~�Ά,ܘ�U�4��\4X����}�ϭu�^�����S�$�s���Ǉ5 �, ���
��ڈ��"K�l��<hX)'��0��g{��2ܨdnX��:Wy�;jS�'<�W�p+�|��2���� �#b'ݪ���Vܝ�����@qɥ�f�Z�r�R�����&�#� }�8E�g�:��N�?2�cryh��sft��X^o2m����=LV.?��4�Z�q���o�e�����b��ݝ(����0�+:���}�#���jt G(��y�?�lv7q�.M�a�����@mq{�w�gc`��^��y���tzA����sWǶ�E�͞����$�r�Ȓ
����U�
�����
�u ���N�Sh���#��z�N��~���[-�:__ ��ֆs����ۓ12Ja<)Ɗ��
H�P(G�<�oz��+��	��bdsv�a����¾A
�'H?3CD: `+j����s\�r�6 3'�W��XR[��`�Pn������\%7�L8`p�)L�4о�dE��V��~İ�$�.\}�����H֥�S���%#��`���P�l
��y�M��T/8cRa��v�I�C>��Z�_^V�2�n/و'�߭\�"M)��p�[D���h�����c/�(��89��u'�n#�����
�t�Ό���/ǳ�8�����$�����q����y���wv��YW�%��	����)�u��:#䯊f/����B5�D�X[G"�� �֨L��թ�񺎞��Q�I��?���Y=������FQ2��a���=x�f!��[����|c3 =Ӌ�׷�_�$�V��!�D�%M�HF����7��.�c��C���gR��'蛶��<��e��L��^����U�Q��ePr�q��O<�H̪'�c��@~]�v��oiܰ/5���?""��/�=�DFIMy5' �e�{��Ġf���y��%���II�_��;�Pz���u��M}ML��t��U�b�?D�C%�-[��d?�J�dɸ�ƷӺz5��T�p��	3c�a�|∕��ЊN��x��Q>׬���������
����#�{�0X� yx�ٻ����p��2iz-�M�u.��-͋����U|�8��a
O�	L���̽�??�Y����a����Ԩ�I�k������:�Z`��\�zz���z�E�~�9䏊s�Q ��a����V��:H[���Ȯ�0_�(鳲�
E�����R�%�JP꓆辸�@W�W��e:`}v��٩�p���z.�}��P���q�ͳ'V䳞��4��'�px f�c��e�#��nǩ��(p�B�.��&���}�޼aH�}���=u���6l�@7�+���rc}���i8��%Sݨ���o��
iT^���F��&���^e���x�v�{F�-�ę�h��6�
;��
�DW{!�̕x �΄��z~, RQj��2���E��%�w�؎f��I���ϗ���_�j��� t.N�R!?b�5�!������)?��@�3yY�g2'�J�%�q랶���aXp[�M�X���Ra�p���%������n���&��ƹ�"������LEk;?�Uv�(\�?�0��_��C�;�:Viw��I$�j�g\�����|FE3B����w�ߢ3>Р��S��"m`cu=1	.nh���*��b���](��G�^���D���;k�A�ZFE���`Mf��ͼA�v�� �/�c���b�J`nS��*N�0�NPD�ƶ��ז���C��;Ff�`X�$e���ߝňED�|�3��k��KŨF8!�SaZys{���n���ML�����H�[>O�V2��E���V��=Wa���l��j��LQD^+l� �@�m`����slz�������	����������>ȶ_�u}�k�Q7�q����p���(�l�ąps�9��V��=��#y���n;J��H5*��7>C+�v26b� :+�-G��0Q��V,4%́�0-���!bF�w $ˑ����z)L�W<1�M���)�i돕�yJ���r�����xϷ���e�({�{
�`����M��Iz��-*��w	:)<r{�Ė!j!�a9�ΝO@�`�Kϻ�yܕ��k�����DT�K�i��P�a�����Q4��e��a�W�C'cS�X�pX�i:���/0�+��sO9)�nK���p���@\�X�EV9qjp t�R�����GY�YC�$�o�F�
�Qi�oM�`SP'd������r���s��z[&��sb�'��aVm6�	g!&\�h���2����c� �a��H�ޔi��}���[:W�pN#�S�������W'�-�Tgޘą�0�A��|�y�	�b3@̡�Uѱ��=���#�=7בu��>~[�:��}�e��^j@r�DK��*t&Ĭ��R���=3:f*2�\"D��/���(�����o,f�܌���2���o٧�m�9"����O ���(Ry@$?�kZ����!�"�`��H�"���0����:����QY,�D��c'���[-��eC?2����U�?ٵPĊ��e24ѻ| ��T<��8X$����;�'7�/��lk��=��9>���l��S�����ڐ��� 7&X_k��j�C���We�ft&|[��7���hڔ�?w��w��8����{uvWrͩǌONt�}�Y��bF�K<��2�
d%c�x�?K�����S��ţ�nE�9��R���s�סƊ�+�O�х��M���^^�*5�pD�7�I�i��z���~���U�mo�V�\��	���2�c�D�c�ϒG)���m��ݗ�pr�W�W�p:�<��0�:(�jG]��9D޲�<����F�
�C��6�Goa�L�!��"���"FUo"��j��O���<E���m6����_�(e|��#�$x�][/�*BvŅ��Bm@�3�2��.���V��3m��|f��Eǯ�\�������Bq`%�,{����E=C,�J@w��3V�>�S�#��P@��֟�B �d�m�0��S��>�w��{Q�t�p�Aۏ���T~^���k/�2��۰�;�0T�EI���T���W���*�m UlE� 7��~;��,���#=p`<P���?���	e���!�"C�sP����lBq�ǀ�8��C��3y{���A�hϺ�B�?&��zr// ϣ�xj�w���5j�x�3c<Is�'/G�&�S�y�lz��k���̉������I�O����$?�)��]F��!�g�v�D��Si0v��P��9%�D�q���R��77F���I����w=�'����X�p��.�B.�8RM�b�Cv�+%��\[cYuyz/����Hh�}�ec\9�2�(vEV�?Pƽ�'G�����㳊q�u��cC�V;�vҽ�)V5���;��dP�%pP9
�2^5�I�{��)�䟮����f|�b�F4_��o��d��h�t�h��tE���$����C.����y�E��<��T��u!�}�Sf���2����Ѹ�N��¦7#K�,��7Tf#���3�zu��_Dy�$��p۶P"��j�H�\U�ʃF����I1M�����G��3 	� |ޝ�}6�&��Q����w���^A OPA}��V2��X���v�tsF���Y�!=�#�	1 r��;@^8�̗j�I�������|+�xYU/�.^��,�wR�U~�������r������{4�V��$n���i�L��*���j�@{�+C��6J�zm�yc�Jq����c�r3,*�X��e\b�����z9{녦�����hE��Ծ7�;=J��$A/��Ca\m�O���ɰ.���N��	 Vr��N	�6�~���	�M�[�/[���o%��φ����F���5՟�/X�n��l�P.�qV�U���������|���<�+�׭W�?����ұ�Ķ�n��X��t��Í��Q��/dܛ8#��W����2�t'$�ǋ�{�<�b?Q���/n�?�l`=@�j��d�����FPa�_�Bh����4A�A�T��]\�[�u�)�Ҍ�r��7´�;n�!����ػ;�:��X@ε�Q�-U!(6�^ϲ
X��}��ic�����踉��_���2P
"FB����Ch&����72��h�=Q6��a|�qi����]���/-�WY�����tLl���A�yu���zbf=�V?��UN)�(x;p@�x�uԛ]�a�p0�؜�f��ֻ-&P#��Pnɡd����|���D31� `٠5[C���H��2(�: �����[.������I?�9�Y�2;�Z�����`��2''>�p�F���Y��\������1/8�W���e��񶭄�|c!��!��ҫǯ���(�N�µ�:%H��@��[|���ܮ^����;倖�����g���� :��5 830�0��1a�,�ʈ��5�$Lj���Lt_|�tv�zϸe�N_z�_/�^w������͙�WŸ�h�)�^b�ϘN������"W(/YN�ٮ�=R+¯�%���F9����r�̑�(�F�����2��U�����z���Ʒ��z���ձ��p�NW�7d�ȿqx����`��[�����Yd\��
���9�q�h���pf(}�'�����OGF�dNt��5��%N�ۛ �Ϳ8Fϙ&�A�K���D�sU��V%�BgQ�Zm�vF�b��n�� 5$H��`B'� �T�]��r�B)Y_
��?�?wؘ�v����y�x��k}���<c�X)���/���-�l(�t�-�����#[�7��<CF��2㈉�FJ�@�����e�v{�ClZ�7p@��z޷Ʃg��x�o��l~��`w��U1�|���TxJM�g^>� �=Ņq���w^Y�v']n�{�����b�Rf��F׉w��Z��C�<`iIO��t��>f��Z0�ʡ�E�<��P/��y�w���*%tX�H)�X���5�(��7�1�to��O �Q��Ԣ�T̂܁��&-挎	2���熴�&}�ٱ��gr\	���� D����F䝖�]��kFĚ
v���iͨ�EL�f���^o��Gۗ?�=*�[��%Y�����O��avc���^�q!����@*���=F(=/=�(��R�?_����׺�<IY}����i
��:�S����@���i���ԡ�3&�����T�dF&��z�!#�ؕl4�7���S�O�ޖ�.!�K��c'�q?3~M�S�$h��_�����Eɏ�<d�8Z�fq���5p����<�M�p�o"�sT">dI�>��{*w9c���{��rV�������O� �q��z=�]�����r�jփ&��
5�F�Z(

�.�	�Vg���_*�/�t�xʌ�v�C^��6r�Ɍ���:dk�L����H"���;
o��� ��(�	X�|L����V@[C��d��n�;�r|��-�\6W7�ha�3���XW�/%!�a-������ʚ��H~�!�B�0R��{3�Q�#g�:`��B���Lc1�X���e�U���hL�[ƨ(�z�!.�}FA!����X��7u�g��J�UbEr��0�Y�r��&f�ǀ)ņ��袨h�Gq ��j��`L��k�JCV�")��GCu��JiC��˸ 8h����-��`����D�i��oM� ��k�N���Qu�Մ���̰!D �O^Tד��e@#C:?EX�%x�S��J2�����e�w��q.ȾdL���o�MA	�4w����]�]���Py�n
��P3g剌AWv��PӮ$\Et)�_�VF��M��>@��5_n�gD������t��\/��U?����O(�P���������i��#�'�Q��R�oX�E�jj��,����o�cpUM�t��|?��+�xC?g"��hT��G����٪gXO6~u���!YOGW<`���);�`�EL8��>���'�8�f8a�S'}P����2��%�t�u�l��Dح�g{�~��6S�&�g[ۼ�ƣ��gÜ��| ���*������O�/��	 H1�u��bL�igMFdh"x��~K{���1፮T�s�!�����ߞ�#��Đj4��Dj�ɤEp�@X����ݱ
�;;�.��M^�K�>=�Y��[�/<b,j���Q:N�P$|��N�ɚ"�$��D�'�@ӭ����]\$�`�DG�$����� ��Ӌ_�U��%����j�Tl�R��M���j��w�����Jvm_(n3�(�/W�⧌(�x/��ay~�T4L��US
QF��@�b	�w��?�Y�҆�e�BE�|��gg��6���5���]��ڱ��T�q
�^�k� �<<�����Gq>z�;�����eQ��)
'@�m�Z�������Vs��H�͋=~Ha~S�	JZ�A��t�!B+ �*H{)�%3뻎�y}"#Wpnx�U/�d%�q���ߏt�f�w�5H�GxH��RP�Ώ_��y���%-~�#Gq��U<[�՘FJni�R��B78Y�h;�g��rd���O�s,H���b�H����I��PN���=�P�\P��W����dsuI��C���)ȏ|��3���>N#������F�R�j�~���dZ�e�x�s�π���Qoq'ͦx/�o�3y��gt��~%D��ޢ3��TjUkZg��բäS��@u/�GTb�cO�F���ө��Dm�P�@�ʷn�d�D��i-$�;,(���f,�q�屑#i�9C��v}�?>Ks鈝��e�웫,�`�Q�ѧaԅ�M����rϖ~��0�YE��}5N�͚�+9�0ǽ���8�*��d�|%�����y�j8*��G�x{k=s�Y����+~U���~����	�9�8p}'��,���%el��W�δ�9�}�h�H��\3���k�ղ����Z�K:#^X8�rr�l�ǀ�15=����玭�7�eDd�\�^{�?(dL���������S3�_7�M��z�*�2n����8�0�B��6��9�pP|	�5.B��\MS�噆_������y�٪���گ#`��(��K��V���Ov_�%~G#H�A��K����ې4w����E3�"!�9���6�u;��8�ț��~�\�a��{ƴ':�1)�
d�Ud��«�X�&�o4�sÉ���p�{w��JO��S>��w�܃�@ �t��F���9��"��r�;1z٬����뤧Y�u6,�;B
��E�O�����>$���b ��?>��m�����	�>��1LY���xƼ��i��C�j�C:/Uk�y����S�ob�&$��k�~Ā�-�܃��XUܒţℛ�ބ�K:�QP.��
�r�-��j*�j�ל���Ay8�/�����v �S�f}\�6�uHʀ-tN/�_%kڂ��k���2�9o����:�s:��۔�U�R��Gì~e��m��.����T�r������kP��糁 �G��ԼRQ:6�u��%�$?k�����\����V@Hra�����Z���s32�1љ���
C�<���G�#�*���-e;T�Wk����;�0�ut)cf ���m1�Gs>�]�Z��?��4�͉��	|^J��{��<.|�d�ڟ1���̊��;T�wp�j�
�F������g(Qj�_��M!;.��6���8�r��no���]J���;�.��sy�S���$(�������H�sP:r���SB���H����3ȥP���^V0_K�ݕ[NX��ݢ0m>�LA� ���D����xg��mX�;�N%�M��J�ӥ��N-U���J�.:� 9=��n�h0��O��H���2�b��(�{��Gb��޲�ȉ���y7xpl~����Z�����ь�7^
!U0L�J��$��@��p�����N�M�� 8rV8w��3�e몹��dM�۫�ndrz<�G+l$�q��{5jr6P�w��|����h��Rz�(P�!R������k����ٺTZ��8���*[����%�3B'���0�P0if�T�l"N�n�i�ı�Jy�FQW;G�ۭc&A8?s�y�0����A?L"���1:���@s.Ƞ<�8;\Y��ހDJ1�5������.�� h,��e��p1N}J�� >��5/h��%���A�yPu�DƦ�?,��Z��]��q��6�ٻCx��W�S�-����"���+(&�A&{�KԷK��G����U(>��u`:�e�@cR��O?ں������I]|��k 6c��Ͳ�?��/�/��T��b�E>���~,wQ�Ԗ�_�e��\�Jn^%�u�q!<�U�Ȯ[� ��9޶��|�F���6�D�nt���T��w�ɝ�Y�TLk����Q'i�uv�� ߂OR����Y1ؠ畁?�֢}z�cE\�*I5�yZ���Ay���]�xe��	�_�ʢZa�k�k8&(�U���*��?Of;LW�Y��4���N�����C����2���zd)��]׿4qh)ZzP�_�Q?���_f崃�i��~
�9ǎ8���|��{\W۞;�W#�!G�P1ӧE�+����Vx�O������WVy�q��^�?yn��,��K��͟�Go{>��@�JR�l͕�.)c�y�:A�Ǚ��ّN����R:����6�'�s�i�a'��������j=1zB1�?���AV�J�ER�ջ��z:�! "��~�vF.*w���k7�VB;YHe�(bP����k���o��'����t�l��9+zЂ�p}0�9cŽ���^�-��V��w��珩PL��j2lJ�)cV3Y�_�yd����N$�w�)���C�3�q�C����=��8fA7k)�?4^��?v��   �菹�B*�X��H]�^�Dk0���pj.&h%����˥�����涳3C���T�p�*|���4=��,I�>�Fܣ��u%�L�7\����G*h��]eW�X������g�Gb�$=o�]������~�^�J�Ѐ�������cғoTmŗ�В2�~L�P��?��eߤ���{5dhOV�=m��^$����C�EM��8�hU�^Ci=~��o;����eU�T����:e 4�>�6���40��Mp�t��3�n�5G��7��q�m��B)��ͣ��(�}����U����sGk(�qZN�F������r$�[�:xm3�&k������IB �$ǿ��P6��U�L�Ti��K����$]g�6z&h��o�Gl�#bw_�.Q��Z�g7:���~7N�&r��i�"��ĳ$��&�*�d62$݄R6o���L�ZzRCvu ��h=4s�O��K�/�@��f���`���	��\��S�i�a���@�̷�{��m�q�ِ�ۖFI��MN��N��[8�l�a �~��C��s��}�a��)[�����VN��Y��-l��Q�vH>z����L�X<��"�lk��ǹ>j�@��T?E�-�~�N�&6P3^��@�M���Dl�� �8�J{)-(r�@��7�ш������޴�-�	@/��D_��7a�'���u�+Y��O ��TLB��ÎI����� �j�?zs|�߱��[�_Ϫ�*r2��!�,�|�ٰ���a��%��01��е>b5�O`V̗yI��)c,�x��'�� ���$��"t����s�x�q���
�wU:��4 |ā��$m�amo�KV�R1�U�wlM���b�V�z���#�h|�h�j��}�%�b�
��i���n��\2g�T�� ]���)GI��j�g�K� �7�wI� n�'�����N��1n���Ⱥ�H�3�6�ȿb(�K������zu�ѝ7�2�	��~n��+���EZ��B-a��P�sd��Sĥ9>��o��,�`����Cjzփ4�'���i?�����ϕ���Ԇ���0hvUcY�үn�����a����s���^�|�	�?kKѤXً����7�=�J�o�y<�L�6�Є����*�T�nrK�fJ����T[����r���{�dz�������,p��i������e�M���)al���BP���x]��N|z�����g�r/��?V�a�>Z��7[@�ߎ�/j�$׍F'^ �Ҿ"�_��*����z���@�o���8�ui��	ؗ^�,'�v�).��Ve�@.�-eE�ؘr���GS�3>��$�Y���T�S4 \�p���A�%�_�5��A�%�k��HGk�a��E�;���,Hy[ea�w�9a ���H��,Jn�0<�R�_2=h1K�l"��̇�P�b`>=7V9���[Ծ/c��h���ǎ�r�d��T��.�/�&h(8���)~w�&�H]<��n�0[t��{GI�����ş�w�V!`GI�A��Юr����#�V3��G5�;���P1՞�Nў#���[K`�K����1�Qo���7���&3ܒ��6C��ЈR�Ǝ}�Vv���o�iYF]^s�1�,���}�� ��bXV��T��5c�h��;�'{�A��y�E���K���(�W�n? �`�a����a, T���)i'TN��"�)))W�P�����sr��wҴ<B����,N�^��Z��hag.,At��Ӈ+���0�D�ضP+�7p;���%P0��J�d�*�ui�q�UT5$;�;U�i/�1�Q�<�li�R����>̛���ZZD����(}�~P�#����U� |V�(�9~��c�	��;��6�:��L��\��QJ2c������K�P5�Ǒ�k�ޥnx��H�8��Je�S]�MqUkBx�>˸�/�+����.)�5��x��n�F
��k����< ���Ƞ�{�)H��1��lO�����N%Æ<��]�������oAg`���G�g^B���	�@����ei�%�� �~3Q��V����B����_h���:d��m��x��Q#�M.M�/�}Q{�,�bJ�ٓx�m��> K]�����x/@rPw{C��[�o�<��=	h����<�2�:�~�˗��d��UX�4�Lz�Hl?���IG ����lw�-ŵ�|��)��U���-5������͋�E�0w���/�pЇgM�c�K�Q~�e
�((�c�D:s���!w��C�tm��h�.F'���d�d���O�����NǀF�6X0.�J�q��-c0���u=�[�Qt�ʭ@j_G�aF���a��U�p����|��#���������^R�f�`���2��yQ7h�vM�!�YiO���/�1=1uL�6�^������J0��j��x��hУ���I�
�[%�7���� �koq�ky���bYF�UVqC�uH\�$��0>H�������~�o��(��9Դ@��q��6>�5�?�������f��Yd ֍q�ԍi�8^$��u�Ȋ]�B؛ü�����p�O��@ x�I��\��{�<ǖ�$F�XI�������.�̗�jU��ׂ͈̓X��P4�9$G�����b��\���������	���:>�h�����9��&��v�t�y+��lw���r�U���W�7���q�P���>�'���D�d#���@�>���'�� +�u�R��*�L�-���s�n��+�c|�=	�' G�Z9.!��̟��{�_������_�k�m�H�
�t4�w �����e����o��$5=w1OŻ^̖� c�x�,�u�.-�����_JhB�������y����,����N�ޗ���t�b� mq���Z�:|E�S��g����>����C��j�A��ڷ�D@(κ�-1Ws!��ƣڐ%r��̼��kR��r?,w��De�<�Vf)y��]��Y��%�8
�TT5�zG��A7΂�:	��d����u��W\.!P�V����&둭��<���`٫r����������@j�!��d�>��+�]F�E���>�nE#褩gM}�0^V	Cz��D)��D���f5��N�X(�!y��� ���W�ցR�ɴȝ�"�(xD(�CG<K��:����$�a��ǿ�/����K-���U�������yBg�gU�P��Q<�0�a�������U��
��,1Ջ��"�V���ڂ��\K������t�Nt��`~���ML0&�#��������L<^��X_�6M�����=��˳�?PQ���GjT��Qh8�L�ߒl��!e�u}��~�<!�1�����H(��K�̝aM����v��ȇ�K�K�8���I*���m��7x�ee�;^��_ɞ`�W$o5g�R���T ^C/�c��3�70�c���{����ty�v�j�֋�{����d�˺�V:0PV:�!�2��H�xfmi-lI�۬�e�� h��qq�Fg3����e�=���p렪�vR=2y�"������d߶��QR�����G۽3��e{Y���.�0F���s��������o���(����A�x�Zd��� 11�e �۟�}��{��{m���2�}D��������\21�R���m��8V�xܫ�8y�߆֭���ǋ�Wv���� �[�!��V���rn��D��#����@�	��q�EiĈۣ�yJ�DJJz�c���1�(�P&�׽����~��k��j�񫃥SD<ڑ)V�j%^�s�:�`>��;E�s�WL�3�����<'�W�#������I�6�r�L ����F����EI9r,��$8���Ҫ�D�K5�s�z��C$6qq��L�������qԥ������]���x����򥚇fL�,�8�}���<cw�����Y�m6�d��xJ9���:��k6�.���~_��ZC�mKP���B\j�W���1������M��,a��]T�`����˕��9��6��g�uԧ�n$k�uX�ָ|=��Op��(�����C֒�T��=�QZ�u;i!�R'�,�u.��g.��˯������Z��l�@���jgb!)��}6$��or�v���Ƞ~p$�5�o�a����X�d��'Q��8���,�o�<r� ������f���}�w&�@�ƍ͟�K�ɢ��~�0��A���.;�Q����N�P����Ǵ�&��҆,�/��S��uݑx�;a�D5��!�ď�V9}'��v��$8�"��%�}�P7�Z��!������u�%.˴��Ӷ5��������c:+d������Nhqm�Y[%J��X�Ố������=^�|:¤���^7�bo	��~g}�f�Ij���*�=Y�W`�͎�����3�?Pa�����(^�����c�(�{�|�M>��zuܳXi̽6�f5�����a�6h�*�+I�K�f~��@���U�d�e������9\hF�� ��o���O�+����Թ��y��CBxE�����a#/���^��IZbL�5��@$<�y6��Q�i(�ۄ
7�p�q9?ݜ���J�����Rɭ����o�- �'q�UIdXA=F<�	:���b_����O`���gjfuڞ��ZALB�������1����r2����u�6�ٕ�\f��R���T6��Rw�]Mq7��0�lI��Up/��&"=�)$�VY�fϫ�=�,�m��ے�a�47�M�M�'�6_�˾Į�z��s��;d6AC�,���1P���l��v$,�'ekJM��X����������{��� ���Mk�Ҫ��Py���@��׶��΁&|���,MRD�ֳ��~���	��9�Ս|�}[�dBB}M@�w6�g `�?���w��d5��R!u�6k�޴	��{�Lsַ���3����>�1��k�5rAJ�?�rf�R,0����MQi�s20����&j{N�����JQ�����Ĝ��@b��2��F$`y�f�/]�7��N����֣8��]��@�	� s�mgQ��j?@�W(C),=�;Z�UՁѩ|��` ��<5U%B(��T4Yڬ�cE��i��bL��Krę�m�0F����˱��
�!��	h�'��P��y�[��$�	#g[r��&��{�%�!!I{��*u��\cHʦZ��Y���O�fvz�-�g^������ ��k�R���W^`x����xB���(��4��ݖ��Zt���<��0m��jf�p@����~#XI�H�O�������uy�I+'n������8kX�Ik��VS����%v�6����"�L#�g�k^܉�!l�"�gG���u��� �9kN�|Hܢ�P��S���Z@�f�C$��WM��6��g�`�mjd��aly>�W�}���)�l ����a�Va�9:4�tfl�]�?:�_nA��PkԿת&�^�;$�&b{�Í���Cna�zz4̀�wV�!��?��^+{�4!�5	���FO3�	p�q5o#�r�q�<c��M��q�@40��0H�����B�'o�� 5�(��{��I���[�D)˞-BN$�u��;�N{�������2lFގ�&S�?���3���������-����p��kg�S���;��st�cqOX
�m�4۽r��`zUl�6P"1DSW��ǋZ
��̮��2�O��|��b��L��@lf
b�aI}Ͱ�=q��?�v�f��s	�%�n�dy����˲x2c���gZ 4�._�7Fй�b�����?GDb�����t2z<4��'����g�h�i�ZM���v6�pR�U�	$� ��AA>6a����ٞ���x�PhW@�!
� P{~�@�3�'N�a��H��kǻ)�'����V�Av�*�mfCE	!��:��|a*����M�{�鋐%y4����o��
3LZ��W̎
�o��7�`�̸d����`rE�M�lU�I��}�\ऍ��N��VN�j��@�1��V }@�޼��Q�7|1�'�!��L&���Y� \�Y�X�f��ٮ�1��p2�����M}C��Cd?"�GT�����_1����ك���c �9Hs¤x�&�S/&��X?�[�=� �u��������$@�ȥ|F5�;��c#�E�Sʓ��������Zl7毶�驾Ⅻ��pr���:�(e�맅D�3�
��M�WE$���_=��;z0P���1�P�uY�0?�ċAB��7˄Q��`�9xd�1��h��dB�{V���~95v��5�dl���4��Gw�r	F�;�!�I����Q�%k/��,���g�NwS��vÈP��6²�r�Xh�#a�Š����0wY�7�D��"wA����Wr����N~w3*����;du�ْ����L�L����s�/df�A�}�
�o���k����q��aS��gd���'ӛ�?o2��P�P8Y]+���E ���C�'p���$5+�Adz����DC��>�w�'�?�?�:��	D�W��4R	�R�(�o�b3>��rp�mΕ~��� ���|g����*�bz�����,��wNPw��i1g�������FI�	=�t�4���zUBkJň�������9f����U�+�;鐯��������!X�!��nF)�+6_��0�{L�R������AS?��1��c���γB7@YF����F���f�N��Le�}�C����"�k�9N(��e��ym���Xh.���87���+���!>lm�[�@q,b�����TK7�X走�\����*⭡Ё����$��	Ŝ~x��`�O(KE6.g��!�*6����3��3��oC���;$[ive{�I���$#�¶�g�(2���N"�e�MfL`<���^��4��A4=}��S[]�}��p)8�bu�xi��ls�,7���]���3՘1�J���Y��E�;@	��D@�Ƕ����#�gT��<b��V���AS'�eZ~~`�3}X�9M�(��X��FC�\��p��q$�`y�?J�6��y8���72@��aε�A$)�r�d����ˋӞ�p�/�WU*(
���,�x�X+�E��'�,rlBD����(=HK�
�<PN�y���$���%�>y�޶��U2���30a�����Af��%�o�VWLfA�|�X�p=�A:	�=��(��n�!78�'p�R�QG���ǥ{�h��K���<)�'�(N�q�|)�`B�S���M �����_�l�V�˹q=\ll���s&]ԪPl���9�$�=�!i%�v�`jU��ٍuB��� ư1)i�?�c���sj��h<27�S'�@W�ߗ�KŢ�M��h��J�4�[k6��Kq��	vG$ı7Cq\N�%���3is�u��$�YR�wn��j�G:Gq��?�'�!p�z&��b��a"\$c���s ��hM����n�L6	D��$r{�#��y-�P�4��Y0�SZ ��T�.�t`l��Zl?��ظ�bF�L]i԰u�aJ�2˒U�DJr7��̞�\A����~��h���C�5J�l/I�D������L��B9�\���)b�A�s��4��}PiU���)��E�ZD���vPMÚ�3�4cw�5��ք%��4��,��9�M�rǠ�ə�qc��6��7`0��3OP��0/�=2^���$B���.��߃�ww�ƛl����5�j!�<��1�@r0X��f�P�@TrGB�)�4:w�RO�`�K�q��ޢ��.���Q�Zq�[��n�$�sNr��%���bx�o�7�@1q��R�Y~�6����֥F;����Jic�)0���3�
(�x�>ѣ�T<m:e���- ��� !��U�t����1D�:%����l�B�Y-Dd�|�?�+���!Ҋ�&�
#���m�V?a�'�J��M����.;��R����n�k�Px�PN��L��y̿M	��H!ȿf@E��~�n���`#=Ǘ*�Rѥ
A,;ވ�&�O�}�C����R��I����ք	�r�����<y��+t�&�����+����p,o�Z�~�����_j�~�y�k���I�Ж��f^��(o��Mp�Ƶ���׆����*$�#�K��9��0%��'�ߊ�q��K`[m���M�m��D�ҙ�<P/)tO[��s����eEMt�*V��f��/<9ےz3Ҽd�ͦ�Řk?w([w�J-jZ>�v���#�"������K`��n�Ч��J������x����sP���y:�kr`:�ҊHI��n .�D8���GJmL�{��@�\{p������4����%���I�%�I�Q�v��jʨN�;?�3�$��q1�S���������~�,���nGw��Y���Y�p	:����ƙ�+�jS�����wf�,�J���Q �	�R��`p��)J���!��\�0?� ��!े��_�9�.�.)h�D����;w��B��DT�r��&yy+K�f&�������%����4�ڜJ�T�,Tr���:����t�tbv�1�ܴ�ނp����\�)^����Je��p�qO�]��U��ӓ���/�~j��"8W��#����B>H�AAe���)��5�b��N��\�K�]*����Q����k�G��<y�W\�wL����[;�Жb���6��8�iBZ�Bּ��5(yx�A��2����M�.P����n�H��E�~��ϵ�ޤ��.x��5
հ�K5��G���K��MfY?��u��y�6e T���r!�d$�u�|d�c�C�"�g_#	�ﭑ�Ա���	O���v"i��7`���p!��������L���<�?��i��_4�wEHk5�}3����|t���J�-����/ˊ�?�g�x�L�ςv�C}@�d�G9ܮ�{G��ł��v�dCT���\~�P�0�IqN	e������+�_�2�u.���;�@�Ӵ�@i��B�=�4���V[>0��0��v���Z�2��/Ε�P����?d�ٚ]�,*�,��*5��U�(�z(��;Y
� iE[me�z�f��ww*��U�2�Q��Ȩ�"��Q��!A���Dy�o�:����J�!��Zx	�2�+�̶f��B[z\"I�E�6�)M^�2���ஂ7�=���>�]ӔU��,ry�w�m4|m+�6���%`A�ל��hq5Y�㢥�g���ZJ}�V,J,�~뭫��Pmh5��'d�7�*�[�ʣ� ���pl���f���M��K��r����F�{<����f��D�R���R�W{#"�6�w���n�%7ת�/��M6��5ǥA��mф����b9�N4۶#���m2y,V�P0B}�^S���-����ωљq�uw\���t��(0KZ�zw�&.w����?�].�칗p��Ѡ#b�W�����dN�l6e����1�l��;g���(�	xj��������ˤ�� 2"�[��I��މ��W�ftD^Mz)�B̡�Z,����7\��?��^DY�:q$̔#O7�=�� J�U�St&��I�g�������x:���j��g�
�FF�(�~}�3�m���n������}K��Z� /�@�gZP�E��<�j~RE��&�2E����l����J�6�_�`�v������-Ӌm�غ�85�+Q.*��V �Z��)u��r-�F�&��ĚJ��I�H])�I�۠�A�K���W��'2��*����� �
.��*�ǜ�@������Ve)AB��7�i�*��lm�syf�q#�G-��k<��"���_��~c�i��ѫT��HK�|�M@��R2��1���?Z�/��8s�9��rHqn����Z�)]�7���aQ됩cS���ggƲe�5�T����~��B�q�b����J���t'3�E.Z��F��TQ ���h���&�qi����6%�ƴ�.sNq</�c=#��Y��Du7�����r@v�=)�FRlB�f��1{5�s�ꢜ�u�B�'��2�z�)G�Ub�o��q)8�Y&g�̥�����hi��I������j�hl��0�O�pB��l|�<\
>�T��i�Q��^JS^�u�	��3�A*�����W��O��9�;���/`�߻�e��硽ƻ���g�te�9Wh�Ԩ��'h��� ��(ztF��E��y�f������_w�mz����r�?�~_��~�L�'�ps��Ъ�U��8��A��u���G"!�p��LnEؼ�&G gNsք	'ͫ�8��)(�T�9(�+d�Z�"��+>�������0'��#���_U<7E窹z�M[4
�x���=���� `�bj��i9�E;7 Hg<@��Ե�tJ�w��I������E��X��B�b2\hG*��E���n15vUD@��,ݕ�{��.8���Z���gI~�.���'L>��n4s6�P�=��C���zY �X�E��[�h���/��
��N+��pR�ww��t��7��KgK�G���R�@'���d�Wy�ނ_�ߥV>š�H$��ٱ�.L����`�T������h�5a�mn���%: a���Fl�a�˥;EC�Q89K�����V��r=��`MT4</j�o�+�!,�~ڔ�����C�;���)Y��EĈ�"����"*��`�mr@稵�*��ý3��<��L�51W:�~�=�Ƚ�!e��OiYH���tu�;�<��fAt"s-��B���U6J F��������RN�/�Pǟ��-�_[A�۲���G6݉%���!K�JԔ���X��lL���^A��}:g�q�H�*��е{/<h�02�}�G�w�V�x߬\
�ش�PavŤF�Y�5%�P+���u�sl�D��?���&G9C��!����c2:2�%�jh�v@S�<�nc5�)�	C2vY��9���Jkk��kY� T���r�I�S��q�m��X��pڡM�4�W
�#�)�������-\I�J���ڃ�.�=��x3C��3���PF2r�,Q˹�.�j�m�-�?��N���\�d�ekN�����a��(�d<���G�%�r*V��	k�1�_)�n�w������n _�T�o,�^[@<�!��Q��SwL^&C�k_�mC��7���0�4�[�2��|�D�:܄��1�d���t��Yp2��WkBS��Ӎɢ'#2�VZD�w�t8�k����p UW���I�Q���&Z�C���<X+y�Z	��`馝7��I��(�ҵ�Մ��G�U�r�%\�K��zev鈸����K�qUN��~�P>6���~�?ޢh|�5���H�u�����4)6��-�K�.b�_!��%�^�qf��3�1Xom9^0>4\�X4= ʎa@+gպ#�Q��7�g�	=v����3p���n��+� �I��s� 8��j|YHPUn�1�)���<m�-4�d��pw4�[�Y�ES���ڋr�&W]r����k
�ЄW�.�5#��h4jꦌy��P���)��AԐ��
|��2��Ǝ|�wr����q��9/�BTJJQ�	�[u�z��V���ϸEaN�N�=����+VBC'8!�RO͞ҹ�^;�R�fa<�+�
�Cj�PΞ3�=j|c[����'�������K�{���ז������b��¡ԫ���I�g��>�w��֖C�u5������d�*c}x��Wqa�����L�����v<�R�@��g��y�^��4@�7|).����1��I@���Y���IF�*�M/�Ho��@,s��%��i����YK
���q��^D5L�T�hО���4z�瀌A8wF��І�� /�^0F����v8�P�������`9n^�!�
	}2���{��N�#v?>.�f������-b�?�����K�L�3"HǬ��şR1TRh�'�j���]m��dノ �Odt�9�˳�1&�o��o}���1u�����4q�a=�/�j}�Q��iW���1�y�9Q���f�3�G��� й�n��>�to d2�ɂ�¢S�O~���߾	:�c2����hQG�j4�~˿�Q������Ó�����e��+d��&%]_T���E<�)6�Y}���bp��_w��!�/�c���Z�XJ?.S�;|SVw��B���Ot������i��򞝨<��.��\>d�h�IYT��%^OO�ݐ��ɪ�6̟�y���[v�&�F$�D`��.�y��V�&?ー7�;��R���*������z}�<ٜA��-TpJ_�H���iϲSm�-�h�M"��"{�3vҿ�Ð�n�w� 2����Q�~̓��7	�@D]0�S�$�!/a:�c�Y�%�5^7 �Aٕ
�u��0c9 ��Jo���1��{��B�O�U
��ָw��w�LYG�-���YD�mX��$PJ@��`l}��lFv,����e�c�;���~}x�^�Ñ�eL�
�0����@��M�%�a��K��,,"4��x�� \�7�mc�A�����;k����~\����۞�t�Ǒd�G HV�Fif��KF:��H��fb���#���#�O^B����U]��f���sYcl�bKn�vN�F_��bF�L,��3r��nM���� 3��d����[��ﻥ�>�ͣl�ט���w3���D6�/���I���d��D�/pyW�V6C2
+m��_�6<F[-!� �M�uG�%t
�j�ͭ�V�P�y�L>[@f�1��J��D1�e]_�^�	�,�`�d��Yi3,�H6�B骬���}a�U�<KTr�:�괂�)'�1��H����c| )������P�d�5.C�IC��A� 32�2ȩ3��@NoOV�ZJ�����V]�,����{Tf+2����Zs��.�~|����Ƥz�v��ɠԊ�+)��=\��,��~�����T�S�Wq�L�(d��:u��%Zaz���YDBƹ��ф+�?A1��P����z��P�'��.l%����>���Ж�I����%l;?�MNl��m[)���Z�ub�7_���$��(�iT0��m��X��L>$�ٴ ��Z�$�i+��;�eD�W���{��
��P�J�uWxoF��d쏅�Ȝ�E������+�8�w.!jW�/d #ƛ�2��)�#m�.��U��8��#����]:b��1b��tC�ˉ2�i���a%&-HE�kh�-��8�W�ɷt�j�(f0��Zo]i��_������#2k�I�9�Y���zgWs����T��`�;x#U�Y�.��o�F:e'A��?�:�A����	Z����A~a�5! �Gq7��(w���am1��r�*h�t�q����M�|�Ew%������ͯ��J4���h|d���*+&g�1t�9ߢO#�2��w�_�#]��`v@��V �[nK���81���OD/5����Q��)0�?\�>��*�aw���'}8c+ܞO��M�`�}~O���y��o亿�,�E� �4؅������J穥�!�V>_�����G����jL����:��fK��ԢCNB�"�=�c��h{@{�m�cb��f6���m��k�f�i�UD��%\ċ����1�G�#V�D/��Y������ZMM�v����?�e��j���xf��E����Ȇ�O~�)����KmH�S߲eM�Q�Se���w���"�ak�}>~7K:��Bc"Hj���&j�E�%��O	שׁ,�7|��eu^���'�Եށ�������|y�=���y���sG<����{���G�m�x;��_%ټ���2�m;.�c���7��4��{��Jj�������W�D:��@��[n��3,�f�B8a\�����p�?n��Rz�s��']��y�(�:�� ��l��E�� ���Y��K�h�;@X�<�����4Ӧ���b� aR�G�G�&��%$}�q��w�&�3ֿ0\'h�2��Js�����I^�7��ۓc�7�G��[�/"5��s�%��ܡNer��6b��QS�-�$������^$6F>r�zB����ZY4����,n���"V��"&�zw�����������a8����j�������xo"�t� ������ZGl��f��H�s��To�W����FЕa�g���f0 �Ό��$c�0�?�iv��-���̨i��դ�&v�M�<�LGN^��=Y�>� ��Rf�T��H4�-�ޤ�����`h����E�Y�$p���8�܈)6p�m�]C.����������$Em!��p#p��UXv�g�_�y�n�}B�ŗ~�Rl/ja���s3j�0<�aN�̎V_���CѢ0֦���p|W���#v $������ӂGTp���F�6�u�<�Xo�n�;|qT_���cDi�4���R�,}��g�~�b̲�>�B��8Y�x�;�.�y����Yh�����ɤ��`)�-�-i�_hj�0o���#����?���'=��v��x2�İ\;���?l4բ�$�9)m&9����|v:�1�K��p+)��w=�o�M�k�_C��w����9O'L��;���p ��S���	���iU����[�"���؁Ht|C����I"�#+�����K��p�TQ`:ߎ���|�_[�H��>��>v}�����$i�p��ڃ$�p����d���<�O�ECP�`SsU�D��?�`W�x�����*!��Η�ڴ���"/p�$]�u������jd�³�q�[��;���S�R��
*0��������Pq�����7�c\V��¸��%�G(,����7�\V�g�F�}����V$�<Sd�.�عڊ�]�K���D|&~��rxk�DG�O�)Z|͐%Q>��-%$n:i�j���	C*��hS�C�����#45���F���Ş�3��G�ܑ�0�i���`�����Ո�>T��K_͡�]�:8A���+���q����c�C��(`�����g@�U���O�k~����˲�
3=�;��lF�ү搟��3?a'/Ӭ���l{���l��i����e��#���L��p����}~�W��$����5�T���v}7�YF!-ʋ^�6>�K�C�e���XvkP�䒬�NpL���ӽӔ{<�Tl��>�wL��9AsJa�!6;��'1:��]��9ʡ�^�	���iC?!rX*$k�Q5?��?6uR��i+�U�O.�H��|y�y�֔� ;X�����7T���9�`��~_�@ Q�ϋ�Iy�`ez��yޚu�~�e��e�<,�l�l ��Ve��	�����p����������>[m����7�2f�g���C$c%"�,�!�;�NH֪���l���	Q�7��C�)	�~��;��.O������#(�%6o/��I��v��6���!�� ��9��� o8��Y��s]�Y�3���0DL��p����4\�w*!)��򠢟�gQv�@pO�8����w����P����[m6#���?�J<�u�"7��s8U 9w�ܪ��%��r&@�Oz>�{��o���n�8ߦ��,3��1��i�]�g&?�� '�����J�1�Qn�(+�E�M<dHaxN�����.��p)�H5�'�� �jB�?ĕ�2ֺԭ������Z�fܝnS)*}|����6��YWv�5�9�&_�.o;������ܲ���R�� J,������1�av�?r�xt?��
P�Nb��w��H��
����3��ӟ2���R1�"�7�*j��v�3���Õ/�G��Z��ԷRI������0J��+�Ӱ��7!��H3���e�V云ey���������P��8}�Ў�X�3��.�������X\υ���3ਵ94f���9�h�ߋU>L��m	x۫�&�ȝC���E%��4�(�9�;�HӶ�O('!ld�~�l*���;���.x��8�VJ��l^�|����t�9� �Z倸GU�?a��b���Z��#B]��y�k���=�_;��x��mw���GD��0��ވ��v5O `ؤ�םշQ"�{Ub�r�Y1���U7w�ƹDsc��ʕ�~���( � �~��$�cX����IW��>/ǜLg���˚CjRQ�C��O=m�nI�f(\"K!ˉ���_�C	�S6��2l�5�����0:j�_]�ܮ�W*i�{�����0w�(��߿���z�/0x�i4߲�����ψ����:-4Gq�C�'����^s�G ��a�Jqm�ѳ�/NYJ p�G�s�3�u�Mb���ƚ�L���M'��..;�vTl���?4�XE�ҩ����^��{��5lK+�W�>mo2,|v6F NF8��2�f�� +5���hE�6����7�8i��ϵ렓�Bz@O�Y�&��L�=��]9�4uv��qg��[���!�7�=ed��K��$vv���T���=@۸����\Ǭ�컽���<�38{&)NF��41���.�dC�K�!P�*�����mw�x���ز%2����-:֯]���P1!̍�c��%��%�mj����9�� ��`W~�ǴA�n	��*������U��eU�^ .	Z?P��� &\�&IB� t���V8ڔpB�
1�SKm��#�l����	�\��;*���鏕¡T)����O�L���t|�>���8���3��l������a子�K6o��XB�h��]�Ø"g�f�4�T언�}܇�5�%�m}30�d!H�ߥu��A���r�AS�yՒ}��a﫚l�M��Sa��`az�"�z����;qWg�3�Ei��7,�"@k�	�XK�GU�+qU�N��3ӛ2�{��S��񂝾ty줈b`�;��o�r��[�5�|�$�����-]��J���Q���w+lXb1�L��ikz/]��?�:��}�6~���;�т�g���P<:}�y�2V����>�Z'�h6ev���9���u��7��̾b>	l�4S�48�AbA1� �:�/��3�����L�q�`�;����ٽ9��f�����PK}�=I�mY �x4A��+#X�<u�G��k�L�x��G��(���f��&���%t�"�!KFϖ�d-
<�� �!����aa�7��wU����#�N�d0��6��Σ��A�!˻���o���v����'�	G��L&q�#�[��6X��]p�[쭆�	���6�Ʀ���6�ۋ��6j�u�Yc�0R���yI\�����p��&�����;����V�Z7����}�߉��l��g�<�v�`�ny���S� �Q��7��M���SҴ4�^�Pzq
H���)D�*L�L����fU6g�G�%l�ՒZǾ�H&ɲx?4�+ES:,H^����Ĭ���vɉJIQ�A��O�|�h׊��z���̓�R�i����sU��wm� �OKz�6���vz�79K�N<O+1;e��Q��|5-˯&�E dP첃������s�]�S?K��DB� [C���>j�A�����2M�&¦���>q�&�̒��8K�	"��CbתK�`H��0��î�Z���`�X����Ra����L�����P;k'٠��7������IsS�ð��8Y���Ǥ�Φ$X��.$�0�0O��w놐ܲ1A� kgl�K��@jq$FrF��CH�{4UWq�N������i�T�'� 	��ٔ!2w�F�M��C���Aׄ�ֽܻ�qm*��y>>��A`ek�`,*�ֲH��%�@'�Y�ұ�W���� 0-����4���R���=x��9`�,����M-��S[�a�'髻�T�׫=�.�]��������S�/n}	�����]:S�~̞I�!��]Zj{`����A0�W|D%���Dh�`�Y���T��9��BBt��)�D!c��Öny}2����ƽ/�*�h ��M:������!�\�n���ـGDȠ�m&�Ώt��Á�h�'#@���n\jgW�$��;�R0�5�a$6�':B�v)��y�%�i/�5`3w�����%��E�����q��?�X�q`#���ov�V1m"F[�4Sl� zB���e��� ?�h'f����'[�jq<Y���-{�!Eڽ��5��!.ۘJ�Z_�^u9A+�U�Ͱ�Ϙ#�;�8�[+�g����"Vk�OY��g�1���p��j�A����S�����m7.&����i]xeI������M0@��1b��+=0_��� H�͝^&���4W �D�;�VB�_ߴ�/L���x�
�)rNG W߰8
��<u��L܂5*`�2�?p�J�ƥ5~ү���� ��%Q�;$�ᣪL���V���,����x��4lX꙯� ޠ @������te|ͳ^�����H��i��Ĩq[/�u�Ta9"����pNL���"���b��
���CCؖ@���K�]�.��b�y�n"e�i�$��ؕ���O��'��(nz��d����R�1ls�5wYf��Ⱇ:�0���D>�@���2�GP�i��P?��7"��́��]~����2�c��v��;��@(2 ռ��D[�<c��`Q'A[�I�{��@�@u�I[Wzܯy������I!6~7ˣ��5֞r]�}'�vy�+π�*�C�˕�ʽ�q�^}�|�:>bU�۠w?�&��곰��-KFx�����B/7��ٜ�HkЏ謁�$�w��٘��-�Ul�'G_���T�h���U;a�ߐ����v��y��D�9W@ry�Hq	�5�~ ������"Z�`��d��G��٨p��~I'v�$��gu#4C-:_�9	� �3 SS��a]��qQ��[�h4p�}�Ssh8} qTXϮ�ƾ#(X�#6���zV�㏾)_���56��T4�ْD�@��M�׈	$$\� Ycw�r�=G�I��xTs覹
M	*�K�9��#����w&p%?{�"�뗔uz��H8��N�P�c@(�h�?f��\���{Κ�^Q;r��I	��;8[��q��o��"�)�Y���\N���D�qEgRx�K�	���H��2����.L��c�9?��Ѡ�˰��,���5��V3D)��4����ޙE\�taI	tvlkt��tGVvq�1��NbasG�&D��]�H�)Fۦ�I�D�1�K�TjM}�"�8)�	u�'���:�~����	ۛ�;T�5? r�Xrw�Y�R�f�Z)��k��Ww\��mL?�"��(:R�*��(2�Y$Y�Jʼ w�'�G�R�� ��`}O�ap�V�։���ѐ|�V?�z��OT`A�GJ����V%t�wꝗ�+J��BgW�f}Ew�n 7�A��~)V�s���5fA��?��8��8LZ��v�U�kϦq}<	���u8�F~���Ua����Q4�j-���
���X�":� b��k�E^�c� �J�=�_2I	�H��VUvYg6%Xr1
�;�`�0������3Ğ*A� OK|6��S�n��\"���r�Җo/��W#U��R@(�[T�.�3D��%�js����#�t�ZZ�̫�5_��w4g�~����G �@(z7��r�y��ɓ"seؿA��6�,E�˥'�`x��2q��`y=�*B�)��H&"[g��m*5��v��Ӯ!���W(�"���g_��}���\:�G��]�K��zQ��2�vɌj�V�e�f�X���	A���z;��ں��i�ICP&�x�3�������\�0��(�[��9�/D]8F_�|����k#!pȊ�J[�ަ5&&;/��q�i��%������a��\�Y1_��)�I@S�3�\��%�c��~:�=���!Ɓ؎�Rv���M�7�/�ýdn"o@|�u�2樂�)�L�L�{d�s����'�3s��,��Pu W<-�/#:�=�nG���Ӹ����D����9O&���h&4w�Ӕ ��F����}f�:�V
Mκ袨��-�� �!EW���D�u85�^7���*w>�B��.�)u�-y�H�����%4y��^_)�F�H�T����$���@�{� iv,	`>�"N�	�5y�\� )'�q�&��μ��{Qٿ���DϒE�~�r�6�=Dyi#��d���v�&���c��{�����'J�9AbR�Â�B�\��V����W�U8��zZ��5-c��A �j���,ެǵu
'CR���-�,���hR81��~^-�1v�>���;)��TXTu�R�0�/ȃɚp��z���|��T����'�;)XC���k�ێ[� �u����b�w-�Gm�O�|SO�ru���±@�Ɨ|� �;7�Uޫ���Ϫ��<L{U0�Š�A�~O~��c��$!�7�3+sc?^Z�8R��F>��� ��H���47�?�S��e�b&�F�X���j��x�D� �z�@L��pxYg^�p��-e�p�.%���C��`� x�[�=c�Rfe#6�Pkl]�6!�[X�pf�\���(�����G�4�|�Ns#��1�ħ�nn�D����=*��o"2�i�t��˂qh0~0Jy�9�IQ���S"Y� ��D�r��b��NQ�Q#�MD9{�<�� ڇ����<| �[$�>�Wl  �A/��U
�x%�7�H�
ow�%n�^I��_�cL76pR��F.��s����}��燩����G�&��dY*����kN�[����=������ׅ-��%�;��T!���G1����X�_R~l)�{^58E�j7���T��Kp���#Fz��R������f��˙7 ����w
�=W�}�[<Z��� 3i�ѥ�S)����Icfb���X쪏��蘒^�M�6��YZEs���,�����gGm�:Exh宧�	�a��`kR��5Δ*�Ǔ�Xd @*�[_XP[�`N=σz.��A�B]�*������}��F��x���Ќ�����}RO}Cz�c'����~�F�'ꓻ��ѳ�`�F�6iH�C�Td_�A�<�I�cgn�yK(Hs�(BQ(����֎��-+93���&f'���M����IGg��Dh��a�o����I;�5zV�dVS��
]Vz�V>�^��Y_�wKW�%;�)�̴���o��`�ܹ�>э�eWA���@J3,t}��SWx���~�s��C�چ�*��-6r$��E���c}Q���фUb_��vr�j���i�M��
*�"�a�{�x��ԇUJ�@hDɆ|����d���"�ޣ�\���FǐQ���y
U�>��k�(W�l/��ivԳ5�ܢ阚���2�L���A��I���~q��m�2�Zw(@)nI�PL��UO�c��q����.T���j�Wx�z.\��W�J�y��h��>�պؔ��RY������G�6�G�lo�b`��a�!f���H[�{�3z����]	�+a˭6�tD`Z��&(��i���չ���Ld)��?�7�v)x^%ͥ�5�ɦ*���C?ʕT�T21b��s4�H�Sliz`�>�(��e��{,��Ơ�M ����DָOi	�pq�i�6X�{�8��`0Ws�)u�a$�~���a$Nd l[+�<^�izt]mt!J�OF�eI&�&?�"�4�e��<�G��gL�as�|��&��g�q�~�#D�V�ڛ_��R���=��RxK�i�����e�)���ú�{��,E�'�2S�-���!)�-6zu�a�oWI'&��ir�Kjs��5��Z����:����
�6-����i��������a%TT/x��u�6+�P[���<9�ϴ���\�!��SKi�s�������sF�p��h�|�h0 �#R�����,�.�L���c��F;HM��p�AB�>�p\bH֓�7ߕ��w�K��%�iE�@u��1�N� ��͒�8��g�(^9��ެo�t�O���H!�傂鍘�m!k��}��.�s���E��V�����!��uә�q9;xbx�j�Do��׾'aVa�=�;q����M��೉����f���O��}rdr�=�^�8y �^8tP~�G���)LY�ƅ��h]&��#���K�yS�l ��3�tZcq��X��T8jJr5�p��kV;�x�;ύ��'�]&�����B_�yz���W	��U��6.)����b��V'�Ȅɑ���{f��e�l��vq�[+p\��n�;yaҊg�d(U,�u���2M�����%�u0��S������n����!��e"�ג�*%[?�T����UhɈv��hV)��})B���ÑH��Df5/� �����:'2���Q��N����7A��/�V�r2�Q��'[�Rj�G0�6���G$��V��1˃B$�2D��X3���Hu����C0`���eZ�:v�Ƈ��B��5Ğ�l!ڇm}�����޶W�M����_C���1�R[��V�&5j�˱��ͦx�"\��:���Rh�A_�";���	{ń.2�n����z�.p��We?2�S����x�L�CC*���aO�Nr@e�E7�]���im}�yk��m_��M|e�As����K�~������ 9�A:O�����O�լ�ĆΗr��/�SЊ5��jJ������x����U��g��dJ�>��B��gc,Ak�)���g%��'jPq	D&D�>7���Msi�Y0����P�x��r�@��� �B+�`���U��kL��I�7}�(KM�络9m�|H�C�p���� nR����B����~M�O��y3"��@����q ܎���،��Wq�p�)���Z��:�BO��mɦ-=q�P'�jZ�5�K6�����Od�HsF�j���J�* �K���wz����-"������N7�����۵���H�8P�t�Wv��Q�C)��_rBT�o��(k�6�G	�$�/^Zh�S��Ġ;F��O�Y8�e]L,�'��t�x���s޴n
��9��UN5����}N���HE�����Wo\�?�7�,_����7�QZ�"�xqs��5�R���?@��
���$ƨ����{`�,�Z�}	���@�Vy;�覶*�^��/�RBI]Vr�U�h}��]m�U6�5')�x�0BbR�6���D�g���^{y�S˶�
��Q�֦-$V���C �ɇ����(2f�"��ߞ�0<V��w��짐�xE0X����dP1�c����J����8�@�k�C(4��%�팦m�57az@:~7`��O���\�T�=ƺת�i��}����x�d��`>=p�p�a�������iKQ���YmفT��m���É��K��_].tzN�j��jz^��J��o�u�ރrA�\}&�Ў1ҺΞ��g�Z,0:ʢH�)����)�����k���3qJ�g�8�x���E��s��nP���-�x/o�����M>����u󢖆�3��z:�`��T��+ߘ���P)��d��E	`F��c��x��9j�������m�&^ߚ�]��UQ���9&��$��#.y�����E�yA�Z�;�[�m��Gُ��*�� ���:�p��7�56�l<r��`]���\.�G5�`���O�?K�*c� =��R%f����g���������,�Oe�-���\ Ύ�������k��d��7�p��lC|[�:��mM�j
KU��_��s���i�,�-��s#�{S!�Q���t>{)�v���-��|��c��c.�,� ��o�=�w��[�*�5:�6BPW(��F)T-�D��UT1P��q W
87f�p�LU��Tkn����9�lX���^� ?��������
���}!�v���'���g��X�3ec؛��NTw��ӫG'��sa�[`�m0�{��'t��	�f�J�������HÝ�0��E���#?�/P�˧��^�Cj5�e0��}~��g���L����*�[ ��t���޻� ��	J7ד����Ƈhe0I$'��瞧�D(b�£Z��G�h�]�Z�h���U�l�3~�O,�.�����ȝ��l��K�="�zMyƆ�򉰖�D�B�b�b�S|a�Dz� ��3$"��=��K]��"Be�Ⱥ�B�������7������O�U��������@���63��a{��gyS�.��K,�K,f @&M�,����5�)�[�����v����.�NA�c�7FLA���Z`�W���S���U�V�����1�7�#0�@0s�X~~���c�ͫ�IvW�� �IΩk�Ggnb��cnV<g}wza>�6��[e��&�j��Ĵ+����Ϋ���wŮ�~������G��^��]M����+��7:��+֖ӶE��e/#�7Uz����X}�A�5�
=⦾��I�a)r�}k�Z{޾�Ф�Z ~e����OX�ʐdk��f����M-7�I�Q�[Adn�S�ܢ��0��s�V����-��3�aj��V3�8�J�X�q}[h{_3�!p��I��"籵!��޻{4ᴠo����E���go���˞*��#^���p����/.�\�(e[�6� i|��D;�>���U_:KVi��^�,����)��}0�0�%V�O�f�>��Jo4�����vlq:K,�����L��[y�}L�]�C��t��;��_�~�M�y��Q�5��l͗��cJư�ꦃ�BFBs^<����� l��@�3�8��m�3R%X߱/���:q�l}kY>	���;S/Ao�X��96G!t��<�R�����϶Z-,�&���"�`�@��YNuvMYۆ=S��?\��G��)�6�08Y�E�Ԡew<�͖���	/E@[�����7$~��9�:�*U�#Ny��:4:$��vb�],4��3��S��b8��������9y?K�����g�GzL6%�n��'!�����)[C���V�6���|X/E*�NVZwl=n�a�c*��3�wJ�3�s��z�绡�q)�s�#`��C6��J+ol2��O�D��'�f���d8z]b�U���ʪc�C�$�s���!|��aH���.����F�
��형6Lu�A�_5q@��!+���Ve�7��Ԑ9�$%��wα餈�Cyޗ~Ws�`�]#tdS�7��u��X�����]k�aP^����	��&@�)�:��
�_W@ �a*�r��8�ќV��c\�̾ZK1*�ap\nO<zF�ɮ����I��������f����H̜@MU󌈋՚m�hI'���-=j�}�%+��"U�b��3Œ�y�ʅ+��A�N+����|C��ȑi��;9�zHu���FhS���O�)c�;α6_*䒯���
�$k��v��q����1��ou�N�2���b�Ob��$�t9�j���A^ͱxn�-�1�&��W�FZ)*Iͥ����R�ô^ ��W J̎=��#��*[�o�$�l��/!������+�t�������������=bA3��^��J�g�hǺ�Ȫ�`���y��`�?�4T
�bĨ>r"�,�M�����߸n���̥�����Yk@����fZ�=ɯ� �0�C 0���-z�k"2���Q�:n��y[���l2��&����ut��N��c��3Ϡc�.iogO$��5kt�0_�?n�@��I���'�G��� �c̲����@�͋�u"�u臛�z� %�-��d��ʰ�2�m��	$����X&5����n��?O�;'&C�yY�@]��$X��l�w���/%4|����9M�d�|R��Ruǭ�O�%2���ŭ�oN����X���*6<>|�@��ױ$�pk���d-��M�q�Օ~��l��4N��l��|�B̝��l�BjC㐹4q�ד���L3d(�$�}��d{$M��ڦ+砸��UM���X���mEfg�k����S�ZRr��.�IS���� ����c��I�����11w�?��
�p��
}V���i�=@��Upn�"�u{��V�u�%m�I�4�S�	e7�!�����*� 8srUx�-Q�$q�Z�$�"<p.0�K%�g.��q����� �J.^��\�6����Po(�O6�� l��������]Nر���C6�~�l�p=�SBj��Wv�?3Fq���FW`����@��~$��2>!�wE��QW��b�0Ⱦ(��|���k�S茜$�wR(�!�]������3�x	M���W@e���@m��j����g�Fj@�Av���J���.w�p~��B�F�#�Ҷ٫eL�w���P��3��-Yw�[Z9��=l,g�]n�2�ZA�(<h�1	�dw�@>�R�M������J,�қ�Yv��0;0���
��/����suqm5�é���4���S����-1���h#�:��*F�����XC��$Na��yVkk�QJW���j�xuU;�N���t4�)U��k� !���������f�j�Ep<tY̮���l�d�Y�bT���N�ϼ�Po�B#�}{�~���а �c�24�Ό���p�w�B�/�+�p�&���J���.1���pMw�md='ٟ���zE�����76�{�<_������(�ll�wt�8������I\.?����Gh�3��NVo܂��ݡ�]�>݁g��X�p��F:|K뤮������o��i+P�[�:";�FvP�R:.=57�fzd�X4H�u���X{,�Kq�fl�i���g����� d]
J�gZ�O��+:f᭠���_�rZF�lwżY^h��ȩ���ys����oh���u�� P![i� ���
�X����I=�6D��^Ղ��u��T�;���j�x��w6��̷��ach��P#<�M���o
`�ڒu���Y8��CĎy[^W��gxi���h�H䳾�@�����y��.��~G�	��];0���Ri" ���¡:ςH7�*1Wǀ�O
O'�f_�������w}!2�l9d%;߫X8,��_�'#oU�Ff@6��G�Y9�e��=A;*F��M��~G��d�~]��J`V$��n�:I�-a��}�D^�:�W�2��ڄ�G�IDoz��:��V�k ���LdG-��G�.�����-kQ=e}L
��-��%{&�K� ����Y����sL�,��\�&�&4��}���|��R:{�%��D�y����h�*a;�N�߂�q��%��:��'���z�P�7�*hs�{϶ɶ����`��pwf$3�U?�?9ɕa|�@������z�ą��f�m�q��TymnU�z϶'����I�]_�?K�V�x�i~�i��:�K7�W嗺	�|�K*.�ŧ�a'P3Um^�M���$w7J��)���)/�0�TBl`�ٛ�B�K2�s�I� �,G"w!^f��K�r��{�`%"Iy�mF��q�ad�ځ�8��:x�s��~��j���N0O��W��4�"dG�X���K#�F�����"�R3M�27k����_���eM��H���cpF��I��ngSyc�e�=��$z?��y���r�/ ��3~��W9�c�s�͓��<i��_�b��H&m�mx'H�e�K���Z��ਲ#���i���Dac��'Eo���0�{��DK���L��~�sT����?t
�k�@�@9�j+�ԣ�m�������"�cc��J�nۡ����2e@`�d�`f��������&�S;�_B�<�'��OM��kI��l�Ը;��}�@v!����j����9p`��]-;"T�����~R�t����u��g�Vb� [�4>p�HD�^����"�f܃M��j��S��R_�Ls���0M�����<��:x�h��"G�k�n"b�X��ҬQ�fy�ƥ]�� A�#���zT��W�H<]ߊ�q��g�ۛJP��iɘM�Ēd�� z�e<���d��Ϟ���JL@kWFp�����g�- �r�6��܌��TqS����T��QgcD�.P���5^��1�R�r]���ڑo��+>���GZX{���O���b�!�Z�*U��+�\�����p�Wб��t }ve����O"RXԨ�p�^ 7~�J�v��`6�If�I�B�s�ˉ�������a)��ǩ���<��5��a�.����BtBjrb�9<ҬZ��QE퇆�}�AiO��-��&o0)?��Kg��Qbl��]�VswL}J/����J�`���9cgb�����[só^{��S���1�k������3����,���h�V��m�ao�xx�ޥH!��wt�/�I|fC����h�����C�Q(��-�bd���P�)����iYŔv9޲�{��u=��"G,��Ij/�T���hjjtI`�3ƇKVEyڽ*?s����`�R�n�|��YAdAr
�v�� �����ѡd���R=�̍��Ϭ����Z�گ�W,�Gl�_]8'�|U�bT�����o�{}�g6�����t:�x��l�)��L�I�_4�lo��:1�WF�g1�#�*��4\��e�N���2���+{���+d���!��d�,�0��+�+D�j(��*M5A�.ڭ��t�=�(�L+���`d�Qg��׎h|)*�b�]�3=���!h�����$?����Y�`���ɥI+�f��Fk�q��Z�w�h���}N;i
�;�XN�1x���`E ���s"D�:��lp���:j�=���s�/����m��ߢ�4�F?��+�l��u�_�U�X_�a���Y8�N�ZHJ�߶_y��x6��?�v�:в�8��k�/�-���I�E�^�7��P޶����@�M#Ψ�>%�͒K=��F� @���=���Nӡk��7A��IyoV��U/��cT���U	i�$�1l��Pzn7����e�cM�1r3�\[�D�kSۣ�$�fZ/����Ц�K���*���ޣ��2�{�_o��"뵚V��6��:��U9�Ta����Ջ��O3�9ڗ�e��~���t���_�n���-a�z�'�EQ�JҠ���i �\yZ:�}�;����p�X�({5��~�HJ��0�ƈ��_�x�7E%1�����Z$���f�,:|~)��Ɣ��xnt�j�HU�q�����W�x�ޑR�Zo1�O�{��S˻��e�ʠ1��y�)�1)YV�$�\ƹw� (U��uǤ�*d�!3�򟱪���Tpm�2?�5�ژ�_:��������� ƾrb�)R�����2���(�6�O5B�1�L��b�|�g���(����E��aȚHv�#�dK휞���{b����sH��^�&C��rk�:��ە��c�_�� ����&����P=�Q7Xf���׺��n�W��JżZ��Q�rjy�\���R�J�?ըV˦?��UFh�D7T�6�<}.��*W�.Vm���D�9���N�@���/�9'�����~�4ԋk�0�6�»1@���L!X�IpV��L�$a,�tӣժQU�I�̛��ヅ�U��$�+�j��7��㒘����<|:���$�^��!���t��89��k�}?�J.���Ino���섦%�Q���j����� �2���r���|kf��o���\��-k܁C �Y�������P��&�����"G�5qmBi����b��}���rFv�����]Q��/WpU�`��ɓ�t}U�՗�{�.�z:����X��G���M-��?���3@I�`���Bw��������?�-G@���8�a�xz�#i~u̅��+�`V����|����w���m��z۬�E{[��"�E4p�I�Jc�h�궸��4��q� �0	4]�`�hJM���i.��4��Klf:E~�
@��:���b=��\���w�*�b�ȹ���L��V�5��Pp3'�P2G�;�_�g��p� �5�[ѧ���b����i5㉑1�B5�:L��F�G���My�j�q��x�i^sq8�{��S37)J����U�ye���YN9s���u�5��R��T�
;��&�5-IgC��7�5�Qǰ_M����-vi�$���-ac��M��@��r�WDN^&P��%�p����d�C7t�y����������(�����Ƨ1G�w	�"Ίh)4�������'�HO��C;�k�?+@��i�CtP+A֬�M�����B��'O�y���N�}ɕ��J�C�r���������}�v�+?=���j*-h[����m,�w.�J�1�y^�ۋ���GF��]���W����#r{*#�~kgÀ�su*av�/�L�\���e�v9�H
���0;�/DUL0Op8тj��-��$q��4�@�ӫ ֝������,�1�c�K�b\F�%�&��|�G}0��IN�A���g�h�{怊{����`F�b����V�+������_�ߟ���M���%g��ML{��n^(�E����L������8��9�QMg����������Z���lXP��9�z��R�q�{F黨�@�s�%%S{�DX,f�*.t+2yDODW��w��=�1���0��Q1�9Le��<]uW��A� �1T��-ix�{�VĦ.}��"��.��Gg��*4~/�qg�P�嫺P�b������D�`e<�{��B]����L�\�W�_`.I�=�:{����2F��<^	��5:U:M���<�`Q�8X���T�h����m$��C�m�V���-��e�yGjk��<iP�'^�XR�:�*ص�<PY�󙱲�L_;���%:�B`���k�{f�V6m�nM�����ܑ=C)U+����,H!J$|�z��2�-ޒ�]����Ɂ�����N� �2�Q0����,#V �V���!��B���V��n;M�(��_�+���7��CBՎ;L1�*���ڬun���˝�����l�%����gŤ*�^&�6XgjVb�uu�8/�Q��9��]����k�S��`�`a[��t�	ʨ���g�dp�(AW�d��[w��c�(�IB��+��EޫOc�8�vK�LG�Fѕ(� .�U�	�����
6��2F�P{�=��ټ^��(̩��8?��yܕ��ͳ���.I��1��&�.���i�f/�Ƣ;h�� �����k�"�8}�;R�H���Y:4�[����$�p?�L����q�/ne8k��v�`g%�ŏ�g�70�񕀧9���z?"�G�&u�^CV�� ���=�F�4L�C�ڒZ�e��8k��x��P$�p�ܜ۰7+s�ORѹ�h�b[�>{�^�i�7�]�ٍ� �Qvi�U%�� �� a�?��Hћ���I�LZ�T��N>��h�0�`���˙��_rl=E`Q�o���q��!l�i�j�u[W����~�)�hj��-�2��yz%p������0���@����PN������?$�)��o����OH
��}�
ĉ����YR�j�����k���^;��+L%Eԕ�D��՘n٬�{��h���rA�N�\S����lK@)2Nv&����t�ϻr ��g�u�M;O!%�pAT�J*瞝�2I���9��Ux�fH�ED4��y�b�=���w%��]=���&�������:2q��P�G�����`����ٹ�Rtlet���$����C��8 �a��Nj��2��.��3�IL\"DD3�i)�ȱ�g�#��:�.50�!t�$R��%QWglk�z��OQ���q,lS!U;!��@ɴ�LtR�� ��~1ƫ�{	B<��i�@�e�����i)���tӭ50����© ׷�wQ>�I�5l�x�_�קA?́��#�vI"��:6�2���'�Qo6�b{�� �`qUMox���,,u��b���0w~���(��m���n�d��h���a�i��ai�9�r~+JW�m�T�"���酵�6�p�os0����/9؍r��2�����:��ɞ��[�� �ev�!ܸi�Er|}��]�m������6���E{O�A�@���[ǇWPg�������b��Q�~t��0�$���[sT4m�]y��7郬w���˂C�@��=N��xF��4C����1I�w�	��lxE(��)#����3b���ļ�aOvso}�����]٢�[Sc�u���QH"Ah��2(��`[1�X�;�-��/��uq�w��հP�wx �Cs���)#L���G�Ϋ�Q��/�~ɼ�B�_G��8�_�qVhxn�pXw/�n.)��svK��͖SO�q��'���RD;��sW;��Pa�'�ō�ǥ�q���ZDV2ݵ���n9>ͯ$� `ھ�[ƴ����
�)���HT(� �}�82Oz_�J��b��֛ze��-p���)��V+"��Ë��VcA�O���+K5����7�62GDb~3�̞�C��Qh�$)�O=DE뫚���\�`���ҡ�ap��vA�g���k��I�^�Ű�ۤ��[� ����fH80 3������G��������ҵך�cb��\�3����m҈S���:2���7���I���\S��RV��И�5����?)��.&�Z�B�Ȝ�,u��]_�VXս	�������|z<nϤ�{�K�dei �9�*�I^�0V�z7�e�w�C̽���;O�[K.��N�v'���d���	��U32=-^��}4�:��"}ߚ�\�6���=%!��T.L�<�E{��ٛ�NjW\�$Ǳܞ��ۑ�O&�`�E؉J�Vi�[�m�����띩��^��\��*���xR�H7<�:���8�]�U|����cd�q��v�*���ws��n#�����!9����w$�50�ru�����ΥC�m2kC0��MH�c=n���n�֐�G+
�|��"X N*���J}�>3,��ǝ���^̻��e�84'�Δ��v5���㈗ɧ<p#f��T����!#�%�v��3D���?�����kW�Le�%�˿�)���X)�ǨDO�!CU�qF���,�R�eJ��0�E]%�t��
,>�w�[�F�M���~?7ְ�0p�qi[C��O���$79g���P��D/�k8��/Λ�J���T�h�١��2p�oN�$<�N�Zt������!��Ү�k�������=yN[;������Ew��M�4<��.��0�3B(���O]���_+�d5x7�uCէ�
 I�>�!%��ؼ8Gi�AL����Ry�|W��Q_���ԓ�ʷ����o&��o5�~�3+H3�+\Ѣ�I/�<|�C�׊��-���M��Y2NX<��$��
�C�ܾD��_���ȟ?yɚ�5����R��GO���zKg����OJ$v6�澈�W��!�a�l@�'�f�-�4��\�F��������/?�9Q����Qx�on���Q�7.���Pbt�ݝK�sR�w�0��3bRg�\.`Cޏ� ��<���t���&\�j�1���(OɃ����p:�kè|H�`�鲝���F��o
���a�)S��ᵉzҢ�H���]����p⥨4�d��˛$��@AY
MA�,LK��c���O)�GNߟx����+s0�/����W�X�F����Մ	�n�2]�p �C�A�-qC	�T6�O�C{��Q	��ǐ��IV�|Z>m2���dXd�:P��mP��=[�����6w�"l�y��"C�2�U���_��A1[��,����D#��b��~r���]s���A%���n�ڍ�Xk�%f���+���9�������cv�+�_Џ������G�6�6�����쨕��{��
����t�C���%C��rf��*6bC�F���I��n;4<�:�H4��O;�L� �@d�I�vhb�S4H��_�==�-;�_~�5'2������k�*;IS�kfI�C��;�#F��#�x�f��O7�aL䔍C"�E������}�H-T�h��;�W8��>SxÈ�9D;������ܽ7�y��8A.��s��/�L�
I�*��-�
	_���B�+�G�&�d����9�c�:�:��!��{yanVr����{��v�>�gX�M�L`����ql���"s��%X�.˻N��,��q8��!:��+I�ˊ�����h{���C;��J:}�V�i��d��P[+f� ��$G��"�l?�c��k���u�y]��8�U�����M���ag6�a�}Y��ڿM�p�Q��F�-��Cg�t�nU�d��*4��9��C̺{�pI�ׇ%!�'�t�˭P��Fs�ah�f�b_B�Q]�w�c+�".^$��\�\����M����&��+R�mgL�}����.�G�!�j����Vt+8����t�p����$kj~��/��A��2�idc-e�k�B*�Y���,�^K_0D�z��ra	�Z�.����D/<cw�Tm�T��]�)��6 ׮6�G�R�j�4$�q������g��ǉ"��p��O��f���cWG�W3U����3�>E0��{
z3vj��F\.T�z�e*!��9?~���J�}�jN2����*�2f��s8cvƄ����1i�b�d�c56{�/��)���o�����t�r�67�*�o�^���ƭ5U���qL^���u��H/���̬�|���C�N�r�(H<��\�$ΑB@� |W�;����.����?ϲ�}�ĤMR�+�Yp�k�(KrEۛ�%�a�����0=�}��D�����t��!���&%�g�-�g�^�X��=΁NJ���k�t3���-}ѯ�Qr��*z|���������&
8�[!�6:�W��0ڋ��VY.����lC�>��,�3�"�����Q�U�xY,nՎ�� {^Ɗ��?�Lo=�MMB���]���l>��$�aOH�b�f3<�;I�S�"���[N~��-oJ]���¬+�Jwa92�ݪ�$��A�����G<����)�JILY�E�ԭ���tXo Y@	H�K���c�$ ���L�8���!���o��h���͒�)�c���5�I��T?���� ��⿘�����#��u��H�a�(/�,T#�^ɽ�y���7��I"4/��]����ԇ3/���h9)�Ҁ�D�[f�oL�c�KA���]��i�L��`jR��.&ρW�v⣇WU��N�K��)�$�)���q���77���sy�[W*�3�S�JK�|��/����}�B.�t�a�ɓ<�<�s��G�KoS��
y�z���j=�������ן^��ZSA��`oA�˻��SΡ��d�̓�Ћ�dիA��Y#!J]S9T��`r��gs�VN�_	��:l�_*�uл�u�J�6 U{ev�6���P��$�K@cK�+^�`��̞�ګQ��u�:�)�}�L�`��Ǵ�Ǘ�G���J�ӌyVKF�����J�+uw�NXԟ���&�N��&�zl��_N�3�a�(�d�?^K���<�҉�1��R�C 66����;���l�,�"�W몐8:���w�6�s:ߓ�>��伤�������b�VvCo�bｓ 9lN9�M:�3���4i�A��yj����^we�d2����}u]S�;ٖs���F�P���h̼Ą~��sě���{c�b�Ɛ��l~.�ݡk��:�J��"�Ѱ@��8��<�-5[�ں�2ƾA�dn�b�_~h4��$a�f'�Ŷ���<d�8�&ӯ�li��O�u�Bpy��� s�S�R3Fo<V�)"���Gm�U찌?x�K�I��G�3L��4c�M���a@�<T�Q(#��5�����ԕ��^����9�&]��fB��C�Lś|�x�˚���Ha)f!�錘�/_���	{�m��4�:��1����[(��GƯN��/��	��Mu��R֙.Զ֢��kX���y�Z�� �j3ʺ �	�o����efZ3��2 ��c�ڕ���W��;'�S$Sb�� s���]Y�m]� nF�{��.63����R��$�{Oӿ�B�XyI��кB�mo����W�l?@3��o�=y�i�s�=��iZcp#���S��6"G��i'xZ��3��c�?G �SP���&j,9G���U������T���|PrB�,;2n%��:��0�q�m7��7�U�%s��b?{��ɉ]�p.	��u#�|��p�78���'C��1���p�9
I�S��9(�T���澈�(H��ȤG��'DX�A%~D� "�|������Q�H�X�����c�ܗ����U��poђq��l�N�7�ŕAM^���)��M[EE�����v����e綐<80�Fq��o�ʛ�:Z��o��i��no�̛k�6E��ԁE-��w�L�l�PAn���!�����o=�˻�m�a������{�6�T��>`�������(�X�`��TL�5L,(�~�˓|L=l��P63I��-1���K�p��]*-k��$i��
r��i����k����d���%��t�9��hf��
KdPop���}x�1�R��ɪh�d\���5W�L����gnDVw^����܆�+MG
�������5���fKD��`��b�x*�u9v&��-���g�6>;%� ����m.O�e4�xT���*oޱ�*(�����Lʌ潠e<���g�2����FN`C�}Q�0�2:����H@�E������h�Z�]�얐<�E�2�[	���5sv���Y��].��1��<�>;�&�7n�@�a'ڼ*F�/�16b��}�2��B�kTS����.�����s�IS�P�д���[�LO5���
v��fl:�5�^gz5��1 ���t�&P6���QVj�cx#��{�3���v���ě^�X��C}T�X���-I
�)�u`��K�>��52/iD�>w8�.Eͩ��ê����'����/6~�jV���\��q��H����txy����!�bQ�xa�:tV
'͓Z��weOY�y�^��]��FN�"L�m˦ڢ'/Z1s^�R��^H68?�d������R����5m���'�Е�������y�A�`�|����Q�Fi��{߻���w�X%\0	�8�vJ���Ȟ�_:�r��7�T� :����LK��k=�G��k���q��������� �D���#-�+1�_�M&c�\��"p�ت7��W��a6�#�PT�W0�C�p�>l�8T�l]��� �DC��2�|�FX��>O���Q���d/�>�&��'d *Ɛ[]Re���)0���m+ٚ/RB� l\�B���|��	 �j�es����jw|�_%o�ƶ�L��U״��=�D�$����Yv���+���"P��%�(��I�?������U�K�#�[W�[���D:��y��}W`���h�̤��%ƻ�^���DyWs}|�D������(s�MѸ �;N�`��:�DP�܀)�zx�(�4v���9T�pè�I�,�Rs�� >Ya'_
����1�`�Ų����m	k�c�gY8W�=�Ot)ݜK� ��C�v�6W(�4;�:\��I���`�Ҭ%��s��\���*���h�z��'�~U���
�͕"b���ﾳ�bc�CZb�>�Qq_�1x�� ��R��3w3���NE?�R45���h���}��m�EY�?7U��L]���M��S�;]���I�+N���[��][��+��bW|�v�}�<cyoo�(��tEO�\�3��9�9�3'*[��v���-T�t,�Gg������ �S�d���TEEż_��g�U�T�C���R����C͟Ԫ2c�-�|3;Џi�^7������(Qj�@\�Q4��kI"��ۭ�ޗ'O�� �Z�R�/�B�{�`��P�Ci����W�h���Gơ�@�P.GKm�����TՏ����mH�f�V3i*��� ��"��63��y:�gv�6=�z듭������3�M!��;�L,�,M08x,-���M��}�T�PY�:����;�HLuC�����u��b��`�̀���-�w���b"���&��gEY\�����u<��}�W�t.��:S���ty3�2���b���*gE��t�^�������F=K��*�'bWqOHhH��ҫ?i[Eէ�A`%�c��W�
�G��x`���'(]{�\`C��Z-cͬps$�PI��p��Q��u7��nOĻ��n���]�o���5���N\���{�,����-�`9%����;gd���}���"l�����)�g,w�~ջda�'O��
|@��
�P�b���K�s��t�����K��+�p	�˸\������w�ʍ���x���H򟩥wxd�LN��v�"E��@����:.�1������ق�a3�H$��9��QQ��cL��b�d2d����s6l�p09��w�8a�S�Mc2
ځ�KE��n�����w�Ȧu�����9�g֎P%`!1Ī� ��d6����Dq�d��@{�j��M�[���(�+�DAK%�f��s"��Ѹ;.MI|��PB����%
��;��:�;��`a�߂Q�jf�*�%�������J����^
�jƗ�Q��NH=w����f�p8�ύܽ|�i���
�M�~5\MN����"09��c�=�;K �W���wlkVI��Mͧ<&��i�Z\;#9�,�w�t��"w
-���Oz��1f�������źy����]ӝJ��� q�|�����mb��ؒ���K��B�q��Ǆ�ú	2�N���L��'0e��,P��(�xB96� L���q]�0�*��LYW�nxI9�C���'}�z�h$���4Is�����γ,�i�f�׆�������7�YڢkN�2���w9����'�
	D��(�|%��o�4�S�ݬ�cbO�ۜ�}�K�[������ε�'1J�"F�V��V�ߎ�z٫�[��߾b��Rrd��)C�!���!����0_��ػR�Z4�W�7�O]U�\�艀��CȀ�ڙϹ��K�ݜu=&�ы�$��rc�B�)�@ ��A����q��O�:U�/7�ԎX���sOVӸ�&�Hh���j�G4g�Qp��yX����S�b�^��A-.��s�̴�l�yy�Mj7$����(~�}�k�^��=1�AY4���ߟWh��6J��������׬`�W�!`�y���3�h%�LM@�z�;a�Y��ҝ�m˖nȬa�{Ho��(��m�K��w�pYҒ�?��fa��c��ˆP�^]�y�Y�z0?#�Y���,-��	����Xt��A?�f�R%k�Ǆ+C�ns&�s���]�dՅ���CsT�&9\V��p�d�z��0����P\��wh��5p��5lu=N*|K!�ñ1��'SW	0˂lm��jF�%�_w�H^���#����t@�!F���C�C����LH]������Ѕ�gsvIy+i�&�2��%��JF0�W��$�)�b�d�gP+���#j�y�KmRS�5� ���ǩ[��G���X��.P��`�1�ϟ�0�?G��w*��Aq���N��;-�w�E�P��X�,kb��h��2�@E{�c4SN�Ip��/RR"��L�G�L�(�R8ѓ�<�mηd,�t<�C�9'S�<�X�g�I�b���<�X������w��)p��v�[�?.ZZz@�P�2%C*w�<�q�D���_0 ��L4p��V��f�X��A��"TVa�bZ:�Rf�� �K1jn���gps/�X���bQm��i��he~< I>����l}+�V�Td�H�#e��`Ҡ�fd���k�`p2�B/Iww���
-�c�;+���M��۰�\�4a%�?���{��Fb��8j�%�!����c�D�I���2Y�A�o���z��.�.hvf��|�#�7h��Ώ�f7Ika�akO%f�iCDln��*,{|��?F����G�Λ�1b��kO�d�X ��H�,��&c���?��Z�A$�
��>D�&�p��U�y5AO��#���K�Ix�J�E�"��Ӫ㞹��#�J��z1���"� s�$�(8���*ŧN�'KG��6}S�mN$�r��Z�S[�y/�C��t �}�$��|��"�@�l���ճ��^ac1������Ycɇ~	}X|�i�'h��?��e���"S爛3������gA5�_���h���W�TR/�:u��Ѝp�)*pn!�*V?�v] ш�Ĺg#n_����wʞ-���=�����>����nM^5��-�.b@�t#��Ea� @�.��>Ӵ����۔��C�C��d�m������u�"�sк����`�K��Bi�฽K����f)�8%�1�*���<m"^9��=Ę3t1�cZ��ؔ���i�^R�߂�)�[��'���[�8I�kM��6�]��ή��6���z��b�d����Z��qB�F�ԙ�1w�z�,��PZ�.Q�:n�~֢�,oe���xW�f����Ԗ�G�o��b\il=��m���E@�QA�� ��򖉹�}8���t?�w�*���H���֋�����(��،�U�J��״�⻵�D`� =���-�5ƛ��_�PGN3��c�75����1�V�WJ(w�"u25_4�z�Co����ُ�e���_�t���� ��t8��g�Q2ژq�R�������G�[��������� +��i�1B|��9C���@��Lcm�Q��V��pH@��G ��M�m��tXI �u�EI�˘��Jn&mO����[�j3��}�j��u�m�W�Q��B-�p��ekoFRO�s�2�Sn�y}����r�=0_F����nԅk����밧O8� ����}�O>[���pU��yjY�� if�����͚�&��4��|��Rp*+��B �n �aE-�H��h|�P�W�?!�%;/i�l�}#�9�4�r���Ax���B~SY��W7_S[�(2�5Z
l��G
�3�=�5��e���������y�\�T�l�y�F�7�ͤ���R�Â�r�鈶��Z �B��|:�>c�Аy�B#��?�j|�lx"*q4���O'�C�W����uv�X�GH#.�?GD�.���i7l��ݝ�_����-;�E���09�g� ��FvPS�उ�]��~-�E���vK����`݂h��]�I�[niY��.� �����5�)��p�p0�DL%�y2��bҤ�'p�I"�1�b��ԛ� 9�8�ު�o?���ufR,���H�,A~<0Ln��V��-AAL��K;]�#O�]w=�
tG�I ��Kn�W�):�����w���2b�]�N��	��}��zr��
���	ß�&�;k�9�Om�3dѥ�qF�r��,dR �/>��1�c&OE4���̃�?����GG�+����,���Z}1q�j�Tڱ_���P8b
Z|(b_���i�+��ᑺ_;�5'X;t�'�7�D	w���[-2� �!�;�^n�n�ŕҍ�?�R��aZv�3���������=��&��9(�Xׁ'p{�Gn��jy��@�&��6�Q�M�%<��_u��9�����~�y���!���A�����?��=��n�9��|ϐ��;��0��C?d��cJm����}�R�t��X�Uz�ԡN@2Ձ}��!��)��O�Lew���~�A�!��Vn�О�B�"[�v�����Kn6��`��/�D9.�7�lY�4A�ZK쩺����F�}
�947�2���j���7��̽-r%�1m`�ҁ14��l�`݈a���<@խ	�8�y?���U��}��~��`�w�����q����Le���VU�Rh��9���N]k{�q��S�n�l��ҩ];�Cz|.�0��ck����n���WXC��G�f�$���;��>HZr���5|���4TO�*�@���]E���\�ޕ�Od���z�.��<
�&Z s�sG�9\~��o �=|@���m��m����+JyP������ǒ�~�*��O���L�Dsz�2�M3����O�-�A�����1tKγ�f��[�9�Η������,��D�r��V�պ�������7��<=�#n�Up/��@A+���*�r ؼ"�����2�R���+�Y(��iv�2�TG�lI�gFO��kX�����?J�
?	��D#���<j�J�9�ĔE��)GL̉��ȁ'�[]\�
�Z�\=<�-��ˀ[�L�bO�iu��(�g���O��8����eK�^ُZR���@���Gh\`).H�����+�Gըg��e���_N�ѱ��Ӯ]�H]伂����H�ٱj���V�T&yU�؀%Y�:�����!�Ġ��EI%)4H��{����HW��O~8�:��'�i�$�b��M�m�2x�w�3OD��?� %ӇTb�1D)"�q->Yۍ9�p�:3+����ZCȸ볤�|�=G��z��3�Fx�đj�����ƪ&
t�>�͎�Xя!8at�1�)b"V��S��  ��ǩ�ډ?,��������c��67�c��Od�i\W���⨟Y�m	+~{�1͠3��Q��D�k������os��+��55�p��84s���2���EK�f�!�8�|�c��OF�0M������h�,�it���Ӡ/V��_���j�j5;���0�O���8�N�ȶcx�m�2�'	��ɀ��i�)�q�+���<1eR�iUl]�
.�/Cj0��U�H��.�����Z�	8�WB��)L�]Q�뼂�=\s�M��n�9�u�&��I�Yn�׉��Qh�V�\��s�qi��~��\�i��������LVV� ��uD�d�I�aj��-��d|ĵ�	���C���d����	-9����O�auN��d�9��%Y1ź�<JY5Nގ{�+<p�`䰘�}U������.�-됝lk��}�
H�Rؙ1sX\��s�	TH������n�r�N�?n�YJ�hG�]!{��վ,�5VΆc#;�e���իMD�j':% Um9q&`-�����xp�G��B�t��]$�e5U$�x�c��+��S�x�O�SSʵ��#�l�o���S�b�7 y��(�q���Ϸ)�Ͳ�=�B���A�m�`ֵ��Ԑ��gdN6ɘMo�N�>��C��%�Z�31��r�9C܆����M6�ݵ�.��U�y�>��:l�:c�Y۝z5f17�l��O�B@vu�ٻ=�����D�n��_a(�!��UX��gg)��/C�	1#1�p�JXٽ���~��O�>���FJ�g�������!x��&4��X��/��V�e��8dI�W���q��������ݭ�РvE�w?6��$>~C��n0܊Muг�@���TC�Pk����G9T�����]���ؤ����'e��;�q�b���D�9E���bj�v���ɃI��j+b���E�w'�k�m��A�Q���mΨ͕w�2���.���2�5�9ȉ�{��(@������q��l�5*9���o5�1B0{tu�:����PJ�K@tj�K[�i{\/yn�n'xg���(凊To�\"���6�	Le*���;���%��y�>UP�&[�wM�sm��A���p�e\�*�y��~(k(����|#4�$�,�����"Z��C�
Rp�vDw�V�cS��B�țPc�a�*���֯�<6@���M	MFڼ*N�3���MI#D	|�qs,P�Oػ@�d_�F�k�e]ڊ�u��9�A�>:F��}�^�sv�ɼ��r,‶bE�+kl����@���i�Za���kn��V�0�j���Q(Y�j�Cϥ48�nd)c�Ò�eֻ�G�

u6�nX!�S��T�?�|MGw�ܦ��C${Pv����m� z��|6��5�7�<�t�ӌ\s�����{2s��I�;PܮB��EwGvX��rs�y��x�Ӕඁ�;�_t�B��Z_��0�>�H�����#P_b� [d��`����N<��Flhz�������.4�n�DH8���J.�}A��k���g~[�v��,I[�6����oB�D���W�P���<�Di74�;��T�.tQ�'b|�� �MA�/�e��;�r�n�t��Iߠ65�tz�T�e�����<C�<���bta�n�ئ���T�K�dH���D�fX�Z�!����3�L�;���-oA�,
�/��z5�Xf�[J��];�����@�*?,���8�(��!�L�K�0 u��;�O6?�N�k�~9��P(���V�0��|�#oT>�8��q�+
n� ��?�.Eg3����(��V�;�����<̀�j$�0<��j%�D���ÇUX�7�K�|Ԍ�1!\����.���G��a���e1������1��wpUΙI�P�=$J���>W��S�����P�-"����1��7���y�i#��N����_�
�%t�	x����⥞��4��驉���X�T^v���W�z%�TtЀ̟Dj���,�8�7�S�\@�9N����W�Ӧ ��C���,��V�kCz������A��eg58�V<q��M�>������=��C�r���az��B�NV��&��h�p\)�oX�[<��C13��ES�s��&�V�'}ePc��S�+8)�b̀��8C���8�n^jڝ#��c3o9��r����X��$gƚs{[�M����0��
�n�<c������s�/7_�C{ٻ�
�" 3�V��k���O'�K�-}D	;�kC�{�bn#�gAD+	�ge2�0|X0֔_bT`Cq�NUL�^@k����M��.�e}�!�IC�T�#���^k}��aY�}����͏Ⱥ����]�/{Y��e�ŋ�G	q��ҝ�� �q��k�"��7;��,��bq"�μ�k�Ep�1gG���:��|"��(V��/`0b4(�q� �cv<�p7�#�z�x�/̖�+q�(�ڳ�� �E�&�>��+^p��Qjw��[
��O��ĉ����==Z+{p�荫b2)�ַT
T�م����\��Lݜ���̕��	S)Ԣ�^�r�+����4)�����c��3-b)����nVj�ʰ������V7n�J�(�a
��zSL���3��o�mo" o�,����"|�ѕ*E��ڿ-�!<�%�� ��Gp��O�D�:�ht�k{�ުc��6F��$ ��TO�r+cI3�ݎ��u�IV�TZ���u%ᩞ�ʈ�V;��E���x�}\e��N�i�^]�����R����oR�����O,?��O��7_֜����lbS���	��O�A��<
Z���.,�>�H��� �VBdO��g���':ɰȑ5�=��xUw��L� �$sy������&Q�}��%GX�������l_�34��pr����IxTBDX�,l�,���L�O+|-8��u6���?�闲�̒�\�_��]&/*�MTM�S�����X��ȅ}3.C�6�� 3g*����L��'~%���&��珣ع��*�6�K�[��(J��;��������D�g�cǙ��'�̝����T-��Z.b;J���u�Z�t�lX�Ȯ��G�1���VP�u����;����xu��?~�X�SbPn ��9>Fƺ9j ��g<���-��j+��cM��ڰ÷F8 ���Pr:�hA�l"1ZE3M��y֊m=�y��Ԝ�������TD@����"�y�\r�ᦀ�Eº�<����s���`�%+��r_����׼=O�?�g�?i���b�z�E���3.n�n��a>J��MDG�9�Et@�O�X�����3b�eLQ7|�=i�=���P+��Ɣw�Yb⩵��{��twc+��ւ� |ů��)��Nmys9�J�SRA�r��i�I˴�d���~���l�x��i� ⛫I�^�lU����~iJ,�'eV�cB�?2͡6] I�\�C�&�����(34��m��-j���]gj�߰+����/�����tr�Z�F�A�m;�8-�%�%�k����suޣ"E����Xs%@X8�d�lǩC?����w@Qc!ՍG�����������ă���&��]z�zs�w��=��K�Ψ��_�D��mo8FU^W`Fz*2���	��`�屝Ъ��=jI΢�2I���0�����s�ދ$����Z���Xvf����(�p�fm�@	K�g"�rӕX��	�a���R��Zn#��8�V��2���c�+��~�6�+�ԸBȵ��\N�������A��f�]��S�L�b���i(_�m�}�����NO����A�Z���3�w����fk�e���i�(t�0�	�7��T���x�(?~a~ęB��&��`�i�[�0
龾1ohM ~�X�k�d�ɜMO����cY�W�ׂ1�ݯ+��1C''U��"mD�ó�	��>#����G���z�ކ���q<�=�Ӛ�V(4�ϑTaQ�S?�o)HVd�0��*�� �+����8�W5<{�s�ވ�J��ǒ����.� &`v�Ͽ/K����=xD8��s��x�P�(&�n`_�:D�u�V�����u�������_����E^��B]e�5O'���*�������)�y�)�A�-|͵�%�9k����=��U��`E##�6(b�% ��$����N}��P�����:�$;)ˆ����5m�|R7��NP!nKPl�Kr�W�V�Md�>+�ņ��C
ka�J��r��"w�
/���+�m���u�qg{/+�g����]OŌr��x�#�9��'xSb�ɠ�!���ڋ��t�ҸWu%��΃9���q�Y�y1���+79��P6�E����Zn�d g�;'@�H��Q)�:�ooX��7���L��H ����oj*�ڡ���uUuL�du2����Gl��~s�XC?Na��j߉?՚�dL�o��HwK�N7�ri,�j�VAA�ޤ�u�R��k�~�j'���wsHr(�/:��Y�Ml�Ad?�Ӱ��# JR��s�N~����R�,�t!�����M��?kZ�-?Lu�>��`�H����s� ������8ҷ"}.�P&]�p�wW��V���(�`�u��'�5�/�QK�V���*,����mC�%�����lHuV�X���
i�0��/ 	lU�O�wz�����i� xYL4+e�*��memZ��\-��~'��r���{���MkP*�����O/Pm]��'�\u�5��kd��B��/=�=�T]~!Y��X"z��a��NO�MD��~��K���
Xo4�:R�A,� �_S��W��� j`�������U����FZ�a���n-�Lz�pK����Ĭ j���b2��&2�"�a��M����̇D%�$)ϛ.)���Wd?XEcj%X!O����j�_�� �|*����l���4�����HS���v�O�{Ѩ��+I�7��������������ĳIEe!�x�qX^w*��( l����"�S$�`.�������&-u��O��\����x�>[x�0�,P{�����T��G�(M�![s�s��x��]�b��kT��D� UX�9|Hޛ��Ef�T��^�*!M����]�oEm|X��P��O����ێ���H���H�<7%z�o *��M�s�*��cE�ys�=)|q(r����z]<��i>� Ac<~�;�N� I��^��=��QZw��5�`��Fi��=׿&�Gp$l���L��&�j�/t͘��K>�z4�Y4��-�
h˲�/�l�-ø�]9����
���Hz(u�>$3�O�I��~t��6ˈ�)2���n�����jG������yS,��w��$X-�[؆�k��J.�\|�8��K�n�Y�|,�uw���˜�r��6Ij��Ʈ�k�͐|�y�c*�wI�i�w(R�x�\B7y�1�(��ꥏ�󛪚��
4�H��0�G>��ʆh^vX���?���Q8�����s�ur�LOc�%���|y4�b���9�PX�H�lpMW}�����tƋ��/;A^����C⹶�{	m�d�Ɔ��0�����ÇD�rb�7Ӳ�0Q{h	:� }g⢮	>�\�B����g7��Z�be����wVP�	/��_IU����右-�w���!*hS��x�bbs^^��8���o!9uW�B�o��8��X��~Ց��d^B�]�e�����H���+�$���gv��)���H���H[=�_�~Nպ鬴O:L@��l�űW#��^���{���� �������V��=�0�`���(��O����� OI��+���\�&��T�kx�8�N��r7'c$2�^���p�x�#��n(��h��l�Pht�Ǝkr	�پ�]��Б�A�m-��W��%T7,$���Gm!"Ѯv�E$�y�BØi��Gx���c�3�@N��̠e/T��3
��@��TY3�W1�E�]ib��f�|�����z�� �~B�TTܟ�'��c<6�d����	i��'����jJ�5��|R<��돤f[Y% R�������ШL�t�7�D��*[x��]�S��K�m¨:�������ZV���3@�J>4�ǫ\�����T�6�k���h���p �wC�Ш߀S���=�п��@x��F�L����Eqo06ӏ�m�r��|�����C��ø˔�rW:X�fW�۪�K�t��O����5I "s�i�1�2��;Ee�R��m�j��{�7��E�]��%�N'�_�c{U�����UaI��qs�kS�+�G����� {飕�R�B�(6�0p)�O��᝶�غ�z�ˑ1�k?�}w��� �DN���/YR��wO���ny�L��� �*�����H{@��f�c4��x%����1NRO�v&�<�E��<�,4�[$��g�j�n�H�E0���@N���`#�&�YPV]�r�b�ʆ��<*] Q�����K<�E�z9�ҧ��V��A�E�C���:2��z�� �!+G��43z��֘F�U{�̀O�$���
t?	�N��LW���n�
h9�_*�29�ض��BW��-���,~KƆ'PߏSچ�Egm"�p\� >{ԛ�Z������R~��'�	6��rW���jS�qd.4�/}06	�@��4Z�k�Ҋ2����F���Eb�F���e�G+���B�>�Fv���Y��-�Vk/B"�~\��七)X�!���Ri�ٮ;�/}u������XOt��bJ���E�yH��?Wf��&��>@0	OJ,a��d��|�7ű�F%D��k��(h@�E���W�Yc��J�!�^�)q}U�hd\x�"��,xpV�80�����rd]g_�a����)�jƼ�̉@�s3�9z�������������U���BgO��e(���� ���3�ө�>㎁ Y��D��"�*v���݉b�2�teX�����8�������[�����2�eig|[�Ս�9۝��Eвw{�¼
�������͑A���V_���	ܤw<��?�#Lͨ-�%�BTp�Ek��!I�tq4t�ڋ&2@��NX��:���w#��3'�Pƿx#>3\AHl�~-&J6Z�� ���@G�nr>8�cQ\�tb�$�*�F�ڰ�y_c��=�G����<B����_�סHM[���)I��~�$9/�8
W�Ɯ�*_esy�m����?�8��+���D�O7xR�zF���^��pU�]�aY�Y�cX[v���(d�Y]�R�Try4�m8�.�,!&a��r�vF�+h���bwP��]g����$�s����}���?v�Y6suIyܮ�{�L�MD$�� |LT�1����pT�o[�ij�8r=O�3s����F����5�5ߘ�~e�U5ad2�:u�ڲx�Y5���TXj�X_��"ߎ������Oʴ}̠�:4�bB�B��gP�l���\o
�^(�,�F?B{��%5h f/������B���� lqVI;���T	N�@��s�@��/��U�(�9�c�]��>U�:���\�zS�Kp��E�?f�+ j �����gPrM�Ĥs��」@P[�n%�tV�mh����v��k�I�#�/c��["��M;�W�蝴�-@�ϻ.bY�mJ0aOz#�1��ڽMg+IQz��:�]g��h�c:�x��T^��	�� N��Z�H�E�E.J	0������A�8\$>AW~'rE���_�C�,ǥV�(��X��#XZ?���(��X��A�m�W&BQ<��.\\�ѿ���gja�4� ���?�M-܄��o��b���9-g�]�3B|bfc@�i�8����"T��!�����9$��Z����#.���(ǵWG""�{H��Š�X9.���d��<G���WTm|օoՑ�C�A�S!;��VmYV�6�����d���n�g���I�r�x�-7d�]�f~0U�zc���>�X�ؼ"{A�N���9��4.yA����"d۵Lʃma��zI��R3�������N��l�p���E���>�d�RJݓC����SA�#�\�.���*�Ǽ'!bTҎ/���4@ŊZ�r��E�? ]N�L��ю/���G]���&KSe�8�3�QnY,��l�{�j�Q))�.`V�5���f��cQ���r�ȱ�ъQ�'n�R�>~PƧwD��!������f���!M�#�%��\E��.ď���4�(���3Uk> ۠�X`'Ȗ����S����Fv$ C�\�,�D|.�;*;Y�"ZW��0Ӆ*w�� ��)� R�K������������F�_?����1[��i|��IKl�&�{_i�{5.gP�<擮�M���d��^���P>�Ǩl���)��y�����/��b���e��r���ę�zj��)�$��6�m!}���B�N^�O�>���l佘�
��!z��.�2,�r�m_
�sh�ǂ[���`4����6�'Y�|���Ulh8�_
�fߛ����.�Ц���i��sA���L ����~���N�H7Î����*Cy�$�`
�	1��YG�J�,n���N4���9����m։�/<��,�W�� sⰉ=�?�{�p����#�.�4�AD��F�>�
.cT���OR����h$���#�
&"�:�b��46y��f�w��v81�~�t�
�&0)92��s�v|ۢ=�𙕨���C�כ/l�c�҂�6C(��a�*ϗ7��
� ��9p��碕��J�=:~�X�A��!��$iWf����Kr��>�n��Lihb��bT��>���CP�<�����B��4ʜ=C�7�a\w�$�;�Vc�!��H�\~�Yf����NЂ�%����f품�I��b{C�0��Tyw�nv�!�����ݱh�g�y`zWq���I���۪bVj�Q��нolJ,И�.�����E�̆��V�3^C���PW�����O�I��&��d��v���(��D�[.��8$x7P�ӖK�K�����$��w�iV9yo�)���]��bC���.+)��C��Tj�꣩��Hveǆp����?�E:�p&�G�]��N0n��fI�����p�g<fٱ{Q]"�9/�i஑���v��fxV�*���L�vh��w@��&:�5!
�2��n,�ޛM��S������.T�	�U
���ٶ�	\#����7T=�T�ʭ:�v�n<�.o��C�⁼��#���$w}:̵���T;ؔnɄ�ƽl~&N��=|�j;�ëTL7�0�s��LGƋ�ϟ��Ǚ�dq��-��o�φ�#�[�F�������1Gmn֔̾K���,�:�%�!�#?xr����� [��>�cI09J����n�����
10�6�J����-��c�y	�7n��&A������=�FbT�d�M3Xx�J)����Yg{�$�nU�i���L����Rk�T�
:�����	_�-�(f�S�8��ǭe6i@թ�hY�U���PQ�9pBQ��q������'&�PU�
m��Z}�^c��<ej�l�襏,1�����#��9t��͵�zHn;N< 0�fD����O�w��^���P떉�| ���؁���Ư�ͬ̄���5�e��hxc�����䋽�����ـ�a�,�UV����9&k8��������\�ێ�B�/�d�-
�N(_�A�����Ly��X��ۜ R��{�O���ar�1g�-Ŵx�
�/̲���q�˷�D�^n��<ԸĂ}�/����M%=�.�%��cy��!�ɑ��#E�|�� ���L��_T��q�!"`e���5�>W�)�-�.Q�4M���S'���~�2��{�)��|�e�tv\�;���c�e��_燼����r��if^Fm-�8���r�A�}�/�������Q�˯c�|CKtD�N'a���
q�o��B<�G�sf��g�E&7��HLJ􁠆z�V�nkCIK������C���xe6��_!4g��r�F��AJd:�wٖ����	����+����Q K(�w�
�5��.�H �4��,б�/wA�I��g�� b�:�tlm�#luL��Lrw�L;s�������w(� ��y����]�e��
" ��/�O�V?r$w*+��M+J��&o�#Ȇ��x��Ƴ��;��N߅Oߴ��z����D�;| r�"\R��ʯ�-ɬ�K	1$J��3^��K}�<�pg�Z�˶/PO���Y�I*��ƿ!� 4iH�QY�H�z9�$s�3�[�� ���H�yM�K��3����4�@L y�)Rk12+R*��(�c8� ��5s��7�d@'P߁b��յ�X�ʁ�a�z��tP����{����<&�&|�ךa�ĵ\��V��1=*�NDA�bt�!���|"0$����s��cX�KyKx�j�v?WY
����*�GX�d�n��˛vjOC� �Iw!�@�#$`w���f���vp�G�͋��+Rrq���J�H���
�9#|Bsh�&y�,���� !�B������^tte^j�lǝ�{��N��T Ŕ��������[����<!�g�Gi��Q�7\��,��������D��G1���j�#,T��!o��Ƽ���M�8�fM�\��Hrڝ�8=������i��y�/-�RD�9�^��V�v��B�VaC6�� �fW4W�:��ͷ��N�w�F(M#8E�퐆�\���G��g4��_i�p>����v�ά��j�5]�����zlqz!��@��nں�*j�����l��	m�x���^�Gչ��r�ߟ���c�Gt�i-������'�����Jʁ#s�xD�ބ\����ʭ���9��d#�D@��*Tz��_�"M�:��R�"0���J�96��!�Ǘ���҆�^C{�KV���y�ᤂ��"	����J���ׅuԂ�h��5U>#T棚�l\؂�Af�X����Ȭb��B��H��M�2��qc��5������%]�z9R��p��4�8f:��Z�����	#V$�㊓��!LHFM�o��9*�<���x�QQ���w�H�H���S;���KoβM2&X�[ڑ�+��xA�ƒ����K����ћ(Z����"�QѺ�q/0+k����Ռ8afu����=�tf��pS�����U�F���P�j9e���һ���Y[�
a������8��x� �a@:P�$�_+�i��י]/c�z Γ|]��������,yo��Hzh2�V|��
��D�E�
�.����!w�/x����.�A��^��>Q$!6S����G����r:V�����~󦇕�3���;�#�����~&"q��<�<I�L�p�t־;�΄�/K0�Dcڠ,ָk�A3"��WN�k����>cP�.s+��'9��썋b$	�k�ܐ�3-8
g�G�\f|E��j���v��r>]͗�e��;MFx�$yt�t���+?ܩƶ�F<�I���|*�!{�@�j�����o���8��-�W�N�ǻZ�2���p	w�^Z\�|a1�k�}�B:Z�Τ��b
��( ��+��P����)��̈�Dl���a�3
S��-��.�c������ͣ���]�n,#���s�uk;�T6+�G���2��Vk���%����u_����vp:��T���� �j���;"��[�� ���Oh�u9�fѝY�Y��j�w$W�*r�i���y=�
�5:�IkjCm��C1 ��"�l"ҷ�����rIS�݂T�7���|w_z&)�Ci��j��fH�C��������$y3���ID����ƹӧăG]�e���*�d.��3�({QJ;Ư�A�1���(���+��k�3 �MdID�G��%�ˠHK	}Ƥm�z�� ��cF�i� ���3�xS2dd+$Ls"{�El|�7&a���F,&�u�e���)���́�K�`-�������QQ���nfD��'�B�9��A�H���WQ�c[�w�Ǘ� �i� �GK����B�E�e˶/��Й�>�KY�ڭʩ̖�S��eb����3�$��Gœa�Vy蘴}1QIi�|�
?y�X{�A�Ͱ$��k�
�I���������Z�9~/E0%�	��Y���w�}�W-"MLc��r�^!�R��)j��j��X�ne��{
=�F�,�x۝��ZG �f�/�[����s�qR��N�و]�&��I�Ur�c}��FmcQ�ĕ$3��8=�[���E��̙��<��x�����W7�N��Y��	�hɥ�v�k ,��/���-����;Ɉ��}��������3��vIB�~T�<��|��H.����� M?*%�>����.@�B���#��|U��3���ʝ*��F�s��[��oʔ��~����P�M�w�]<��-B��#\=B����M��.>k��M�4OEl��*��N��f�4�-��^I�Ū�@Sx�i*@?��X���3.!���jS|i�]l�����l��E���
1W�Fb׏��R�x*6h{/��c�Б��Ǆ�(G��������z��Ӈg��	YMx��)x-�:��9v-�h\��_c�!�e���"�k�$X�*��l���䠛����O�\m����������Þ¯'�z��:N�S͠�)�v�Ӿ�O��+6`O��S���-@[L�8������f8y�㡰�7/Y�y�{y=�2��^���R�pN�+�}��͎]������6�&t9��#�V����N"p��p��*"�����F�(1�!�U���>�+�Z1�a�����P��\�� ��j]e�:�xU��F2�P��B�7���
ø��V()��F��/ڒ�SYb6��_��V���ӆ����lD~��-Ø���	C3�6nvdkt�ƾ��5�_b��	��f�C�n�%+���fQcJ�D<�C2�J^��W�S�kΡ�6E�+�f�Ow'��� ڒJ��&��Xrh'�m�ns?|�$��Fź�Sڢ�+ӟ)�1���b�*�XO��Y�W�;�;V��7�Ch���:����t�;�=�l�w�p�'i3�G��s �x�h+�0��s�	2?��s<G��A
�#b�}�%[%�������g�"�VhF��n}�����A&�V�vV	�eoT惬�CDy<D��"xX�jw��ž'��y3WaP�"�b4b�cd��<wQ����_�_r��Y%B�s�Tsp�k���)�.g����[��$D*�9@�X
sV��+�x�'y�[p8�u�+�c&�G9͑��]�d��wXڂ܍yI��_�|H9<�q;?�H)|�:<.n54��d⦌�~��ii�l�K3YQ�Z�6!�id_1���ֆ��Q��K5��Z_���6<>mz����gQ�SZ�u�1���y��f�
��S�~*t��0�x��ˁ�h��;P���<�l�o��V�L*�U�Q���_T!�`,���2�O,����G����h�ǋ�c5,�xA !���%�P>����})兢�mOj�ă|I���ix���f�2��p����ߔ� 4#����=q�ª�pe0��\���ǫ��mv,�� $��2b��PeZ�m�e�#�`KU\^�x�u&`��H�>��媛����7F�D�+:���ט3G���-p�qN�hB�Q!Cٷ��A�i�Y!лPuM}�Y�o7@~C�E��[ĩi�[8�6=]��~�"�\�U|�ڍ�A�F��P�_���-c���?���5�i���$F����1��9�VR%� v���7š7CI�6�������cz��!��X4��sr��J1��ӂ��m�hN���WR�Z��_!>}����iL�۵V�;5�9�8�1
5��=',�֩��Hp�W�n)��س
7[Ɇ�|Z�l���Ѯh��C<��G'w��O	���꒸��S^�M����ihg���֋<ؠV��!J;A�?-�68c�ՙd]����p7Ů�u=���;Z��$)���&ۓe�2����5I���8f��J֣� �F)�}�c�sc�wbm��؏�jYg�����;�9�@0��(CAa��!�3��������v��gF�
G4"�Z�^�Ilh�t���݅k��^]h�D�gcX����*��?;�������wb���9n�(����i�R���Ɖ�=掆��D�$�ʶ6
�,�%�$�yl<Ci|C��O����m,�\{�hP�iqO���qD�kұ���� ����
�D<��=b>�� u�Hp�?�?�M}k�W���	��:�Ȱ�J�s��/:���i�j&Va0~"Gk��9'"����Z��P�:M�F!���H��m
bK��r1[�!5	F$e�o�?����[��~�̯m��	m1$� ��lC�>���ً�ܟ�t%��kW^ݨ�'n�9b���N�~L�|��3͢c�JI�����O�L�6P�[�U��Nc0��| .+���EȪ�M+Ǖ7�4�� ��ga�;�����PG�=�{��>Oe`�sN��ҷ �Ǜ�3��t�!M����J�8k��^�A�$d�;Gt��P [�g���%�d�0�M�V�C!��X����2��u�/)�s+�w�5�8ӊ��Q^�L�V�w�}��<"Eb�PD��83���R>~�u�����CV�p����8��@�֊УV$l+]|��n�,�+��c`���C���C'�z#�O�e��XaxiU!�%M�D
��0~���6Ɲ.r��h���w��k���"����8�j^��dP����e�/�p�d1g"���탄�T�4",�4�t5�Dn������0�9��6�
�FŨ��$&*36�[�~�|�s%-��t��֕�e5�E�)� d��@$Vn����Po�c@�UB���d
sg+q'j=a�{�t�)�5%{�f�R�Z���%{���/��v�4��ުM�{��d���*��"Xq�����;U�s1�t9��j�N��+�	��E-,H�����r[��Λ����{6g�Ho.�oǧD���`�dQٖ$�P)9�I^����7�O�t�,�	�Z/�@@��'���0W���[���c�����0Y�ծLL2ھ�KXv4����C��;�����M�L[���~���a�CX����J��ن�\Q[_2�G��v|I�˩:�R���%�:QW��@,�I`�����`ۥ�ވm#	W��L2��A�4B[�FU���e����������Y��L�v��i���q��񗰃W�5�o8�"�O�-ik#�7U�������yO%�<�k_����v
�"�7ʱ�	h�L�5+ ��oY8�G~WǏ	t����̜Ώ��Ch{kQ{N]�AMW�AԀ����_t٦��V:IWO	��y���N����~�B;�^�	a�K�d[����EUՑc�FKOj��֡�e�	ݾ�.��V�8��~�Iy��RC凜e9R�����)����{�|2���*��)Qގ�tO�5��:E~��)�ú{���h����~�M�T��>Z<y�����C�&)�x����][��m�o�F0�m�/�־��l�z�I�����u+�����\v����.b��l��#�E�($�%d�!&����$(_ǒ���mI��*8��^�:"wq����
�D���Y�sm�t%�g9.<8ћ$=P�o��C�;�6:�J�J ��q�;G G�Ѳ&�Cis�r��9Ay췙�ԕmS����&��������!=J`�;cm������G&���.@!l%bh�C�.��v�/��xʴzC�a�m����C/��[�Q��Ī̛(4��Qgo�g4z��I���b��$}MW���� �nb��������G��
�9#���� ���#�S������1y����[E6 qI�.Ϡ0+�}�0M��kW�t�ҁ����k�t���a=�k��e˝���n�-S�p��<j���2��Ae�E��)������@��	�f��jЏ���Iޱ�-	��G����-w�ˎg�O�@��}WH4���o΢�9��O�\����8�*R�ѽX,Ό:�%�߄	c<��-:%=����� ����$O�zG�S!�7�V�Z��j�����X=�@fyl^*��偰��:��?,�@-"D��
R�� �qe8���;��\X�X�w�¦I4'J<��>��j:�����p5cݔ���B	�����bf���4ǎڲ8�c8
f\P�{�Ҏ	�KR�KҔ��ꢑ�`��\��DW�!<iu�\�@U���_��T�7������f��b�2آ�Ǒ��@�|?��ˇ��n�}�|���`z3� ��`hw�ȱ��}�q�|rW�E���mѤQgs�F��St��
�4�7�?@V���@h �^�����e)��b�ŀ"�R�q�q�;H�2���}�*Ĕ�I|�ٙ�����j%!_2�*�ԍ�v����������T:�I爒A�pIKo�����G��%6"�NԑYfF���Y�����oo�V�I�J��L��K�j���=�F(��MD����?������a�����(����������P�?Vщz�Q�`g��F8T�^r <�k���t_U6K�iC��~n��$�$1�=C�[}^����e�ީ����e��/T�L�U�H�p�B���z��X/��g7�_u�L��)4����a�\ax��M���k_)�d�d��s^��M!�V:�|Z�cT�{gǘ��4[҉�$H�쥮֝��NhR��|4	��J����2�!I3�%H���U�Ͼ\�X9%;V���y-j�x��m|�8����n����3�Se<tUM�/�7:��0��.�=0x���1ɋ��d��4u������-�H-v2�8~64ԕ�"K�/M�U��g�|��(ʹTs]��;q[	g���7�pio���)vs�Gr��K��2g��h��w#5�)� �+�P�+_c鴬���Ҧz�Ro��D-�haS���@��Oo�iz�Z}D�V�r������7y���o"qC�gqF<�I��o4�m�_�ﰑ_�$��1��Hn�v>JzْcLo����O��"�Px�g����V�o��� ��u���Aq9R�<�n���cnb�<5AS<|��o�W2���@u2簊 it�C�ϙ��^d�r��"��\
2g�%m�E0��Pe��¥�v����J��w�����
b֡H����"
��&t+���0���5n��H�._�Y�`��R�͈�͎*��z�ڭ���@�p�����S"g�{w���z�u��;���f�ed[��p�2�2]ױK�0l(vA���~�`�e��V�����X2A�|>%�r���/�hh���j��a��2�@|O"���qƹem\Aib���̹�Qﺉ��x$��g��a�^�S!����sF&R��6�0̅����@p�������	�~M��y7`11-w��o���j&_\RS+���0�VU�`����@�"zL� vi�H�m�6�������2?$˯{-W�1͟H�]^*J��T����隙��B~֛�k���SP�8Ĺ$Bªj��w �خ��$,�, D:%oK/��a�O��{x�#@+w�P�C�Ľ�d�"q%�r�WKh����L�!$�C�H1�u�W�@��R�>���\�s���������B����@�B��U ��B����?b�V��^�!�f ����%>Ɔ�T�4���g֭��~��<4��,���:vT
Tc��>��u�C��#��H����
u�h����)γ�B�c
^���)9�o�=��G,G�����=�[��ۺ��S]>���ua�����A`}�8xVt�}I��� ��|�@�)�N�_3�$8Iy�4Hҵ�ӗr��cO:)7� 3z|"\w9Y�3���J��Wz�������P9X����t�<��1P[�����r_俙H���޹_�GÉVs W�d��3�r?�i��ZܬTIw�AƇֽS��B �)ܔ�r[u��o�c�K!!8����Ga�Y/U�}�!�1$�D��c�<���t���$�������v�����yK��1�jl��̱o �俅���H{�}ְUI�K�Yu�MFsl��p��bU�[c���W=Bp�,im�� ��HMdbE8��NkP�̌�ʘj��˺��N�	c�������-w�[�L>4�w��i��9`ސ�pi_4�֗�S��5�I����@/>�Q|�^��|к�1�����7�H��5c�r��ě~�z�oB��,�B?@���p�p�5����5���k�$���1v���L�O*��:z��P����)�=�4r�������y�SE݊I� �S�2�q.�:��䓼!Ia	״U!_wVrYw~|��X^P�.��>V�{�`��b��$���z�M�{3�Q]�����q�	�GF�LҌ@�矑�lir@��P
VE�\� H����f�eQۿ�{���ܽ+RL�>2�zj�a+�J�P?%g|y�� g5v��a?�@��rHZ���r�J��� ����g�g"����y;|��j���2)H�V�������
���=�DiXj�2��Z :��:[�]g=l��!�P�A�)Xf��(1�m�����b-Ď��H�0.�Ky1��V)G��tԁ	^�/|����3���2�mk��o�S7K�h���K6��@-dN��v�������Ipx�01�{���<	0��N�O):T����ai���%�Zz�k�$}��q�f����b$ε&,�W���%1qQj�J��w���`ѡ�q�����H�%i`fv���<#��*�ߐޣ��$]XY4i
�ؚ�J ���"�U��ձ���P3m�4�m�q�U���M�?��j��I9��Q|�Q��&�jtg��v�:�k�P����3qފn���U�����Yw#�@�9���3gIկ�وX�pL����d<��%�Af&��щ���vp,s�����̽���Ҍn�jN�A�/c��b �@����1�|�2C����*M�FO�J�G*^������}�I\ '�p��������5y�zj�$�c�#2���ա�!W�2]��V�eh��6� +�9�\_� �a2�0r�=�6�	�Q16�/$��z2�9�<���B�,I�jf�tR�߾��Pe��?;e��R�ӯ��A����<Q�3���N�jz]^�?<Rmh�q\!>2�5�#^�{��c���(�R�75�����=}�/)�1�4���r �/�SR(dg��Ut{s��6a|zz�������)��ʳ�@\�m�����1���jhͮ*ƞt���/3o�}�2JN��7F�@���b�Y�=��2�����Z�d���H�f儑.��h� ��g�BB32{�ь���|r:٭�6�^a��b�"&dv��E/jHF%�c �Ó��h���N�y��d�};Ȩ��P�/��s�&�y�[�%��nA6���2���%6�>��TS���/9�ig �d�^:���wl�|�Z���e��Cx�9þ�V(�y�s��-�Nc�ũ����ld�|��ڕ���;K���eS퐁aq�I���S��;?k�$��dX�T�6���&���QC��X23/��6��� ���H�	hD�n1�
� �����͠*��?1����֚������3��O=BN����FO�%�&�_ Ezu���k�Е��N���!�
�$a���ҋ>Y�(K.�p.澧�����Z;�Do�����dz4����=J��������9i�ç��b��Ƿ��m�d��*Q�a��I�x�^D��}��3��3 �� J���w�F���Ϡ�FHG��i��:���&��I&�,�:3���
��a�#«�z����?�k����`w���O��i@w��-�6r{��|���G��JX���Ӕ�ϕ � �Z��oP�
<� _�
%�~�u$77�ʽ��3vO��UǱ�u�!�'zdZ����[^ �d�(=k���Y�$��`�,�a7���IW�V޿�z+�P��y��������+j��;�4ip %�$����:B����y!�R�\ Τ���`��j�B_����˕��,���~�y,�����V��N[
�I���H�Zˌ���? �Uyk�|;�\�g�=�d���8�`�<[	�<���z��Չ8���*��+��d����Z��>@1N�?�[겒�<�.�E�+��������pi��8h�V?Zn:؇��e�*�l7θP��8�C����b!0�~�7��̪���un�J�vo���"�RsE�w����+*�Z���Й�Zv���W~��_���T��'��:6q0��/��Bh��E�v�g�(MP��G�;О�1�' �e�/�{A�N�����~�h#�*&XZ',��%[��o��Z���p;��N�FsC8R�f��Y�9%p��P��k��ďՕ�MTɃ!�#��)����As�֠e��A�Ib�AR�3^��Erz���2��F蹄�m/��)��@=�S�p�x$�d!|r�����@etO�,�x-�ɡ�e+��A&��(0�UoɅ;��fΟw��gs��Ń���lJF���!����E���ph%�Q�� 'i�|��'��3��u>�4��i�i 
��j�7:<gى�K�H@��� ����_MPƶ�(涫� �^x��;����q)�m1l�@�3)�bV��>Q��G2�-D6Y�ŪQA>��a��(j��=�]�\���S$�ڗ ���c�� 2�U'[�� 	VtwYe�_�֕��D�wLW��s�	�ՙ:k��E3o"7$�s�li�� �Zu?��cB$>1�Y"��$Gr4������WICZ
�{E����U|�p��@���F�a<,�9�8	�U!=���L��pT�2l�4��G!?_t"g<���SM|N�~C�ee��bnZ��n��"FwA��"Tb�p����5j@ei9������Iii���MU�FӖ�L��`UD��ԊW���Q����=���Lk�i_���1������
6�c���a���^��y:�j�śU,��FҚ>T��I0#��<��jA^�s��_ˣLg�Q�-o��5��t!����Bٍ�3,��`R�(���I�e�4�(2S�gBUs���IKx��G�Y�9���z=w�˞J��@:��������h��F�^�_�7�3E�k;�d1JJ�"�  ��g� �W+#�~�A�]�=Z�3��K~����I9�K��>� ��;��%sY�z��ޒ�)W�
���#����e*����|�y�u�M�!�Y���Ӯꚴ�q�٫�����j�9'K�����`�өɯ�(��n+ ��]�u�&Kk��S��L+N��6��N_rc_3F1M_��eBf
#'�e2�g���P��yM}��W�a��ȅ����P�bs�4t�L�I)'��Y1�IQ[��>�ۘZm��⫓��]��E���2&���w���F�T�qS�uY����r+�B�7[*�J�y*C����?I�hOkB��&.Aڐ��L4#�
�k��>��ƅ&i�K�AW�v�`�; r�t�H�}*���^�P�RW!}���WpOna����8��Д��M��P��b�\����+��}�d�*�+?�y	���J0. :7��V���M|g}y�����PK�Ā���A&��_�E�ZD�.7���L�#�Ba�b��-.���<5BW%޽iU���D˕̀�z�z@YU�g�F$�k�s�oJ��}����e��DXl��A�;�ՙ�$G�m�n`٩�2暒�K��2^k���cQ/��
�LpF]/�M�l ���=qc��!��Q�*z���O#֣�Ħ�T��]p�94���n4�R��v�X�>����}r@eNh�B��ۂ�e(�8Ӂ�꼟I��e���t��kH��ti9&w�Aփ�C	JXfQYG}ԛ�ʍ�r�Jd��V��o�(?���O��Cm���'�&ZC����%c� �&���2�j�#���F�I�i�Y4��j�5�#���^4�޼z��d�|>,�� ��x8�+��L��n��	u���5�\��a�=��Sw�?]@޺�(��·w�ǒz�lHV�6�~j��U�(�a�2�L�1$u��@B��⭇� ���F�X��t��T��\��X95G�I#��-tT;K����~��_P;��)S!��C��`Of�'RҌ �[��A�������R�7���o�%h����;���(� �CC��EJ�Q[��������cC�CI���Q�>�9Ί�ۑ��AB�)�VI^�I��^k-�{�rwd�&Z���N�!�Fk���k>�S�8Itk�a��^M16+ �3��y�)�_pll�^���|	�~����|Pt�Zǧ.˦�Kz\:7������^��-����r�jZ3/�����G��,����� �ٌ�d�I1�n	�����I����#i�W_�M�h��+�I�����:ɛ5�BϾ)�2�B7�Gt4O��7�h�W��8{>j���"�<2.�(�
�1�gS�:u9��芷T��*��m�Z�v$�|s��'�.k*�Ⱦ�}̝�ф;��@e�/"�Z���_���+zoY2���	�a}p���B�2zw0^K�/,Ղ�k�!Xì���#�4���^��Rj��z5+�U�B���lpd�@$�ȹ8H"$��T`T��1L?�V��*x�o�]av����r%Ԋ>�pI��xn�SI��8�p�-���F>���zǌf-\���u��o<'hN+og��U��������33��)m��-99��G{p'ci'~~��n���H��9�tÉ݃��?���/q�z�VB�xd|��[�ÃS���s��2neh �c<��"�\gT|��-��%�-TV>� A�$���6������h�P�X��i�,��8����3���b���e���Fѓ�T��4�I�{e��M2��_��૏􃤶���*ُ`e~/�^q��')9Q����Ц�X����ք �In�5ĔI�h��bm �>�!�F3j���������6 T��`'{"8��XAHJ��� ����
��i�s!�0ܣ�n�|��+��F~J��d�y�rc�ySh�U��*�P�1�������9�#�Kf���R�ז�0�u�l���k�� �1�7)Ly����t��+0�0趱�K��LP�1G��q]�S�"�X�[��y)��lEz�?�yKp�E���fAυ](C:��<ڂO`[�V���d��7���K�ӹ�a�uo�`�o��sD�$@TU�v��G�iLu]X��kg���e
/o�p����O)i}���'��H__SnMΞ�=����T�����p,�n�&B+��<�Hl�]j�[n�\���]�|ju�N��HG�
-g��AZ��[�0����c��d������Oa߈��.�����D�0�">�Lc�Ë���b��ѕ�E�������9��Q��:yK�PO�J�A.��4�����3.>po�vr���m"ST��A�\S��e9I�`cr3
�����X<@Sfy<DC�Ӑu�ҵT�!�@H��`��l�z�A��D�b�!�[�i+���v�����w(]�����y5+)mH�}�B3��q�T�kGL��tP�4}�y����i�	����X>/�J�U���DO�6D�~o��W���1P���� �o/V�e+0��5�1��$y7U�~[����Zs�SD��Y��3Y�08B�� ퟧ��wq�]���F����Z��HU��K<h	I'��r{�E��V��=+D	%"���������1�A��G�AS3�kYFk���F�bRQt�%�R���		s V�T�o����ۂOι؋1l�j����s������jC�NS�b2��\� �~q$�w�/%yk��3{g�ܒ�p1�&���U?��y�>�1�\���d�o*�y]����;�0��G�,x-�0+8;@<�'	>ȩG������0~ܴ�^Z�\��('�ʨ��ЕRqL�[3�Qq�n/Ün�}��U��Оa��({A)�ĭc�bj�u�
�I\c�2E�5#�v�aO̹�j\W�/㲹��Q8��Yڈw(�QG)H��{م�������m}zsm'vX���H1H���
R�5	T��o�[�W�-�Uo~J�m��*�����װ��h!,V7��u�y��(+ʴh]P�s�8��P��s#���L�c/^�pE�3�O�(Į��9R��)��S�x^$I)���dnw�+:���%\�0�j�fзY���
Z�Y���\F�E@w�(��@埞^Z���E�Kʓ�T20�����CL��]j��z+������n��y}��B0�Z(�?�5��1��cݒ;�p�qm��9������َ*�ݪ��7���y�\-;�)�]{��B�j�)0Nhb�D>�=��E�	g���6��~b!�0������u(�'l��ɝP�F@��H�V����.8�����	���4Qu�]��ӆ&������Xbk�������?���-�V��8N�g����9��h�έR��������]W
;���$�] �)|��g ՙ�3<�������H�V����~�<�%�����34G�\9N�*�8�!SM��p8��/i�Qw�����L?���ZS�,�roAo��.�eT�4p?�C��b�&���[�뷊���_S'�"
�e�l��-`RqDB�����v��^p�?a>��{��/e�K��O������;��
��Ť����AN�@�6an�V�_E`a��=�1
�ޜ\4�L6$��@_�{:���lwP[J���Z��y��<0�K� p����O�@#��H
��}�N���&�ڱ{K{xU��1��w��5��+��l9#��������/_�]
-H=l}t��ú�*� �G'&�@�@�)H��^x�ʚ[��ɱ��;�k�6��W�
�%�,O�_�tmv�[�<֙\����0�Gp�\z_Sgq��a�fϴ?�������2��ʸ�/95[Gl�Ur0Q����8��"(sM��;n����ln����U���kj���aSe���q�7�������h����1�R�B�_H��U��Ž>{�1I��LF���]��Ӭ����hC�p���FX�fK��@C���y�{�Α�Ƴ\�ݡ�r�I���3�H$���1�a"�5���O1��r���3�iY��H��H�����|�ڠ�ح��tA}E�����������qf�s�����4�l	�8�i��x�u�J�J����T��n(G���s ʟ����CR��3�Q������ �C��+_�lLw��%�/�ø�2����	�Λ�E�+������/ue`�� �-�$��Zm��`w�{�$�no���)hE�w������H���eM9�J,40��寅�F&F@���^g�K�S&ƨ��G��*�քPJ�,�䌻-��@���L�������m�����"��¬0/��K�Uum���&YN�S!��yO�ܫ���X����_��L�rX�v�������sz�X��\C���Cb����N���Dm�r��^X�<�ۓ��_�˴|mH#�-�&�a���M��H�J<I� h�7yN�W�O��`ӗ�{�@(��$ۤ���	�X[ �#=U\w���x��
m���4����R�&ȫX��%'d���c�w�ల�q>@����j�����!���=r��V�yMt38��W�E��rb���>+�Y&��0K��,]���4�ݓ.Oo��Y�/J��v���k�Z�g;o�ĔL	�_G�h;�mi��U�s\�K�{Z�n�O�|�~s��IӞ��V�>��3|��T���~��"�ً�.��q�A��i��~I �t���F,�gQfx֥UV�`'+a�.MV���z��|���en�S`������4�!�i�	w���
���$�KD՘J,B�f����L��cQ�N�u���v�u_t��/A��S�����n&��y�w��-.�U0Of�ߔd6��|��JQ�rc�o��U(wS�^c���������S^��2�#,�n�ڎ��W�!{���}Fo�S�%N��M�gA�":��AL��wmH6;�F�����`�a��T=뮄0,��d����OaOa�Fk@�=9�U�&~��5n�N� ��և@�3�[=G��)S���4�0SO�z�]���I��	e� ~պ�Z##�k���!�����=cS��lѢԢ��������,Qm�#��D�2�q��F��I�p��Hq�ɳ��t��;.�O�7ٻ����u�Ç��et�� $�_�X̒^'���$�9y:������o�C�Z��/�����.��r�#)�w���D.G��g�!di0<-�<*�����nQ)ϧ��w��|G��\Z��Q�W�lu��4K"�tyJ�
���}���FsE|{�=�<_Q�H��9��xX#��}���	�������<b/�G� �b~��)A��4 ����3��>]��|p��1RG\��~�D T{î�<]�I��T�zG���-%0����|� �?�RQ�F�+V�9��o�)��DEl߱�GZNm�r\d&R+xR��9��������\|�~�� ��:uӻ�X��С�����)������d	�H�$��
t���u�i!�s-f	
�ҩ�L��݀�mp]��U09˗/b͕��N���_{ݑ}
Ȅ��M���?�t�&sa�r�M�����X�Ye��n^W��d4��%V>���l�A���� 5^W�.�h�F��p�?����n��|�Q��)s�mIu�|}/�v�c�8���B7��lc�b�+%5�,���o��@ h\Vt%ZI ���h3f��N��q��E�[t��Ǻ�B$̔�9��{���y�WR_dAG����� ��V@�(C�{@*�T��lǒ��:F��8]E6�^����Dg�����vl^lA�i?�C�s;����*����u!��eO%"M�!�t7}�l�m��p8!������s�*E��%���+�A��9V{$a)P4l-"/���ӎ'^�A�j�Cm�4�,�9�����h����l��0�֙�F=;��nyl�^i.!Lh(?C1GUo ��W!�f�H��a*��ndg�HC��{Y���o�}�l!��d��6祤�\���U!��C�Y�����PVtdO�b�}�h�J��|�H��b_�a]�Q|��6��P��pׂ�n�=	R��V;]rj^�
F��p8�(Z��1�A����X%�Q5e��FoG���̅�C�
Tq��Q�����M�[�t��i��i�$ﯙ��@�����K����k���4�KP�ث���o�}�/Б7�t:�'��v̰�O|OY��*#��ڭX(3gQ6K�&K!_T�״�q�v��,V��1��z�Ӥn}3e�1��G�-�Y�����A!����!]rJ�'�8�����@���F��� #��O$�&o�ƣJaU�d+1}
8��¥i2�̣��� �Hm?�M5����M��� �a�����xER����}H"ֈ�xz;h�6wR��l�O[)?m �@M{�($��4�2������"�e%�r��h��|����u��$�j�����Zq_S��m��,���Z�<8�A�q�(/���m�#��*�(N����Wk(.:oA��(�O����o���N�
{�9]��{v�8پA�6�d�������RV�LK��e����V�\O*f�T����D�㘛EU$�<T�&o�����.`�(K����п�K�Z�z����M����ѥz�_C��ٌ�*4l2��CJ����_���m��*�XZ�z>E�^Vo>��u�8�p��H�t�~������˨0��TUuㄤ/�xv��-�>x�s(��b�À=R���lu7��m����Z�3m�D��d�Ӯ�	��\)>*nx���P��5#G1�k��٬� �/[�=W��H�]9뗘�!��a��p��㧣LH}���k�in/�F�,:�U!��B�t���hpBv��������K�)_�3��c\��:E.6�R_R.�mP�T�����#�/\��%���LG%��Ez�Y̓_���ϑz�Z��N�E���Z�t���*�"�P2ʩx�n��Eȴ����A$wYA�Eb#50d��*Ь�:�h�f�u�����i��Q31��Z�M ���a��Nw�LL���+e�@�l���]p<1{L���v��]BW��^�	��u@��7,���zBUa��;�> ��4�3��?q��yއ���hQ������g�)=�֠G�W�, E�1�a�;HAMm��U)V-��N��-&�d���?����}\RnJ\T�h��n'u�(`]:H$3�*�zcS��9l���ܲF�vo�����P���������VF^,�r(��H�ڡ��w�vF�؆��~5 䝋�ࢂ�&��nbq�L�F� !=�nb���	�Ҵe��=GT�9��2WrK������k�Tn��(�F�G��2�e�z�?SD�l��X*B�0`�e����_��OÉol\9�Uj�C{�� �J��m����D�k� ����=�|���"�^��u�X�|���/�b��G���=�V�-m��qN�?k�� }��I��v80�eqC"$e=j����ҫ<6(;����������]���Ϟ,e'��I{H��F9�䣍 ��L
�c�(�2��E��S3&�����SS��y=^���:>V���}��Z�p�F�J��*1>�|sj��W) P�ȹރ���K�+�;n>��P���B�_��l�X­�5����"�rMKf`�m��X��Z(hI� ��ZRzS���o�-;;�c�i���#��
_ϲ6���c��E�H�X�q�9��a,��6g����[�/P~�G<	�ñ�M���Ǟ�ɾ6f�Y�#�*�
��b�|PC�$&!@��~��	]\L�Ct1��C%	�P�2�})u+�(}N�S�l��j����bW�aA��W*AqL���Y,O�t�.�Hߕ�iG�����o|Z�J�������7�<4�`��)Gu��.&�z���
�����-;�~-�$,�TO��(z&���z?L��z�@z,��TMnLTuv5�2/R+%i�,ݦ���9�bd��aC>��>S5ʼَZVl؄=Ќ���JN�-={E���̼Žq_���qRe��;��<���'�C�nc9�K�����ɴ��N_7}�-��4�#2���`Ca�jk�]I/����Q�`�������r��V����c�=�???��x\���7N9{6ԮJK�z1q*����*�	2D�*:M��sʩ}^�!�x�_[GT�ن�8�I`�M�C�	8����v�-�r��x/Oy��`�Ӆ�sX�����B��G/���.���/�WQ�Z�zy����%{s�~oz)F��#]�N`��������]G��3��i��\��US�2���X�V���cΥj��3��Q��l�Q ��4�÷#t��ɪ���x(���S�-�9���@��f1 ע�F�		�"���4�J���'r��R�D�ā�Ћ��u��>���Qd��G���cz.����R��UP��f������������km8]��s�@����9I�4�o���75zqz�u�O����Tq���ZPT���)�%��ؕ�u��zň�s;Тqj�ꀀgAZG��,�Z�mJ �zl��q���1�	��wF��C-3�9("AS2���0͋�&tR)�%����-`Ph�G�V�Y#�m<���Xt�!v�+6���C�Y�������p�Hj+s�6��Џ�N�^_*�+����7�B�䶪�3��'�J����}y�xDq.�>�L���V���C�V$<�֦�k,�Y�zW��������s�Z)b�?���F�Y�Ea"�.��
����cg�Qۥm��KiW��w�*�[k���]� ^j'�n$�x���q����] �45��'|_�s0P{/�}Ӈ(v;���5��XQ�{1S�s0~�M�(U*a�짰]�8�(�~�����C ��2��+1��c�["�/�$��*%ne�����x΅�,�FX�x�)Ģ ��=���9��ȩ�=�5!���
+��>}�܆��sT�[��F�\���xF�lha#�-��������|����w\`�sK�)�^[N���$��<�esSK���!U��:����-zI�F�����mZ�v�H�����?�.�Ҷ�V��|���GUǋEܔ{���_a0%sY֍Iñ���k�h8�x���5�5�s������!����2=��ĳý�ѯ1\������e�+��5����(��#���?F[o���,��]�hQ����^Ĵ���}>Z1��~U�r|r�W�C��a�$��4D>��y�5h�3/��鰄��hӱ�1f|�z�}����]zF]�|��Z�Z3� �zG7�`N��p I6�� ��g�<�:�?{Z�AŨ�V��Q����]�F�F�xi%��s0���J����R����4��q����j����'x�մ��y��S�:��S����O*&p׎��Ͻ��S��XI�sm*�L�қ�b�X��S5��C��_Zee������ T�OW����#4*����8(z�T9�ɠb�����Ɋ�t��W�<�s�P�太�U�|;��qe?�{���Ln-�}?�'�[!�SV���7�"]�(流��n�J?>���������,|ƥ���vm ��Jw&�J_�BIu��QB+!/�8��G~��I�u@1���	��q�Pk6��y��g{t�/ ��S��6>�2���nv0��Ѿ�<���"V���x�Q���*�F�A(W���T�9�D���� ~ؠ�8�f���i���#���ff��~s�K�@"�B��N������gYAt���b�Ǯ��)$A������!7bL<�B��%�M[�c�X�_�S���7�u�-�Q���ԿN[�RW��}.#
-,�K2i�z��^u�g�f���j��^-ǿ�
�]�I���Tıj�OJA��4�q����
y��g��[��	|&zu��$(s�ꑓA|h��/6��6h��ڻ�������I�'��y�N�2�9�a��4��=}~P����h&uk��]���
�O{�É���3po�ԗ{]^g�8k�[���{�e��'7��F�Ylƺ������?5E�W�б���tL[��S���Z�0�:�����S���n���q$X��<Ӣ+c[B�D/A�C��W߾^O������.?8�C��h��}����U��0�Y�Q���-`���C��R�o�7�g.Ώ�=P�wB�m0�+�^���ۮ�as`����R��4�I1�g}T�w\�PmҎk/�g�������a&Մt���I*�O�L�m�=��`�����6��"�(D���r,k��C��j�����	���(�p�i^��bpHx�
������3'��"�eWp��I���D+�gu�֫1u@�}�1��5>/j[��z��7:>��R�n��i�j�s�W�&��AEx��\����|9>s�(a?BY���{6Hr'p�ڃ�p���nd6����.+�u� JK���d�#��������J�`���[�1
p��w	�ļ���>��
�r�$+�?�9I��k3iY� 6І�	\{4��H�у�䠠�=W���ہ����/��&/8��M�4a1�xl�Ÿ9�`c6��ţG�y�6�Lg#�z�{+���~i�腍i�JP��f�d���\M����6��e�/���^��2�[�K��g|M�� �����Y����8��fڅ��i����m�	7_��KuZ�A�����B�-�P��g~,x��[@6nݼ��!Ky�I�h;ᨚ��Lfn�awlQ����G��,m��K�����?� �W[�]x�RvIô���:`6]>��E�M:���{��}�<w|�`�/�����Vp���%�����&�M�����\C~��>�����}�,ہ�el�7������J�'�;k�2Uo�1����f��,]~9*���~DX�m?�|P�z
�rH�72���=�M���eG�0�²�π��K�%H78a�����|Bf�������4A��m��w:i��Pl7g��)Z��6VpY�0���6�49��lmȼrS�÷sq�u.�pMő�_>�H(�au-�f���aN��L:���U@�� �Z�
���In���
�Ϡ$�|��>W���(���9VS�2n�9o��Ӈ��Uy�a~_%%PѷzE�
�Y�pE�T|̾Z���Z�g��՚Z��"8�㌍��&M����!��]&gT�Z��,���k��m�`?1��rU1�0J�A�-q�3������[��y^����e���ʎû���|��I�r�8=�4N
�����2Y�3p��ܛ����������
�^ ��E�0�����J�S|�;�������|���_��^��񮍫�{�羭Es���o4\cS��r�p�����d��n+ +���w.��kK2�c�VP�:�A���W<	�/.���*�'�0�1����8��������OP�����Oo�m�:��Ȃ�H+�9�i�aw���;L}��28�2o�B�<ټ���@�$P��Z�Y�g��f���y���UQ��A�ƾ���_N^�l�စ_�%̣�
����+��㺦�WŇi��Չ$D���<.e @
�b�òGF�ϗ^���2�^�?��ג��l(f�%hͷg�6�t�=� �L�?�	y[�|n��\������PG��Vھd�Cv�'�5�TQ�m^��_��
�U0$:���c�5Ŧ�����E��o��^�E0oY#�ే�Nv���F���`"���H/"��?G}`� �)�������IOe|�����6���?��m�k�[GG��-���[��+�PS?g�CN ��h��ۗ3�P���M:KG���}}�7�8�K�|���g8��|q��o��WAC5�v��K%���zƓ�v���5���r�����U�e�o�ܰ	Ƌ�[�
�^��8���q������S��#����g
q�핊殗��sy�)]'��57�s�E���{uQ��3�]~-�;E`�u�_��z�d�SJ��r�
%�Z֌��f�k�Ri ��)X;+v6�~�RU��ؑ^����0'9,�����?=�]w|N��\ h����.�N��r��u�[\��O��4��Զ��`W:���9����܂��
g؛�ѳ��s84�Ts�~�\��Ӓ/�����������1.d$��nd����!m�>���h��p"�f��QGy��r���$ݖIԿ�������]kǖ�.]c��h�»�T1o�w7־�.��c��r��G�o�U�=�%�x$���
)QDuE1a�EJi�{���w�J�uܐ�f~�S*U���H�ڈ*���Jq��9�%[�m�ԥp+��������bh�o+��Ύ��W����e��JƘ����.E��Qz�'�L�L�MDS�u8�ӎ|���!��?�������y����:���%�]�Z����ӵ�-�R&�L=�N��O+iQ4j�{\�N-+VV&{�0P�c?"�*A? ���<�(C���G0�>:�k3�ү}�>>SJYֻ����^5)êϺ�N�����Y&�90a��
�W�\�1NC��-����d(�;���G��������-$��ն�2'��}�]n����+t[��l��IT�=�&��'ώQ��d1�c6��W����]���Ӹ���B��iɦ�oO�Ry"T����T��4�(�k��.,�;���z�zY��M:�[�4��_�����k��~GI�Z�斜јbqq~�g��5�Us7�LƣU��]�/�ƕ��ˬ�KdAQd7�L��+SfBZ7�i��~��<�A�]���\x�n��F��<=w��A~X�V�ͩ"ܽ=aO\B�	���-��w$��z݀��e���������#Oe1�M�a3�`j@᪹��{*��m��3����?�	4�!S� a����/��i����>�(C���XUI�T�a�z�7���7�Z�w��a�z�j5��6R%�"�?n��8��NEA�V�뺰ڞ�`a�K}!i��􋜵Z
���~��jg��O�����#�"�'հ���E����vc�M$4_�J�	l�-�'�R��u��d��x���ŕ�GA�J��7��^+#�r�[D��C$�qhuZ���I�7�'tRX��P6@O����]��[�:<�\��w_$N=s2�9�۝����=�-q7�	�;�Z]_0���y~�卅#�bG���)��وa�����}\�P��:�.X���0r�?w�>u��kz�|*搤�D<���Y_�+b�y��D�X�D`ŉ��w�3I�S�X��y'�׫�fတ@�g��X�B���Wȫ�Cp�ysW�;-��F�yq�Xcũ��w�nV���p�s�h�o��<R{�ӁTE�Ҽ@�����f[>wF+nA�G�5��r�9���IZ/Xڟ���`[�Q�ν�K�:S�u����, �8YY��>J���S(MCEv+Ko2S�7��o�DFx(I��}{���ٕ����)렎'c���5�����.������\Ō�<�m�k�*�P�7��U�p����%�A�K���I/7Np9?X���z�䡓R���	J����C�a�&�Rw�,��?�X�iq�U�լu�4��'AAZ}�Ӹ4%��òd����hK�E;�S�_f6���.
0K�Or}h�+9����z'���(�˦�T̬�� �e|�w�#]d�+��&� ����E6��'+vw��aHT�@2�0�"_A�I9��(}��t�4I?1�K�R?�f/5E�SJ(�{^%0���_P�RG5����
��~��E��Ub������-�mNA�|!��&\c�tyH(��/���x"Q=Y��)%��R��F��]n>��؏��*�[7� |��Tv�(z!Pf2�V�jµg�k\:��+�1T4TWޔ|���K��]�9~6���}`�>��i��q�%7����c&�u���3O>��k=�\\z����Z��ɫRs0�\����@��)�����:��G����=�o��7(91a�x�WJR߈9�s���'�K��	g��=�z�&��|"��{�荊I����	E��ľ�[Ĭb��<>� �otL��I�����}+��W�m�����������c��3��ٟ,B�i��M)�/u+s�<BE����V8�x�񝤑�������!���4r��`�K|+N#$�'}�ȹw&�V��v�+�c�ׄb�%�.�]vĮ{)����WX��x���+��SM,�D;�(�-$%��ƙHԳ�&0F��ľ�(��Λ��T<~���xH�=AK�>��N�q�����8���j��'?o���R}��x��}�eU��z&����&v�Ҍ5>����ErV��(��c���D�S��r�}�7!d���bp���H��B[6u��QV�7���_o�OtF�l�a_�[�(H&L�$��p�N�E:8*�`F�Hl/�)���g��FX��Bg�7ն�X���E�������=�V���ׯl	1���d��ɿ�$��b5&n{��FJ2����8|ߗ�@%��@g!]QW�+�I3���-B1��?�/.ኘ ��V�t��1)�~.���%�!!����J/^J?G~��iY�6fQ��uH����ƚ'����v��n'�wDM��ܠ�ͣI��^30v�l��q��������!�_z���zRN�"Z��g:�\,Ә��}�=��q�hNP/�F�'6i�����ij9���5�e����>z>�1�XWq];�������SM��[���6��I<8T�t
g�4.�5��Ab�W�w�R���:⚧����h����JҁP&��x9���و�?�.6�~	�٧q��ua9�yA�(�$I?JJ�����1�kj,~��?�� �"���S�4 �ﱱ�(<��hZ{� k�ƙW}����"%��q��i�m���b�4 45Tr��v=DTSa\��ٺ[��|��/'��~1(�=��9>$�@���J�rR5#8��}c����e)i�ב�2K� 0c�B���<tfq�*[\�����@Ef��,N��j��8��u�[��1FA��f8��dO7ȸ�ʁ�l�M�(�:�?D�2�	�&v�y�84�+���'�5���kH�	ޗ�����{p�ĭp�0s�ѯ�2,��eY�V����M����}-W%�!�%�:�x1ȓ��7D|�}i8�de!�c��5�Ȑ���
8s{O�Nń<%=l�	�[���Q���!CV��������-�>�z�ſg�Z1MG��U�*���Ì5��:��<�!�M�`dm���Njc�q�%���Hn��$R��W��6���h��S{S��2���{�ƭ�ڐs#���������K��"&;'��%W�|�&,�2}���x(�
�.Ks����AWx��t�������H��	^�FR�%�� O���yxz�7v���8�!sO-͢eRP`-�"���ĩ8�*/�!�Q�h����Zq�X���͠RJ�;xCv�M��p���o���A��SF�9���z�Y�������]��� ����}?�y�|�x�W��݂_�^���4��yH*�8��z��}���W��;>�ϖ���?�م�����/U�+�f��T�r�)h��wRv��M����|[��:�^D�F�у\���(��H��i�lj����P������w�g?�n��p3��q�? O[9?�Ē��B���#8ڎ):�S\�f�iX���L�^t�A�����Q
�6(���ߗΟ*?W�������yS}��%.�]҃l=��kPZ���Ñ��(I7�֮�6V����$� �ոɞ"}H8_���I�+J��C���5h�Ε�U��X��cm1'��N6$,��h���X~�]#)���v)��UİD�&I�hs3j�]q��l��=�E�*�$3���jGbV�(a>��2X���r��0������J��2Z���f����N�Pk IP~����e,+pר�
�t�u�yr�����U��/��}���ݛEg�Rp��4��E�ų�U���h�L�iey�4+�MP�����W����Ϡ�s�k�i��]�����#��%�VWюP1���v�mlX�W$�L�d��x���d9���N*9��v]M�h����&�
e�62���\�+�=I�l@u�p�<�+�䀝�Ն�Tꏈ|
�4J�0 �%�^�_|��&�&�*�z+9��3p�o�W���%
��(�m�	x>�� ����������{'�/
���6y���M2a⥙]����ع�,�[ �.cQ;�a���x3�^���[8F�&=��I�y�ͦ�Zr��
j�ĖV�&4	�[x��f�<s���:�u~Z9T�=꧎�HKaT � �0���s�f�������8��@G��\*Ag�7��� s^o�Gi� xv�c�Bh���4�� �m���g<���"M��q0^��G��m�=�O����D	N ���=ޡf*|����=E�d0/3fN���H�������RI��U��"h���h���W��4+[K��A��B]VY���9F<���[�u�/�}(Ag_�(?�D������6$��O��dw&�H��ƺX��U��b:īlX�	A�k	EbL���e��G~�$6{�&oK�ˉ�s���o����4!Os t�A럏KP2�+��6_usk�)�Ŏ��\�q�Y♱R�?lO��L�Z��n�����6 [�q�G/��#/�2/1��� �	 Y�s��A���^�6p�u��-�K��W������
�3���vs
��<���$2EʻE K��y�s�5�zoi��	9j{4�H�������/WN��uc�lr�o�C#`	��I��ܻ��	�"�K���p2�ł�<�����(y�������UG"rj�v�][��ڤȡo�28l8J����y!��ң+����Ճ��p3t �FF�u:.���j���΁`u�q�@��rH�!/S��v0&�!+��;��w00���[X���q5�n�}� ԯ�U2�g%DvɄj���<ϑ߇�4,&�T�T^;8��
C��
��R[p��U%*�s��@���Vh�3�.����Y��k9� T����p1�����^5@\Of6�����p�I.���B%��+_�����)��2�w�Ob�8U"?���8�c�*T6;�Մ$H;P�9K������T5ߡ�Y�'=:Oȑ8��h(�h������[쯲ɨ�$^ܐ ��Lׁ��0i>��u:�2БA�P��+�@��}i]��a�d#�xS�ΐ�ʳs:E��9����x�\X����!�^�N���f7��0��Ȭӎ�)xp�vc2���[E.T��g��|����RM��_% [ݻ��<x^cy��Q>���߻��Vt�:������U�E�7�Yo�h�h�i!�nc~���8�1���%������/%�s�=&C����-l>,z_MЖ���l���bS=�l��P���g��7����I��0-e���"��$��m�vD�L��>��W�C���s���)Rb^�=���é�^�J�� "؊os�?xE�?L�J�X_X�_��L��B�p��:��k�E2t'�;�K��Ut��As/|���|�"��s�&�JBE���D��e����Q�����z�]���G������x��v�Cj�!��;ƌ�0S<��}w����u��9�}k���O9��`����-Y��2�4�B�[|ފ�I7f{���]0ݙ��n�F��TG�������a?�r�����tN�T�b�4(/���bb?$�W���#0S��)K������=�+i�W�0��zCa�+��0x<������g�
Q/:륦��n��ڏ�B��u��)���H�k	*�߹�1�9iT��e��O>*�5��tR��\07p ��-�ww����h��q�\�>����m���G#m� њ�7�F�@�Q
��0�˞�02�P%���|�,�7 O�գ��R�;�& �Οm���!�w&I�[�
�1l?ȵ+��A�OU�}���0��k��&�CH�s��d'F���u.�;%�Ib���i�c��H�.ȹ�:�!�y���핉�ڽC3��K/s��94�s{�G`P�G
�E�n	�����ݜŒ5���a�V�Y���� xۥj�gIKƾ �S�;kE������f`�,�u꨾�Ȋ�tS�x�9W�j���F����Ճ	�"KHJn�x��"��؟l��b��`E�F�����T�0�ӷ��U١@[�t.4�R>�R��6�g	��_x���K#����jy�$� �Z���9�A>������h-^�@����)McЏ3��E���_w�� � ��替�9 m��;3��0ń�~��Kkk�1�%���m��]E;&����(Y������n�>�B�w���6�v�r����K� b�(IM����"z�jƠ���v����["�m�����f>H���,2,��ȴ�D]���]�]/���ZB�a\��t"�H7���)Q��3��y�c@B�}4XIǶ����z&h���x�>��l<z�8�mG���R��'�Ƒ�d=����0z,o�����:�/
X߆�ܶ�7V;���C��n���]14�����H�P�wu�0�6AV\ɯ{ڊ��E�q�=Ӯ��u�9!�d�Ar�8�����m�GuX��mφ��*+���3eRdI��ι``�Y�������������E1J]���o$��3/�L�����e]*�Y��	}�1zw�_eMq�x��tە2�o�e̅^���l��qI�-�&���Y��`C�'@.%g�0�	�G���yC"�G�S_Vì�������Cx���DD6�̹,o�Q�^�>�ͩ�Lgb8~�x�{_dh,z0�s�-��O��3o `C����(��8	3�?�tEϝ��<t�i��KAWP�ȎC�ˣ�.��ֿ�3߱��F� Y�:O�9��l��G �8����3�w��wy�IGA���t�J�+n����Mn�� �S�f����yq�ڙ�"m��"����E��D��a�w9�k�)���=�s��y�S~;b%f�f��rP4ʦ�Ȓ���ޔ_���ߖ����2u_�c�>D�pD\@�\�N�<��J.j�̹�H�8�wn7Su��8+Y�q%�G�I}Ll2�WV2��iۯY�?1 dHë�F7��|�8�!��*�4�?Ou��9f ����%�p������9��w5�pX�|���??�R��zh	}*3�C��Wď/* a]�&����;��c���w|PT�!��0���W����柸�F0��M�b�S�"��˅��3�L�Wvg~��I=���E�^��r��ڲi���]��!�\����4��٘�ن�Kr�ü��}W��x҃�3֑���đՊ;%5�q��7Z7i�6�q3*���w2s��<�Q+ȹ�B"M�έP�5%RΚp'�!��4/�Mr�Y���r�]�6Z^*���粃(��Lt� �AQs�H�
 ʹ#|c�'0ɽ1 u>T��E�Z����гʠ��\�JJh�.�q)h��ގQ�����@B�^��ߣG��")�N���9)��T��Ҁ)�����A,9z�(")趇��4�m��yV)U簾C_%�me4�����`��A�4K88�\R҅�S�u�2��)���IBPX*J�I�X�#X�X1�)�H�W��OX>8F� o�S ��a��M���^]�����M;q����6�D&�V:ВE����~�ǹaL�.�L}B_�������RGH���_�%zdz�� A]����Ҋz�����ͼ��/M$
k�<-o��Ueӓ�1�y�����y�ds0��w�1���}XpN����[u�Z^�[gn������:�"��U�:]g��k���4�uP���I
��<u���E���Ë�0ǘ��<�.��Y$i��h�����H�;>���������������]�/�����:�!��ԁLdޯ�~Q:�
(���iEXD�o�i�v9���.�+���i4��Jژ���;��#
��xs[֦�ɬ��q.?��΋<������ڑ�"�"��_FRUֈr����<�4����I�ݡ�tQ#�E��q���h���|����_�Ԓ�=a�iS������$���0�hh�cͳ�q�+��և�����y��(��$,�D��h���]��V[߰%�܆H����fv�JL�b�V��J���϶P����\}m��H�D\���]Je���+5��%.��s���`A��jz�:tGP�;�#�'@;Ѣq&n�M���� ?�"d�u�o:����n �~�S�5`br>{���z�)�\�V��4w�l���#��6��� �x̠i�RR���Ҽ �|v���tf�s;600����ys%>���ԡ!���.@�s�l���2]�拙�>���4g}cJ/j��Vj�˯p����%U#	�H|�Q��t���� 7���nԸڕ���/v��ꢀCm�i��(?Y��]5��H%K����q�X{q�V���4�q]E`��0wn?Ϲ�y�mz� 1�_�9i��d���[��%~��zF2�2:��~7��]�g`
�0��F�K,#Mp�*g<;��̶-���9�K�t&�o�f/IĸҸ�8�u�F4	��3�q{D0��m�N4(���W���}S.�'DgR;ލ�:0�,�k8�nFL������n�h����"o���l~��m���r7���~�����|S]!ͦ�B�6?����`QskiۗZ��b�r��o�"��/��R3�O�$����,Q}�4-n�i��s����2#I�%�h�����4:���CA͋T�� �\�hc:ͳM\�G��	~��"����}:��Ѵ��њ'1�+p��i U��$�.u߯	��D�A���Uб��a�{R�7X.���t�0�����){,��;�o�%����0�n���J�C��l��*�6t%/Z��)O���B�]�*���G0��~~S�S�ݖ�{�Ric���rt��K�%B��ja��a	E�&�=��B�W7r�Z�x ?b�ݾh���ٳAP��*{���I�M|Ji�(;s�om�3���h���z:��L�����_��ta�w��ӿ�N7���T?{��q�{X��o�����t�����$<��=
�tb��=d�	����D�Fݛ����<���$�{	b�H�zug�R^�y;��C�|�RR,o�N�	����	���$ ��n�ޑ�����n�c�ƾs`4Ջ3Sj"�_�=��"��s��^_o4�h���с"ho��/�c�{B֖Rm#����l����%^�#��!�����d#�k1�)C%�Z�GҲ-�lf���N<�7�=�5��-���呑d����̭��(�x�K�(k�����I}n���*���-�C��Đ'�}�����P�%�`�<���w ^�M�_ �m��-+���V���
��z���F.}�N.��#+����y��գ�v7q�xҢ�ۘ\��|��~;9�f��9�Z���u�3	���3�x��^ws�F{f��c��*{\S<
=�{hHr+���\Ҧ����3&��l�����
)`c� ��X�C�B)/A9�BGL1���U��@����s����8ȶE]��a�Z�)���v��T�v%r�*>�rݷqj�f�s�DR��>�=V\��yfM�u���:���?r��6^��Sc���n�yI2b��:�v�	��E����cm�F0T,$�9��Nbmf���<�O��Dd,�P[ߦ����1��ۥ;;�[��Sd�.�}37W��:�A�[��s*hzH� yV�r7��s�\p�'��q��"�
`�7��
�5�x�@t}�5������{�Xz�L �u�mALz�!��W<�['��4#a��-H9#뛫����Rq8D<&�K��p,ھz�W���e�����g���if���7T3&J���$X�|DH�6�����p�+yj�
��D�Qv���5�\�����=ۯ�H�W����6p/]�Sc�|���i������.���)�z��x�!B���ܟ��>��$m����T�J)�'�Y������8'�X ��B�Ym�@o��{�Q���C�F�B�	L�\���oV~=ŔXx& �mg�*�@�EtY\W��h�z���PbF0a@H3����#KN�, EyL��|&w�^��خ��/���B�������cѸͼ0�g֖w�4�� � ���	�?6��5�a1S��c�X�LHV�uz��-L4��bS_8I4�1����2t����,ɃB�W/Ws
��`J'x�f�W��Q�����{� /���O�����q0�|ό�Sw�w-���0H˞Oh+���t���>���W�� �:�����\��/���HK0��`�څ�$��q��YL�)�I��AԮ
�Sa��`�cӬT�U?�1�ͅ[�"�pnW����}�Re9�c�ʁ��0����Ybr�h&]���%� �D&j�\ڹǈH���u
��7^��<ۨ�k#��7�Z�Z8хz�"d�6�E��T�p����SHgQ���˽nc�K��M������E�u?�m�Q.��M-p��w��^Xg���g���4�o�<�:�#���!��ϑ�D�P������,]t�v�",+5�R��l�SD�IK(���)`�#{!�P��iX	�lW�Z_ؤ���Y�#�KO��$��Gi�X0��v�*d�`���Urx��imf;��,�J�p�$>JW$�L��&x�h�M����-����qB�T�Ac�/�I(�E���3�<�]��ÎⰝ9&����\qqηܫ�*�Y ���1]'��o6@�T3�����wxG�圓�r�3�|~;��4)jP���ӓ�/yp��VR�1��%��w����\�,e@*��P��7t��(� ��:P�J�Rcw΂X����7�(Xs�aw�r�8$/Z�����f�W��`v�9��-˓��v��)q���G�)�6,����w��Q?��, )ե`-v�;����PA���G�
3�_MA���@�߉Z_\]��w �Ðv�'.���߂�
ޚ���獶96�,��rTbpAsp��k�&8��@+y��[f{�m�� �ӷ��L���k�M0_�g��vUF��Ν�ae���������mZ�5�����g�)ZF�0/D&'=x;�}�g�O�u\�U���
��ʹ�< ���,��d؟Lݨ��}|ϲ�-A��W0�^����p����q�6��)a퉬�	í�������u�ew�;��L;�6���q�� �)�y���]:H�XE���>�_�eZ�K�5��u�J�@i�4�k�p�K�Ț����n�7���0�u������9��YDVO��f��bt�x��.�&�/���On�+>���y�h��kYs�GjH
0�*�p!V�/������%�)5*����=tu�P��6�"�Ci<���+��Sog�$q�7���J�gBSqlabTac+��Ӌ��ŝGa���_nf�uֺ}�n��w�bP9�\�̠y(3� ���X'��%��k�YǑ\9>�Cڝ�2���k�y-������Č|�#_��g�7�./���:V��̀�H��&���IIƠ�Q+5C�p39�$�u��$3���1�\�-Cu�z����VV-lz���X����:�~/V�?K��ʬ�Ä�7�wZ�{{u�}�l���;C?��Z����-M�I����15�mPF�;���8�L��`5|k�C�����=�%
Q��/�l����J��@��
3k�GU��0i�47�7�!߇n�b�g�	i��h�`��+?���;�zwS1�!���D=s[�j�`����um��Y��б�;�,*��oT��j��b	�/nd
�C��л��ªK��F�4�!����ڼ7E�_���˽d�]p��"�Ѡ!����߃F\���,N�n"����e�7��Aa��?��
O��Wc��q��|�M�q�4��Ӧo�ۆV!�M鮗򿃩��Ξ��ï
W��u.�Sݫ����ۼ��F��� ����p�4,�Ɋ
!�A�t^ˏ��.��jmn.4�|���%%��,�	P��MX^�r�@)��1�{z�eG�Q#Bl�r�w�'�yc�0�U�4*��Sj�R`��t{o��ZY�4'��]d.�@*''.�<�a�!�Y[T�5���1���c���t�\���akzk q$�r3~D�΀��O����z^!,��X8�?L��<0��ف&�)0{���� ̞#��V/�%�^���EiOme�C�O�o����E�Q�[�@	��I��"*�����jy�'��^����^������	S���&��*������Kb:�\'��q#@fYY+�#�� e �� f���m�.3���m����-�9�a��Ճ'v�i��F��ykf�?wXm��]��!,��T����x2I�$�0c��ʦ���4���8�"���S<\p3�>���P2��ZB�1�f5O�UayZ�H��Z��q��Wzt�\�2I�S+6/K��;E�+��"�Ѹ9<�I���e�������k3�ͯdn�kγj��JeI #���ַ
��Bw����Z�H�`")���4P����g&(�z�C�UQ	 n�h�g"��orw9A�]��p��;S�cC�Ԕ��X�:�?�����m{�@M�(N`Enol��HC^�㧺����� �?�Hd��Y��շ��M�ˢQ9JQ��HL��~
WgS��{fEuh6��؟�(����QNp~��Uu��0>Rs�ݮ�Ou���"^��lÑ��6Sk|��6H�A::H����rvt�Ȕ��c���Մ˖I��f���juP�j���1��oZ#�aH�н��7�kK66C�I+l��/
@�$!�_�j3 �73y�tVވƏ��j��f�Y$��PsF�Y�_	���-ìP]&��2�$�XUɑ�>��.��[�R'&5���9�s��kGٶ�j�E����yV�Lt�0sy!�0F�^��-U�R���W���2��?�1??��̙��`o-�n�+��1�Xה5��6+"P~��$÷�YTi��G���^x�����Mp[+P�ؤZY��e��䐚���\Zt�\k��j�i���A�A�n����%v�"�+ �#���N��k�^Y}��s ��,q,nӳWŽ�%��>z����˾3ڹ.�E��#\�^H)kaJ�hQ*2���XL�D�8���Q�^(� SH�ObZ��"��=���&�x�UB$�� �;���7|]�1G�Q��H�m��bwJ���ڻ" ��qX��e����<)������;����I|�&�Ӥ�Ҕ?6�%k�V|�����K~�R�Ƽ��F�GNcë�d9�.-�5�On���Oە��x�b�:'�q±�\٭��(z �j�"�Z�O�z��鳸��'���m�J+-�n��A��N(bִ���s�x�z����*��yNb�9b���y����%E��jr�í��{��)|@�۶�4X.����v;����Vm��
�O�w�=�Я'�����6;��	�G��6�1>�3��������N{�:�m��e��WD�!~��NE�6��fT"CG��+w����(ms9���;PW�(;:Q�N��ls�N4Z�À�`θ�p�J���]5�X�ƑQ�I��{P��A}C�O�+��,9��_"][��cO��<V��:���B����-���9�ï;��r��8�SO���f�f��lB�����]��a��P��k�ۼpW�ͧ�R_u����c���n
̶g�m�V�rKͬ^��K�Pp��tr�q����K����?�O�����]����Ak3a�K�M���QD�� Q��9F2A:��-rK��?� w a+UP�X�]R�7��'sڱ�SА�̸˵�9��t��`{{� ͱ�:�ewP�iG��Okm��l1��>���1�ϯoK%;��)�IL4+�f�#��<y��t1� ��`n�Q�(�:�ѷfR$��>��wT�fb8��>���gi���XCO>�3���3�*8�o�g�%�1J�O1���S%+�����0}&��y2r��W��A	WN7n�{�]�\-� �d-§ 8~q$�Y]|���y�!e�u�xt�2X�WI�Yi��[0��>�����~�z��d�j^��2���J�Q�B�O-���Z��r$fj��;�.A7	Ǩ�|�I�� k��B�R����s��ݒ8�+mE آ�In��}*U(��N<I[�zpaP����C ��O��80�VG�	�i����<k�)els�d��n��\�����Q-�ļ],ml���J�Y�3�[Ɣ��S�fݦ�g�� �KZ�	���,�������h���]��[��	",�m}JH�Q�����m�P����m�(s(ܜ�zVu�7cK��"C.#�N7Jf��T<@M'	]}�Z�bcȜw�̫�Tl�F&���	tM��/����MR�5��#�_���*cV��I{-$MwMH4�����h�i���_���r�?��NKm� �����gQ�Tr�N4x�a�lӠ���d�.ĥ;yC+Z>hں���(.ѠEϠQ.�WM�*6���0�%�o�cz���Ev�)[��y�S\�K�[ŏU�e?��&h��-'.Ҟޫ��2Pl�YGR��F���;c�k��Ӫ!yI�`��3?�&-]i:�����K��ţ) ��7��q��V�4�Z��-a����f�>Jz��1�Bl�~��0�����(��9Ss��,St�l�,	��u�U�觥�hsU��M���ւL�]u��1 ��H�	�
b?��O�ېv��;W���/�\l���cIM�?�ќ�,�g�@FV�`g�|�%�?�Y[ZKKLE)��G4�u�tz��GjT)�� ���}��t �G�BY��"��&p��P�\�u�M�h��1*s��rF�m���h������(Z��~��i4�tB��#F�;N�v�!v��&�LO���Fŋ�ȇk��
h��!f����4����	�m���vGf�Ttw�6��v��*DGc��:��ތ�S�p[;6�d)�AGm�_����mp��Ct?З�Y��H��o�n���i�����vJ�I"���-|���0�d�l!�B�,S��}l�G��Lm����M-�5q�*(�G�i�3I�N⃽����j;Kv�Y�L�]�@�\D9d2Fd�U��/��h�*'���"&+j��i�6�͓6Q<j���[�O�t	�����ζ��@x�ϨWd�����u��j����à�}�m�Ek��!;5�]SNЩ���"�ə��'��5%hꛇ?��pQ��dW������8*�c�0k	Mh�Q�LN�Ĩ�(�њ�2 Y��i$6h�r��D���7�З�������j����:�+�5?#W�r�(jz+�����C�v:�8�����+7�qne\��Z'՛(b��S�L�	(jJ����WƴbU�Lj�r)z�q�xg:xR�q���弎L�rܷ ١�^������f��Q ���&�J��`��7V��NIe�V���\J�z~�!�L'�7�PW�n��%���ؔ���\9�z'z`�ˈ�X��>-������ѶB�5�^!Li�ڕ~i2���X�����S&��l˰��Kܪ�a}o��u���O���gfn���c,2>媓�.�����WXi�j�g�A8�^�bO���Ü�2�͉Vo-cY5��G�4 =�qO�3�w0���ޑ���f�����m�X"�3�S��˃�f�Ա1��5�_Ķi�r��t��a�i�ă����W���1N���S�M���EW|$߬fط4���5Ht�[�B�+Ы��a�O+I[�R{���Cg��C��Mo
�\�dп��8)���WEI{��+�`3��E	N���'�>c�a��J�nn[�1��PF�M�a49�910Z.(5�����i-`�ݒ����ey�2�g��n#7kc��	;�0�.ǺW����T���j�>��k�O��\����NT?��m�O��j�D7��%8�Ƴ�n�����aΔ�߭h��bid�t�źt�&*c�B�gԱ�B���!�F ���[��Ec %��VZqI�@���,?~��=�(6zP?� R�i@�K�<��K��m�ē;��t��[U����N�Om�)�6�"x�F��&4|5eb9W��9�u�Rz�]� �3�$���
��ꋬ2,v��%Z�$��4���]  ��g���5=&�di�6zΦv�9��n��~Ѡ���qb �q��!�y,e]Õ|�0��U�*=ei�k����!�Pp"�zQ[j����| �O�c���d �F�||�W]Ҽ��r3_����J�݋I5wE���]��f���_q��11�K���7����fy@S�-d�Sjp�w���N]�����N��][��~`E�6&�(�I��U���Z>p���$�F��	y���'T��^d�\��Ԯ >֬��s�UV�6�)zm��У�04W���B��|?���g����|�	���!c�,ab@�Ǽ<]�&e��V��+��Abpu�M�֝s�(VQ���Oi`��򐱂T��wA�N�{���1~k~W̬���["�/�	��s 3���y?z�I2�}���{K2�sHAĉ�`�|�v��������`Z<�c�U�n*>f�~ɑ�ff�f(gO��9�@�S��j���U4���.�4�A�ќ-��8���=��V�]X�c�C�:��+�ݹb��&�t�B�5�-��-zewuT�B��SV%�l�K��+���3W�:��o��M3�*
�N%ZBz��p�~� }	T+�O�{����`"�~�F���^R*t�д+v�
X�< Xu s�'y/��� ��g���M:��h�Z��?��@���Fkl�'&�bq|�4���fl��>�*�,��EԖ�-�>�FE+Az�J�0�aV��'��f�Q���C���W���M	�^���PT�i�iᢹ��o;k2ܖ�>ų9���j�)��"&�]2u¤��9(��*3�n4��x[�{��W���fK4ְD������<�����k��a��V���,�k�V`����ݺY�Os��w�m��=��5?�:��Z)�e�#�)���O�� ��/*~k�M��˨B���Bb\j	I��Ϯ:�p��R�dݬ��e���JR���7�7��ya�
��9��Z%���`�YF�Ќ���
c$k�#�EA�d�UJ�z��\J-����_ruM�/'5���A���Xa{���)�OA����D_��7)�c�U��U-_u�7<1D���+t�-�~�~��!�uӑ���k���Y���yV��g�B���U�u�B?>?uT�j�^n� �
�%)�#�؈MbI_>��1MӜk^,�#w�+�<�4 ��K*�T�K���
��s�Et�*�Z�հ��Q�\?���G	��v��v(��h���"<L�ڑw/�y��	�N薬�ӷ��}�����	0;�nѧ�
���l*���
���R����4/��( 4A��	 $ �z�GEWzOEr�I�r	L�VV ����ep���DPmy ыiE�sMu�����K�;�W	�m4�e`l͖���ܧyޯ?fi��^���LD�ߏe��Qt9Ѹ�$)�q�D۫X0�$����#�X�8�_`����̆���YZ�y��j�P������q\DE�P&^���_	�|ΞE�X�-Q�ZIͱei�Ke�gV?y��Q��§67'cWJ�*��U���֞��8�'KL ��ky�Bn���+TU���<]��-�KЕ��.qI?,�㫌S���	B��5�a������
���Zd���]Y�oG����<{��=`t2���ߺ�͏F���q�׿vW�=+H�Js:�����6�g�[�`t��D����/|���a�ļ�H5����+����sP�K)�I�ɍLs�k^KQ�٥�oY��U�����Cū�+���x����%��!������9����Ƨ��WC�H��S&�HB� �ɖ����m0��V>�#�����-pyGG���p�A��}L�H���#��ie�,�L��-�S�Q�� Tf���� �T
�D�ۑc�,�,�)6����:��#���Иd����x�|Mb��7z0H9T;%(z2���*�FN�y���2'þ�+sz�dKe��9�'�����2^�t�vG�ذS��~��u�9��5;�ё�!S  ���B��őT����i�x�J��t�7\��� �����U��|B`��N��Cpz3#L����L�$��h+��n�ƺ���(��ں�@t�TOմ��Y,�[��kCۗj'bΤ�Ǌ�tZ�S,b����5�1��i�_����8��E�u�i(|4Sx��^3�(�>F^�I��.����i���s	Fq:)����;���n�։C��1PE����I!�����H.��}��+:�'�+ط_�h^si4A��q���.? �a�N�9�@���y�)!A���1L܆�b���l�)�X@|YDT*Jm�m��%��x��z*��)	ˣ��Dͪc�j]�lιJ�\-d�.;ǂ����0ߟ�=c/�����,������KrI9�O�(�0���o��]��OK�d�y9N�v�)�i$<����:�4�GB�ںb��5eF��<0�h�f-c(2(�*�-"��Y1�=@��*��Ts�I��y<S:��:���7�2�jV��KU��Yn3��k�'� j��/ܘ�����YT�X�eBę�!�}*�k�_�rH�3$��0�B��,�7�*�%�7�Z��d��Ӏ�,����T?aǍ)j)`v�P��=8 �:0kY�~KעS�d��K�b����oF�����
�-�'B��I+@�P�(��+��%[v�I��U6"@]� �,�=�/��z�h�q)`.Q�'�h(�?R���	�Ԡܴ�=�q�_�����#�u�lvM��w��xZ1��P%�eH���F�_(�;���@�,�SG-m�<��}�v�]}$�:�ە��ͪQ�e�Vk�j���I#5��=+��OM,A�aL��el��C ���pf����f���f %�IY"��x'02a��M%��JkT�qnp�kQ8U��`5����ب���� ��},�0�
�"˅�v�e�Os��.���	�Mɋ�;! Do�s�ݷ:��
�yK�F$�¥�*˗z͋��Lܫ�k�F�%s�f���J�H�v�n�d&s��p����9+�(��0���t��乇e�֧�{?p����&`ڟ<��hD��Šݘ Y�-)��)�"�)�������69���N���U���q_}�f`^���n^���ӄ�Iɱ���}?4�$+����������o�rO�W�P��ɀ"�r��Փ�7�ӣ�xI^Ұ��h��ח徸h��3Ć$<�m�R��%�m(� Y��v�,� ~�*JX��ր���i2�}��XZe�k�[̟��Eq����	�����<Ͼ�1n�,��H�(�p�$�������M�9=�I�p�͹iO�û�0�T��I���_�:d�a�gi�������x}��9f�f�N�f���N1�nk��f�$?	e~c��,��|C0��j��<Z����zQ8��� ��g�F�S���&��d��\v!��	z����AF�+x�^�t�3�@2)AD9������8ys��U+o�=��SU�uL�ޞ��9pr I�'i���	x&`�Asۦy���xS6u�G��ȸ$�z��y��>��f�H{Y�w�7��Ӵ�[���c[�7�9?���o�����Q\9Q�z<�P�[u��E�G2"��>�ڇ�Ǝ#��ϳ�6�������v`\A�O���mo" ���-����z���F�[���䒱��߿;A��A��)5R%-#��� S�g����*K]%�Z&�w ����ǈ!n4mU��㳆��{�`�X� Qw��9჏�-����%*	�)�1䯴���2��l� 	�w�/
7z6<VR����%��_d��Q[��C����u[X>��vn��Jw�붖vX)�Qx6�O^N���xS&Lui�Q��n�%�*�̭  ��s��Ԫ�P���'A;��ZO�a�����R��8�N��L�F�*�}�:u�Ř[��5Ih����Z-Ӿ�*�O릍����$괕e���Wt44$�р���-#y�y-'x 5Z;
0�*䋊䥫q��8z+����U\�:D���dg�t�a�C{|W��5z�)���R<��D܀�A?<+�w��1��/iy�ތc�b�nPn��\� ��4�n��[*id�@���ma�A�&�|��p��s2��~-������֦_�UKz��y�����D�G��&y���7Ȃ%�d�6���E���0������\�3(Ξ�WM��&ftq2a�~��D������\�$i#j��7��W��_S��5�m�.�Q���Gfs��Xj�jMe�4y��s��Ԡő�}e��*F�q���5	�yKv'	�s���9�u��ॄ�ìO_��^��� If�	���ԥ�W���b$�˃���r8v��O��O�`=���ڜ�E�fG�/�X�eD�*����F"?!;�����A��ݺ�@�E8�!�[�|���i&/��>�����p8�]��K��i?�R�����
rvhp���u�#�̝h�m�M}j:��Ŝ�8�Rl���>��A���,�޿��s�98M��}���Z�^���S��w�~�>#��8ʝJ+��A�-�x�����#y�X�\�B�e�=M2`v��b���K!��,1��z�ۏC��|?����8	�ʺ�x�c.��C��H<�����g�#nM���׊�%?j��u\X���_���-�Nׅ紓�����vE�lٶ�zr/�d�}����c8���F.�zr��mw{L�EYV�C1�~�g��S;����S��ȃ󯗀{�_�"dcq��q��;�j���1ޱ�AZK�̹��I�������0#�|���(BLee,���S^7�E��N"���8^�V/ʇ�U���:���h��?���lQ�ahd�	�u�����|g0f,ݢyjs���Ƽ��[j�T��OWzҝ<;:�#�Z��.����P{���ў����]9�C���⮠� �<A���L�,-Ԉ���ڨ�\�B'�56>=�7MO�I�7�^�]�l\�\t�`�T:;��DI�,ú`�b��y��Ćq���
�d2�P���
��zm���]3IQ�/��6�|��o�;m��IL,��|�2i���R�[�čِ̪ovi#Vxa�}9)��fkӧ�C��uta�7ؕ�&_��Q>��-'�w^	�;�A��{�w�_ �8Y V@��2s�J@M��8J�b!..<C��uԝ�/�.��F׊9���yrkR�o���-��
�^I�)��/ax���REeLy��&Oz��3���O��Z#JuZ���k�rOf�\��LxC��>���~֞�C�O�p��@�nA�b�on6��KL, ^����{����K��2F
�d�j:�|\ڂ&�Ŕ���J��ٺ�(f����Aj�PQX#�K�,���-8�_;fkK:�91�[����������7���bJw!�_�4`�
�T	wU��1зgfĿM�9��9�bV}�wM�ţ�-���\�F��K��З hJ-*��#6��	�ԙ�HS�`Ȁ?c4È���:o	��l��CIM�ʚ�a9�D�H�DoH�^X���.�H|�`0���l��#�ڀ��(~�������4I�@����ǣ�0�{6�t�� I��GʴK%��H0�tS'�dָA�癏8�NT���T������Q����70(��*-�8����M%�%��D@^4]=c\�W`�[C���ލ��3=�IGHN�rX0�Mť˸�;Ȝ�qR������c=N5�<�d**XA�6�?��2��������I�v�(f�F=MG�4��5ğ�E��^ù
����ϋn��oУ���Oz�x9 =ɻ��asR(��\r�Lň@�1S��V�����E�lKC�����GJ������U�vi-h�f�%�z_bG΃L�D�<{=\}!��>96}bk%��E��۔O�^s��J�%������1����%�҅(�';�9Pa�n����\'7�����(U6�w�e���G(�$��VE�i�p�����ȉ���B@��7��L�`��O�Z�����#
I�����:�!�����)?�-~���zFs֞�]y��`5 �smX��Ђ,��j�2ł�K�~�Z�,����m��1�8�}�Bd�>Q3��5�ғ���WV���{�_����w2���Qa��ʪq�@ϫ�u3�i����}��ز]�5%�P�?��h��s/ 0Z��I-���x��΅�俳ȗX	�E-�������|��&}��8�q�8m愫/�r�7]�wN��c78�w�;h��0��f���`�`�I�����x녌��]S���%+������QY���Ϙ�7�t��P@�0@Oμ��([4M��\�z�g���6�x/Y��t�)]�������jt쀍��ޑt�l]����/hSJO�4i+����^R�AWP����_gK,��Ȧ�&�QZ�L�>�N\�+�_���$"�PU}����k�*ZSU�Ak��u�����lH�K��q�H7�����'!D�9����T�E�w�d�͚��[_ ����u�/>�AY3��W}�d�JzI\#,�_}W*����x�2��v���w������`��Ǹ�at�Ni���z8���,͢�,j�,O��j�� �ĒcwK�G��T��O����ǍeXq�BN=!�Z�
K�қ�xL.-�<L7`�ު���ݺ4�ǖ���!�4����rO�wsQ<����c�����\��af{5�+��Ȣ%A�)�a�9eƿ0x3�>���BB.��������������u� �o;ԲH��/�] [�f��e��C���J+�?����P������]���^�|l�ʺ�h�]{�~;gu����B�5�P�8�E�:En�&?�����.�7Z���\aa='�w�n������U�����?jP[\�i�4@s����K>�>Ҁ:�(�+�)T��¯n�a���@Z'>��/�
�"��uŬ=�ˠ���#�M9K�͗�q+�`%�#d���jnf�L�;�T}�U⏐����qi�t�����E��/�h��.�nR7u�.�d�P�N?o��_�9%Hx`���	B��-�N)ŧ �8��[ň�`r��A���k7﵉�O�fM��6QP���ps�>���6b�PԏsX�"h�1���I&tP�H�Y����gP~�����_۶;;H�}���_4�U�V�Z_>:?�Ɖ�A���
� �$7���+kZk�X��r(��+��X���r3��q���y�Xl.�y���+�e6mut!ellu�.�tc~�ٌZӻ���t@	���������^�}��0i}[�5��\���1B}Sb�O��q�lb��I�_N��S	�M�"���"!':}�^��>�B����	��þ�(�6���D������~��/�NᎂH��?�����,4cԙ�Yy���&l0�X+B�X�Dқ�	�����m���S}> 3�������y�8��7gK̽R
~�X�l����H� �;[T����~���@9�b�u-���m%��6�ڝ��������Rc+�N&�o1����9���	44S#3��ٯAoUmH�"�|{��Я��9�_�^W�S��� ��F�?
v2qA�g4���2�a�
P�� 3��u���GE�
STc݂!�VlƿBt�+�|��4��(���Aۘ�?�����R��;�z�F빃w��` �<�x�r�[IJe��ũE�Z����_�O��h�
W s^��w��"����0Q�|L��5����K�y
�4��:&�;'@�6���q��Ʃ55�\	�d��_U�:\.�=��- }YW7^�b���{ol�;������P�q��n���Q��B)�|��,��Dp��7�P���|�lo����.�q��i̕�e�yn��a @��P���p��R=#?ѨCx-�,�ón�M�o�sRŻ�@�6u݃�i�}�Q�Q��W�	3��t�z���A #�7h��?�������d�����M���}�Mx�Q��dJl�?x�\�SH�x�mfMrL"�4��f7��iZe甆M�P
���Z�h��E��k�(^�x)�D�+5T �q�M@��L�8O�P��	f�a<2����Էj�m$_���Mo�A,n;������957f���E�}�b-��9�I��'��'M�������v$��xo<���\y��7��LOJ?[U�n���9���{&���6���2�o�5H���q[��9��������1��zzִ�^�'pj}m��ՙ]��̡���8B�*���"6�Q�t^����u�caW�t�z�����#��t�A����?���$E�(P<	��	ϋ��EF�Bw� �ؽam,,���mK��:�+�_L�rx]Ezء�����R�zbal �� �]s^��}�٥oS$Vy�
t�i.��jo�a�dԑ�tMj�~�w�1uR��dF��¼��á�:�`=!�ۿ�ϭ�̥���:}/�{(���}���U^�y����M3�����d��I'���`ఌ�˛��?�_���WC~����zE�~ĥ�%M񙣅�5�6ĆrW(�*����?��K�K_ؘ�h
�?zc��տYW���+R�Ĥ5�n{_ Q�AUSE%�n�o���!ր�y� ��_g
5��U����T�j����U_&����F�wA!�Ɨ`����s8g��m��ɕ�N��\�����n���!ʘ��Y#��lb%ײ��8�h�.8��(�� \B��@���剏�b-̞`{&��PP���d~��~<8�PN'U�%f���b��P�ֳ���i_������@�w
�L�@n-&��w�.+�M_��L�H�=�;�Y�@#��8���K�l���|�6���PO��;�-��am�YuZ��/�u#s��}�����}��鑕�����?���%��^j|{m���jrЭ��]�vJ6@�
H#�r^��Ň�[Z%.o	O�4�߾N��Ť�s�h�D��	�'t�P��k�|_�4��y%�A�ISs�v��2GK�&��'_�0�텾���3�ۻ+�*M�wA�<���N�W}��L�8����(��_hi���}�d������5e�J�Ɓ��^�3�x\�WUcD]��#<��Q5s>�H(��y.����a5v,�K��?����h�B&�S��u>��OCf�!����lj6�g#V�I�}��a�ÎG(bȢX!����� �(���I�����^k���\^��s����ҧ�w��?�5��S��ň-m�Қ��^� ]D
�r�C
��7P/چ��'78½�<�2ZE��0����Ϟ;K E� \_�����rx!ү��]�!��Fϥ���� �Ȁ���-��C�%��m��m�Xw���C�G��%7F�!�� f	�B���,��iE�>-k?爯.l�Ii�EW6�*�F��|j�gx��B/�bֱbvM��e1ڪT�����4���l7wS]QyLI-m��>0Z&f��"H�����$�mδ?�� d���.���@�N+����m}m��I�wD�TX�o��37�{��������g��'���	V&���0Y'�)�WY��V��UdϪ��@{�.J�c�C���̲Qn����K��(�E�����~=��[��c�xb��o��1yHǚ��.��4
�W��n��>CS�y���)�R��f�ě߻�9lLK��H��$(O�5oX�ְT����.j��N77V��N Η�d&^���R�^�W6�43�I�x���ИY%���ש�*T��xEE�)�C[ٸ�����JA	��}ɓ�y6C��eЛ�Y^���%�[E��/&�k�B�-5�%ZTǗ����l����ʏ���޵j�P֎�s��*��Ͽ˝&�=Kзĺ��^�������άC�%K�m�Vgӱ��R*����z@Wȭ�9M��w�!��VS�Y��1�.��+�ϔ� �R�^�!���[c�?y�³Z�y*��~�'�˕�K#��%�{�N̷�絣�lД�HS�W��5��!UQ��Mc�6�-G��Tw���Q�+�uG�����Ԯ�@���Ik�N-��D�;�ι��*L�rC�Q:g��r�!��3:�7�عWi�F,��_�*X �9�Z�=�>�U������f���0�.��lK.�����U�����׃��m������´�DP����D�!w6I�XC��$� �F	���w�ᄧpE��W��P<I'������&�~r ����:��5�/�.���c�e�*<����J��)�l�v�"`�G�@�h���E�;��*F���s�JH8<"�w9�{���0a$C]t���q����,D��R���9�A'�~P9u�,/n�F�TnU�yL^�,��Gif�t������ZH#�j0�:e�^q����/@�fW�CWg4�;����B�-�ug�q 7����T����b��r��o����3�6���qй��`����&���ԩ�J�e���s�pP
]�~1�\Gf��q���i6ٶ���Zm���)ڠZٔ*d0Ez�'�Yќ�_Wg	���(y�`� ��{�y]��_qЯ!`���������~�vX�*C���Q�R0d�;��LI3ez���~������j0T�1=2�҆�a�Z(��n6*;׷�w��� �.\�k7�SJ~�gv{�S�����yQJ�Ig,��Fl�Ko	.��y8!�G��Yi:�M"��W��U
9�ϖ���f���X�8z�����V2J�}0˩(�+�Ց)�Ā��ca�'=���f�?��<f� 	<%G9��S#f���2���S������R�iK'�D�Y�X�`���Dv�T�So	��Rhٚ�:���(�&a(���/	�D!��86�%�Z��:���렻�#�g�~��^��V����|�2�|W��Ǵh�����^i���}��_;��Q�VSՀ��n}[K'��l�3+`Z�zg�V�~I�{7;���2MXG��=�̽'�,�ɸ�
^h��U�ȹ�/yn�
�q"�<���}�����&8��\GV�pf��m�wdmb�H+�c�L%"W��AHn0� X\��$����[0;�����O�x5��)������{�e�UaS����Dحe"|0�|F��X�8��R/�vp�b��p�=9������I�^,��B1�Y��z蟘���˸%�%��]��ma���kog6�d�����$YɎ�$�(�tG7pi�0���83%<kU���b��v��mE~����t�:Q���V #w��N�����0�{�J����V������.��U��ˢÁ9����ѯ�Kc���W9żD�qa�b~r�A�Jn�+:���QV�!kx���6cg>�U�'���_'d�5sX�s������野^��L�,�td�񠕘�@��D�(���@J_���k����E"3�bD�k�Tim������|�e'9��"�xX��{J��w�4=��´uc����K�M����<?f �fj����͛�V�Q#��(������J�酟r�����^v��f�C�\9x|=���s�x��A�� S@R|��0��Nn�I_eK���H��%�" g�����<SL�)Ut�L�F��)Z�sr�&��.�.�H0�ޙ7<*,������*������=̺^yK�/��H&�H�d�]���?�T�# E{���L1��6�-�H�[�L4ɝ�Q8FSH�e��������C��TR�@m����INqrL���33�P��0ČJ��ZH��%h&��#��D��>�����v��S��l�"��sɹ�����^~�+��4��.6�ܧZP�m�r���H�Աn�3'B]������zd'�cԶ��N�����s�����<]�@�BbT(�b*P�	\�!X/�L�j>x���ʐ��#`F��j�3%'�~BIW(}�t@d�H�55��_sB�û[�̟��U3 �w��9~]5{v�	F�ݍe׮ YTs�g����>G�sgѯ��9< 턃�lQJ�p��a�J�P?v�Ih�=�ׇ����<���P���g��� ��O;n�Eܸ�bV�2��g�ξ_gΎ��z�R�sn�}0��ŁAs��-Ӕ,��y�QU���٩�1��k��cnǕ��lz�s���R���� �dAԝ@�xf����JqZ�l����_H(f�o'�	ϸ(�	�a�#:�N�9�KիtouCS����kyw�˻C�~{��pHL�Zx�c_(�9���R�������G!�Ҧ�Ld�q�;�B�|_�̥��@E����iM�8��:P� a%)B�Mg��>�xK�\��@��9lLҚ*/�*g��1ڈz�fb-[��~44i׳��C3X�1J�݈��͞�5a��+e�18e	o�����%1���/��$�!��:쐏��GA���j�(F���}�Q���R���9�S�����h�7Q��
�"�D��C�� aklwCW��%�J� ���1Έ�����
&&�������ʗ�4��,�y�T�Ɣ����3�l�|�c�	��$�j����V5�Z��y}%�H+L"�<� ��w�g���)#�R(�&AN�L�D���(��������`�B���v&R+��' ,x����\C�@ڂvZ���d�0p�Q䙠(��d�/o��?;�$B�H��D��tXU�H�����A-87�2�|P ݌��v�E52Ft+90�n��/_T�LZt�w��^<
�q1�6k����;Ȯ��PE���@���O�ʲ�\X���e-��HC����g��0���Dūu����zo?\��F�|�}�,�� �/� 揔f��E�exw�l�#h� ��^hU�/��U�O�����<����E�j���a����4}#td�e`�H�O=��4��(wG��I�%uc�[Jl�+��0�|���Ǜ�S�b1��}�CV�Nq�V	��3yg�"L�+�X!��e�Z���*�Z$_�����;~h~�$�Oǰ��5�X4L7iB#��",�[��q�SF���v�K?�SH�ǋ��o���r����Z�?J���:I�{_G�HY����&��dA���(si�. <T�-�R��b�s:hPy抹n߱��"'��4v���-F�4�}ґW'=$��y�M2Ta���Ғ	;��5��� j� ��d���f\�e�h�M���1��@��������ڔ�(�j���2[����f*ȕ@¤{��Q�j����M�8|U�vt���3�eY��?Ƭg�&�eb#������fjls��>�e)�et ��~�e9�����j�.��6�&�v�����6ugF��G?�Yl�U��ld��;Ja+X^n�h�S	]On�^a f��q#>fד��u�/`q�t�Q��Jv��g��W^}֠Sڄ�c4/b�,@
H��6��C��.�����ηI���b�\(���խ>?^c�Ń�g�m����s�+�9�IE������eWCTc���� FCʣO���"RBq���0��ml۶��T^�E��5mn@)r��l;��o�S]t*B�4cn�tU�Uݒ�؀:��S��趺�P���&y��+�1K���l����R|�DK3Wwp	�����B7P׌V��}}Z��5b���������0�����J��Vw����x�x^1F)r$:�
����y�*ߦ.U���k�բ�@���G����j� �?�"S(��������D��>Q�=���pס8P�v׺h�@��4#�+���P��U���>�����Ӗ�A)&t&�}�~�2	
�k�N�N0p�"E*�vG~��VM"<�9؈�a�J���p����e�ᇌ��
LO�EC%�+���y��حݣ��Ji�p���ƛ0ͣҹoZ��p-�X��W�7���S�r�A����>�]�ћ����%�?NX�n-fi�&� \�?(�(���/U|��=�C=:i��n�z�<R�❭9�ׇS"ÀѨ�U��eQ���|�7�w�Q��j�B�'D5����๽�]��Ѳ��!�a�^n�`��U�k����o�d%��=*�]���岾�B58�\�@[4����~�	z������ G�Y3�Ÿ�<<������qI��(��H�oуY�����4��)��;�`��h%�ⴡ��;0�����+��P�0�G�П�z�5�_���j�tw����C��Kљ��jkK�Jچ�q�À�3��Mȳ���_퍅�a�.�P�E鲔��R�0�͉��S�Y�ݳ��P�ߒ�hZ��0:���j [�d��A�nA!ƛ|3������]��E��#x	@l��@��l����E]4�w5��/#��:��=(x^eY���~�LU�'"���?g%�oP�u�-�* G��Q��}��o���X���B�,5�܈�q�JTC����%dY�!z�/��w�%�T�Z��,��B�#\���;*Ķ�\����P�bE���݀��G�'��J���� Qd��(&�L�6����s��JqQ��*4�&z�dz���X��A\S�3�10�L�H���I�{5�t���z�G;���i����ۣU TK���|dU��2"U����G>����({��NƘz�>�T�(�����ơu�T}��ZO��Σq  �iA�	����Ù��#t���� �+U�2������W��P����t�;R}dK�������⸮��n��(�%o�,@��Z����J`���x>�I�=�&{{P��Z&_�&{��1����Xٻ��>LF���t�rX�F,)�i���� �?����Уɔ$U�c[_&��k����cD(ω��2�M��4N�i�G�M>���r5����XI�	3�U���KuTmq��i�F�4�U���f@�_-x½�i�LA��*�sc�9?��%'�A�T3�5�y�tP��T��S��7���!�0��zq)�K����Ld[Щ�ajr����.�H���/N���.��B,f�Nj�E�O6`����@�����~�i���ک 6�AF��zL"a�hj+Խ�����t�������U���	�W����ޑ�a6�3��0"5]X���@Q��[����a� 4}H^����H�&q�xA��^�B�5��	�ޤ5b��ꄆy?���g]�Vb���6D�b�L�ǔ^=��<c��Q�x4��fwWH�į�m���"���>CR��U{O�B�2�&	�aV
�	�|��mi��=,G��L!�(H���I��#M�c�Ô�k��nv����t��,O�0������e/t-�t��(�������3.��t��$rou-��M��@{`mq��]��t�U��5�c�\����� %��18�\Wq���&�.����^A��3���Tb/�J�"/�����k��ludz%��MG�{��V���[�5�s�Bt��v6<\�B�|�U�1	N2�hLz��#N꽖3s��Kw�r&Rk�-�g��·q��K��
��ӽ�� �R�Od��tK�����e5���CC<�M���qQ"؄��Z]��q?$����*�d~E��~�B(�X�RF�·F*���*�o�\k}|����#�Jr�*�>�E�n��/}m�H�N��� @�&.3�c�3=��L3����Qq��w4
���mp�r8��.$�T"����]xX�Rd��l�y�!,:G�&�w�d>���p��o��%�I��r�{�T���2`��l))��B0��b��2Y����iRx�+nVI��̃���d�yb��δ(�2ZM�oʹ_a04��!���2�(���{���>ύ?���zg����Cl��1���"�%���Qn����s�ar��G�XC՘q�����t)��Tl�9%���8�Ge�	�ӡKvVD�CQ�X�[���UZs{kǹ�-#�O"'A�!LK M�$W��p��ti�`��VؓC3u�oN���㐺�!��+�o�w4ô+)	L���M<��T�˕�oƸ@�P�ɘ޴�)��k�ZĆU_s�'��K9	U�ϊ���M@�rQs�V��e�<�I��-��R��S����E�${���##�D�/ &���;�(�}�Ū�F����_E�f$����ƾ��}lUF����9�SHT�J��ݿ��.�r!��7����@5f���C\�:����zv퀠m
s� �9*уjU�4w4��.�a��O��&�K�6��	���Yɖ'�[�}9��6GW�¯[+M	�"�
��r6+���?p�Ywh��l� K��Ґa���a��dSI�����ϑƕ�"V+,��?W���]I�5�����形�wRl���%�Y3x�&#f,�Z�����{�yԿ������
�̋����Y@<hڒjq���-v�p�V��Cvp�J]W����;e@�1�1�d�{�k�Q��)���g�+,Բ���y��=hv�@"�hl��=�C����d���b��`��bNmv,�>]X-4R���Y�M�9T�;t�0.C�9�ȗ�O�a�|��H�c�\b<�?2֥�b1PX�N���YӋ��$�Mi�Y�`��A�\q���������i�tL2���%�'�r[�j�"G�m&�*w?��iW�a><�&��O����ޮ�����[�����G裊��a���W�?��v��o׊�������'�.���>����w\4l��3��V5�&L��h�B��0{T��p����i��-R���I~f�ݚ�qH|Q�{U�d����_�x���ʳ��G;����p?N��.�
#�c �=����*JYz�J���N̖+tq>�)��;��B��w�Pr��C6
3�?��3������{\�����U'��U�AN�Xl��썱v���e�
�ᡟ�M� �t�P
_�ޭW�Vd��z�%2�2"i��0(��U�W��IXCu��^��kyB~���z,Q�j��/
�Dt�q�*#L�x�(���P�4����y�%��q� ��?�N߂6,͎�X�&�Dx�w�(R��7�*.W��@���"�[�R9���n 9���L8`M}ѓ��#�4ɗ_09��P&"�b��?��_�����\նpQ�Y�ڿ��"f_� 9��s� �����{aE�#��aT�Vx���vp�X}.6}�Oh�a�f���^]��I\	�I�A�|O��ifPi�`���*+��N#�V���g��d�����g��P�����RA����m�-9>�bD�s���M4�)�zw?��O!	��{�Yd�M�x��An�����-�%�@Rr����Q5T	�s0O��;gTuٳ����9cA������EY(z��]�2t���88�g���G���<�~t+;!����Y���h��%�=�`H|�f�zMG����]�b��v+m�7{X�gU`bd�{R��t�(r��ťSV�^��V�H���ȹ��АӨ�b� ZG���5��>jP<Hwk½**�`������&�G���5�^�ھ����AD cf�����+���AN��_VJ4�5�<:���4���6�U��錒����w��M$��Ԏ���%��$B����^�_8�)�:n��x|T�����"��v%����
u	�xr�M�[�QA 2M�?z�w������?M<ƐL̈#O�%`ͬ��_�7y�!-�yY�MM4.�#���?���S[�
Yu$��/9u)�dS�!.��x޸W�3=X�d�3�㌮�1p.���nD
MI���I��0�*~��܂Z[G��(a��-���'�4d��ꌉ;v�N���#2P��Q�ԡnJ�c8�F��R�Vpb��<�;��2=@֭�ے��"������e����������!_)�%�>� wH�/2-�?�,��`�W#��#��5$�KI�����|\�B���g���E�G0�y���x��m
~Rʀ�{k{l�;MW�Agi��n���1d�C���;�c����l����q#"�odt,E���z�U@J^]�*��w��و�❠@K�����Q1O:�N>���fe�Vس�˰rv��P~D��hz��xF|���qw�k+	�]o��`'o*�^I3�_h���kI�.il�@��<�\�B�H��"�A�x� �._U�GidXJ�%w�S�ەt����tg߿�v�<4�_���^������P���)�8�i��f�<�[uy��� EK�U��>�e�� ���oy�0x1`tuk�������x�(<~G__�0O��T��7E���H��ELY�Bߍ|)������p.pt�]\t#�����?h��--n��cS�����|m%�J�ٝ1x�d���=%+e�@jO���ܶmӤ.O�B��7"��8��;�&�X�k�f�`u!�n�k�4[�2�Z�=M��أ�z����;�vI$t$�\����\�|�Qr�J��e�Ǡf.C&��۱�2�e�� ��R~�:aT�?'x��o��Fo�<��� %����O��j�vRŕުu��ag�-��%u�{~�?q��;U�{���x�J�͒�NEF�a���%�3���B1����>�͏����!r��J*B3w�_���&�5)\z�>��F3Ŝr���z%i�[%�
�y�W��0ʌ5����~�P}L�u՝�� ���6ݔ�q)��G/���U/)�<����(��r{t�ڊ  [e�)7|p�H6��~�	Ƶ�6�����<rt��.��;,Ա��Q2��Pt��땙b�P4;�ԳC/��R(^G5*�^(��Cb������0d���wC
7K�� �ƴй7�P�)D���^����I()����i���҃�|k�;���	����~f/z�N�;��	0���1K�$�ȨHe0�����Yur�6TS��&�g������������GJ��N����?��m,�H�'�%��@�%=@���ɛ1�92����QV�g�m����ۋ��6ƶ�A}Ǆ�d�w��WEF��a���p0��'#�`sy�b};�����#���#�A�-�%���G~�9�r÷%��{<aE ���~o��,��#�K1��s���˟t���������C�Π��e(�_J��+O��~1n���[c�1�(�k�Ϟ�k�������1���$����%J�hf2����`���[��4m��hG-8������P7f:�	�Cq;�Z	eߢ������1!�v��	��M�0-߾ǖ��r��'�(����[��/͕7��X(pJ���n�{��O�v�=hg�5������3��P�a9t�OL<T(���8��{n���ճ�m*���»퇽(K6�ʡBA�])+���%����-Փ��J����=x�y.��{��4��iJ ��ұ��G�ߋ�M��-�vHZ��mL�*��Xs ��v-�_J_���@Zt��bM��{�����%���z�Q���ɻ9�����\c��*XB�P�����C����Ah����Y�4�3"E�<3*���/k!"_��:����������7&X�"��.$�#9���^E�|��k&r�ub��}�)���6>�f����V[a1��j��\s�]����COp�z������W�v�g����WzV%]���ƨ}>�G)�Ay�\Lc��t�9�_V�ln��P��Jc�Z�6�/�5E#;23�d���.O��W~ZU�z,?$������ܤ��۫d��Bg���9�Z��D��>m\�f�ZqH="Yjۄ]��DL�
�.�Rk��G�lj��� �uP��5)Ś��i)� ����Nz���ףFC>Vx��R�Z礟{F4�\�M�e`�'�����}oOJ$�q��<fɦ9T��/�l%2M��C�W�G�$�T���?Z�=��a�W��_�G�����(aI�K����%������z���#hC8�����1e+w'�y��ފ�v���Z�QXn��af�k�h���� b��@G�v���'e����ĕ� �uL;����3]˳y�{ 1�r)�?�UVY�O䨷Ɇan����&��}i��B+���#���h-�6⠭�w�>�r�2D�V=;�\"u9�M��m���o�-�٢3
�E�J��En���Q�&��*9�S�7�,������G&��.��>ͨގ [:��u�;�	��՛]�!1�F~bm�0xA����,�[��Ҫ�=�Z�'	?��|B��u
`�4��/W�5�X�ǎ�#<�e&�4wj�滮qm��&�nP�N*Sֿ9�_���;�O�e��p��'>}3�y�w %�2P�u�v:�]8}��h�"�z^�I+���	:5�^V�`e�>��r4�n#�OZ#/��A���U���,]�WȠUf��nq�m�]�['7�K���ӡ��LJYq��885S�.w��a�g�t����>T�m5���r��Kb)C3W����r^������OW�<L��z��L|K�S*�@��0MA�^���@���yrA&"�"�U�,ƭ�_�~� I�_��5�N�Ȍ��t	$�cL-߁����W�*��@%����`��D��d�89X���㱄����'�)R���VC�89�ʙr2I�f��1�jZ�p���@b"������{RE](t�YO�w��g�"�zr3����H��ł���}5�5s�:���9�rcR8��C�X.V�c�H��s^���9�\\��[��)z3��6t��"'�ӯ5���-�5�3��J�re�ð�j����w���M��G��*�t�����C+ʛ �wy2G����W����;�K�ψK��YϹW j|�^@B}�e,E�\F�{]V�=��9��s���UN����<��(�ݑ�R���F�"hlR���B�"�!1⼿���Fj(��8�^����.̒Q'�I�k*��M �3a���e�3�?n�K��S�-�:��
~?��J�f�q��$�N��_��z�s����J�R�89�������SM%P�o �wJb:*�$jH�o��7u��/6'��#_����ftI4�i�<�Yr��R�G,{+��$���O.��D�8;��L�v϶�q�WS����ŗx*� 4���a��r����qjN1&օ�K(��b��� łc�|�J�0w�P��"���[7^��H�����B�L��b�mڎ�U��b5o�&$`���M_�[�<����.v��{�%@�N���1�"p�,��S%Qk��cm=6��|Zd��Q&>&`~��6+l�����]���#Ъ"�Q�5�#�ɒ+�;CW��ȭb*�]��:���oM�?̴Oe{vT:ɋߪJ�G֑\"Qsr�P�q~u�1��M�~�����?��l��޻�Qc�r����b�Z\g��筲�lUr�T��+x> �nd.�C�/+���U�w��qw����]u,QsQ�_x�4Ep��׫6T�L�}[$�+@(a�`����\��4�9�֟�]��7���˼ѕV�Iب,.�f�"s��R��/!�d �����x&�����ܰO���bZe��@h��r�5y�Ț�̽!��[@o�uj�8&'��G*SF����=����Y[i��D�x�}�^Ŷ�\���~����)P�g������TϞG����?�:iT�F�wk��^ޡE���lۓ�4\��v��,��v5�\3NL5�9,�|"ǀI)��tI��p��RK�v�c+`���<#� )����־*J�STЧ�^͍�>� :����'�0~T/n�.�Х^����E�� ;Q?����3�A����4Xg��آY�LzKQv�y1�ɋf�ڦ���K!��?��rG�F�ɲoN��^�u�\d�����a�7�����p3jC�!��]z
��>���{�4:j	�c=R��t�z%<j!���V�*>,��f�t�ЌG��@���B�7]�4ۑ9�!�E��ftytх/$�r��o+P�w'��.P�b4Ww����]�(8�P_�[}�J�⨔wR�����#�(^�:_³M�^C��R�¾�ﶪc�{�kʌQ}��N�;����u ~a���@7@��q��=.��e�o6��&�{掚�߱7�;J,,LvI[a��ut�=@��
���BJ>��{��ԳbthI�J��{Hc�s�Lfy��&���cY���8�Y>z��a���
]3�ﰴ[������\Cz����d�˟4¯��Ͽ\!�\-9�6����M�'��Fɇ%Xq���h�☆�D��kj�t�6�[�|:�bt��]_� ��xDHF��G�������U�F��ȱ��"/қ���䐋���#�fC=�爿�͢���vt�l(�r�0�G�;�[��
�o�gӠr�XL�LZ���}���rSme�,W�j�b$�ȝ`��L�aH6"ޱ��`�ا�1h�+��?����R��(�5}����#�p��>� "b#[2�Q*���?�n�������﷌Z�9v�ǜ�38����f?Lc���ԝ���o!,�
$�JPd���wޚ4�趢a�5�"_���dCǑ�1���wi�k�D`N6�Cq����y*�8T���%b�K-(� ���}���4������>^�G�ܴ�t� ��z�T3>�apw]B�\A%���Ft>�شY�W73���	e��_�E��6�b�sy:�X�����z�)�:�yP�ᅋc�d��5Lp���n�_Tڛ����P��48= ϟ�US'&��T!�$-'�L�_���Z�6.b<M���6l.��k�=��3�U}ʝ�~��Z���qQ����&Ѣ��g����q��5J���#k.�-����a��$��3���5׬z˂�[#����F]Ԏ :N&ɑ�%����B}0��o����I��d:�(�Vf�Q��g]�&^m!�����A�C�g�yx��f��'��>�� �B�(§�>ӝ7z�'���������o�U��d���=:/N�`�6[W亗��{yг��Ů
RbaN$y�����Iy0��|e�T��5�LV����C͍؄L�q3\B�=�j܄r\�#3������Y�y�jb� ���<g�*Z����dǽ#�6~��ە���}���t>�PHH����n���H�ƃx�~=[��^@�����w�$��?�.A�l�#7A�X����pYҘb�]�7��7�G�A\{9���l!w�м!P�h]Kg"+s7�������21�r�!	̩^���N%�h#���[�ӗ�{ښ�Ky�-�yG<oy܊�\��͠�H6%���^�@d��\P�+Uu����f�ft�}�BB�o�7�`}>�U~$���=��X�ʚ�� ;�_�3�����q��Mř�������΁���:ۍע%�K�h�`��.yl�ff^�p����#d�˘|�i�����O���VJ@S�U%��d�C��.(4Ld�K�	j,\(�H.{0/g� �im+���B�u$X���F�:xg~�-�X�}?�'%s�~v-?�s�!Ǆ�-����������+�	���w��/��ý�v�d�C��TT�H�	n�'�:�;������_�W\j�>���zL	:����G��������Z*CM��8����p�X�3��sG�B^�����3�2��,ƕ�JX?NnXR�xD¸�u��[h��I�aDio-*�1�Ų����,���د;�����65���O5]�y �pM�9��ڋ��H�<���^G0o�<@
8Վ�," *��wz�.��������4�p��wL1dQz���,�<u]���"��!�x͉����ߨ9V�JS3��O�8_ep�^o.۬��U�h��^��'��Z�J>.�i�I�H��Ұ����TK�nNJM�Ӻ\��.��W�+�uD�a��K��k��.	���§�dBbM�1F��s��^g�3h�'@��9�۪8r�?9M	���kG���a��Q����r@�;g�?����;�jk)��h���iY�
F(]���������,���f��wrb�}���`�$={�8�`EBCP�m-��.���%��U�M�T�{�ݎ���*֛����I��_��b��s'Y3�"�3q�}V��5�h�;������\9�Ra��V��jQ��diP!l� _�Ǳ\�ww��ႍK�����>��2�l�@�C�̻+wU��(���C�|��>�
'��7�+���n�j](��d�lA8<G��z��߶�d�Q��Ƣ�����lν�eIAX�TP��|=��M���"jv�o���`W� O�y�18mYq1�B��Hk��c�����臨��rgx�h:)���x����2ǭ7_h��@���3A�p0���%"��p<�RLQ/��v����ǐ���H�&�P��kn��I����¹=�xv����^��ռ3�՘<!�@����+��;�~{�dt�)ϋ����h��9K'�����9L�m(vw�����v���vva�.*	�g�anqN�b@d9t|���2��T
��EL=4D+L�f��2�wv9'�|(Z�^���W�P��E�����:pS�=��$B��0�����[Y�@���&�8�]��?����Bo>٪�:J��K�$�3"".)��q�f��KN[�K%Dp�<�h�"�@L�b�Y돢��GT�ǘˤa��?{-���x�:S鯒͘&��&�!�W�r����X=�z�S��D~��[T���x'�F�E��QI0���"���C�O)�t?�G���4AF���OΘ
X�*�^;�o�8�	�X��^�/9�#�@բ- ����ĭ��!����Mkk|��\W���f}eD��>p�����::j�8��$�ۜ������ƈ�*�"z�_Ӻ�n]9�G��#I�=��O�k���v1v��Ҹ�Y�+غ���Z���~��b���gDv�hy�,�bK��RΡ�{��U����<n�
�O�Q�k���M��v�I�ܟ�C]��b�|i~#7[}�V���B�1gW��e������Ωљg����,ﮕqz����<�߭)΂��ݖ���X^m#�N��M�[��%� �� �}�_?�#9��ӗ%�E>�WB�n��4�^	>Y�w���N��	�yWo�4r�IT(�C�^���@���)b��<5�MM�`��W� �on2L¤~�/ u����qk�S#��X��tR&<��>����.�ȯd�W	�M��W7X����KP��f�|����=g|T �w�YL�*O�jOD��A�x�s�$ڗ����ځ��9�ܬnS��E?.��-��BtcS���צj�P���<ˮ��u����"�5�k�zpZ{b���{�ɫ�I�o��˲�E(�8������<o��i�����a�p�ײ�^]=�;�Bf��ϘP�'b���C?h��6a�X ��˳*�[���T��S	���B����`9Z����1N8	�1s�]��R�K�f\/�ݐ�̲m�]k���2��ڍp��m�|IA�Jb@���R�MY��y �=��}���4���VU��t�N�'&���1�+��x�,��Y�bc ��w��$������&G�*�6+Ȩ���8�T�B;;d�[OQ�!EHr�ʺn;eDes����u�2[I���0�,���B@�x�m��TW1|�����z��3�����f���T��Qo���� ���5��v#N��%��}� �&;T���c��CƊ\��V�0���Skb�VXA��/z=\yz�_�[�����`�_���1԰�S�W��$�w"=+�%�L��B�1��q)wV>` �
w�A,&����x���^T���EY>����#��-\�4��ňr���1aC�8nᯎ	�5��׎J��$c1T̓�\9�Ψ�1u"�!9/g�$F�L��[��wa��p�'��� Z���NV�̽{���Ю0�^sz��Ӭ�iP����9�
�v�q!�m0WC�v�]N�}*p�&P��y�.��s��f<���glj�L��1�[m�	�60����?c��Q��[���@��g��:P6Y[�P�Z� ��Ne��"׈���BH�MU����w�@�����~S3�x#�oq�@���E�QO��[	XS����1�#�tgS'�S�K��!a��E8'��\��7��P��qv�k� �]�EU�ċ�59��1.�Y鉍�u��Q���'��^��n��(�cG/��.�Ѧ@��N�Yz���/Qݮ�ñ��᩺~#�δ2���Z,8P�E9�֡��.]q���b"����Ӫ1���*5�{U��׳��ϟ�M���d!;˟o���S2z˒�r�6�V_�����کζ�K��b��<��������x����@gZ�x�i�q�,1�Q_�����#��p�?5��n�r$�!�3��;7���q1Ǉ|��T��Sr��%(�ӏU�IlM�Ǐ9b�39��d�c������G8�?\�+�
�.9���Fӧ�ė���5�g����1�m�Wh�^�*-0�����v�\\�0нHP1��7��8�X��a�ƀ,O].q(���Ob�H�)ӓ,~�ݤ�;�
h�P�)�β8;-H�����?��͋3�(���M2�X��mM=�~)�0��ҵ����$"�͎T�>�0[�`W�%�j�����_^T��u��~��Di���8ܖO�"���L�^Dl]�����j�k���2эEp�����J`P���u�7�fF�ǭ0�T ���~� �����0d�����m�r�ع��_����^�� �	
�:�H�<J���n #�)H��������pj��{@r�r���S?\�`�Y"��ҭ�=�7�c@��P[J�?�
�S��-�Ȑ;٫�6���@iw)q�c�ѣ��eN8���2r,,��B���y�4
u�4Ş����Jʡ��I��]3���nݼ�}�"�=������%~#͵�x[Mg�硿�(� �l�6�����ފ�>>������+Ҷ�5�9��U(�э���<��`֫,Sd�#IC�Wx�;�s���iAJ��`��15��`Y�j"�k�E淖�06�V?e,�{0���|*jW�� >���	���)ɕ<M�ۊ-�x~8Y|.�Uqf��%u#w�����y������eQf��R�7�t�	��O���Q1�cڨjt���ˏb����c�.>������
އ�)H�����k�9ЯS���z);D�c���A�5ˌDq���J~�����@��ی<�`�G����zY
�,:;yE�+{�ex\s��NW�k�)n_a�Sd_Et9����_K_�T�{�R�.C��?2�pf���b�c�Ud�����K��}3A��i��̈́>�B�!�20M�4��� ��M�t$�9
����h���ʷDS�>0��]sV%՛���$�a�y���sO�$g�9��Iϒ��W�'ߋeYG��� ��)�G��4R(�P�f�V�E=�l҈�X�(FݛB�@��yQy�x����2����I1j��,�/f"勮UЯdP�E-X;W��л�=ā7,�W���j�/3!h"���ˋ��*�j(O���yVb��qR�<�o�k�����*o�Qi`V��I.s�I�?r:���r���$��7C/��A��%jr�l2�̧�5�?���`~���X摎�x�m������v,fD����E�_�j8Z��R~Oc��R�?O���]�~���L�i*�c�Gqgs2�fv6��-�^E:����i��GuY���^'������.<����S3������X�z�7������Q-CP�;�_
w�m�D`#��
Z��A��e�($P�gV�^�/��a��Ϥa�fɧ�,AΩRJ�2o���&���dM����7v�ĺ�v�Œ�(�;*yؾ�+o�)���p�m���yU3p�x3�P�!Z3�1$�0DUZ��E�Rt�̧��z�U��G�bA"��t�
��q��y�D��Br+�W���]����j�}�2b��D͟^M�+��x^i��̻����5�g�U����������>Of�[��]4�c��5m��M�<����[-�I���(�[x������t
H4�B��(Y�����GitEme��ʠ�������y_]�WF��-�_~	|V�n1�4dfߊPl�J2�(_�=J|?�G���*0S�Ε��#%�Pέ�땠'�� ��ݼ�0��n�
`�O��LDr�B�\�xg�[�5+�5���`�]Hs/-�����ei�ym�K*k��h��|]f�a$$�'�ۆ݀w�p�N�Q�/+L��Q�+2Ժ�7sz�����sY̗~3�S5�`��"�Gr6B6�-wyްn��	X�ϰ(5�[��PϽ`uW��m��f��εN���R�� 0$�);����� 8T��H�ZeN��ߛV���p��e�_��5�l@�(-��0_��JL�ታ@4��r���vO"���&Ը�������t��q�$k�O�UNZ'Ʋ��;���:���Y;�S��+����o(��o��7"��\(�8»��.�����(�������,���NFܗ�l��!�	�������
���f��N�����J+�0����i��#ǌ�(�۱=e��ӳ�Î�`�w�\A��|N��
%����˺�5��G�&l�g���1�����YU9��ZyQ��Z]ǖ���[^+Ʊ�Q9�6S?��
JCf�8�ΰ�<,��1��cO8������CkzbꝄ]�ɺ�߱��dLh��Uf�/Cf4�O��/V�i�h��6��8_� ���]58��\l6V����s/��}�z��!��SJŪ)/l5%	YQC(�,�BxF�'�ۼ�_�����g��7�?i��:���(@�q^��qM�O�o����9�i%���Y����$*;���s���jr�0�z�K*�㗔z	(�~aݓ�b)B�g����ʞ@1�����|��W%5�}�I�����!!{ؾO���껭����2!̛1\7�C��y�j;T&
|Z!�7�"/�i1  `�~�#z��9٨���.�)=|���W1n��q��t�<����׋�>겂4�Er؋է)��}���"O�.���=�.RM.�`���S�}��r�zF\|п�յ�Ok<X�cD+cZ�5�-�Fa�3/��tl�w�<_�:g��Ke9dwacҋ���6�e�r��P�Q]����6��{���2"%}��o4,�f����I��T�|�n%�{��q_�2�r�v纆�=������˃]U>�a�ڹ?��z�z�%�G[�d�j �r[�O�ӑ����4�� CK�Z��$}���$j�"c?~��7���w����&���`���u�g0@��+��HZ{
|�KN��nv낍�[��Bh�n���(dyΧ��+��b���)�Ƃ�� ;`��u�s�O�!M�9�Gd��2����|�>�h3[`ͲX�H�H����m:0�$�<�P,��n#)4��%����whk��J�*|H����M�z�����Ϛŵ��s�K�0��rJ����-��$���q~cA��BsV[�k�	���&�|ː��7,��2�a2RT���q�h#������@j��e�����L���K����~�pn#���}j9]A���P)��9m��I5-Te�At[�pӣ�`:�,b����߅�۱�5��BB����Ą�̻U��԰o����$����8���5Z�$!񠕮��;틂�̴P�4�\ؠ15�~��0�g����-��\�)OҳH�g�
dO�q�P�����F���u�ۓ��$r�${��/7"=r��G��M+ph+VAC�	TlجOj,�-���8��ţ����Ce�a�mEG��ZB"�e��Y��k"��h.�%�Ap�������>i����z6!Q�3���j�H��Bt�z\���Z�o�������Ft�7n~�X]} ��cNWG��
mE�^���G���K�V�C���y��eӅ[�s�j�Z'���Pd-*_m� �fɠ�>�N�&�.�K�:�����̶-_�dNf��E(1�pO���W�$�:"M�_-ܦV��,�ڊ���,�ah�L�d��)J����y=7T�B�XFm<��}�t~3@n
��;L1Ւ}"73��!%C|t���n�5�=N�-�@��}�J�HwXJ@
��xJ�I�~����\�>E�ذ��(���_ۓ&�Ԧs��1vm�Ӣ�b�8�ȉj��>��NXӠ����I27��z��>��;���F�{[�'c��%�,װc�d��^�8�\��N��jIȍ�Q�7�f�r�Z[��+3�6��n�\Lɖ!|̡/d��`���ٯo�g�R�adY ���/l�y��^�,Eƪ��� �&.�l���w^i��w��qrƍ��!z���?���렾�Uh�}�YÞ��v�ުa5��� j���w�ZZ�᥂��B�,b���FS��1�]�F�v� "�U��%�k#Tq	c���%�VN>�L��@��j��RԼ�/����K=�����W����b�kD��WIȰo��c3 *�DL���� ~Jx�Z���˾�£����K��U��m��=O�Yj���$��H�up��;� ����k-:�۞�J�~Z�6�ָT0�xt��EB�d����l�P�K�B��־�~�@^�;s��w��GZ9"3�b��wb�g#��5���x��n���H��.��o3u-��:��ݨ^� �Pw,�����?���b]��\��_zR�>��r����Z��K���7V'��)�'�x��?sή{��T����gC{��t�/n����O窉%N��SSz7݆5��Z-P�+�j@�C������A���38:��n�`ʬ��c!^\.;�>�˦S�P��8��*��d�<@�Fq�N�qzj��OaZ$Bq���,4�EV�]��ӗя�i�:�p��٩M���J?��A�zzU�������{�|�>�ǜ>v�V�����A !^|yU��0�ʲ�y�gv����^Ӳ�������.2DK���K�Fۏbo�>4�?�
+���u��G�?a\�@�""�)�O��o%��}1v��,����ؕ\�a�8��s���B�+ �3U�)Ġڥj`u(ԩ�| đ��|D��1��u��1I f�l���,�������zp��+ǒ��?
����K:VYAC7b$��F����]L��Wf���~��Ӿ��|F~_����!/�����z���<ٝM	y�m"�JeG�B()� `nw�7;@���.dЦJCv������8�幎mg���Uz��|0�|�wD�]�$�6OJ����dR=uϏ�ha���a4���0M�/�Z ��A>@H^K�5hvPU�\\bv��BA�O����V�e)��*�����m���T�|���N�A@�]Ē���|������û���iƱ�5U�O�x��=N�Kα�l5�K;������:��<s�HN��=[��\�2ɉ��Ŕd*t�������U��o�����c�3d��Jv{)���e�xY��^�I�{���ӡ�V�u��wCf<�M����0/r;3��~�·��j�n�r-�n����X�ذ����۵P���t�6��W��~4Ŭ�x��*F9w��0~�;����Fs�d�49�spC ?�<�ߤ��%��`~ۗjg&�C`k=��eӓ_�[�@�!>�ť��d���K<|b��y�h#3ӵu�~�����(����Fg���`�Q�1��� /0<�׽�߭�4��K��B�`�Ng�_}>F��/��!�Kq�$�+at�]N����v흺-؎���^���┙��7�#�
�!��06x��oG?B�3=��oyE6���/Kv�	�Œ9��3qc��R�d*�U0~�f�U�|��]��N���L��;�*h:-$I�b�� ���
�/�d���I����UI��@ uk �M��� Jrzȟ�p� �E%:��K�G��Z��M�X�_+�U��[����9*����42df�D�9��[�K�Mڵ�c퉔���/
��ƿ`1f+}�3�O�*~��p}G7ع���<c �鏪m;t~�����pj=�mU̚�����U/�v���}I.�I�>�B�������w�s��=���9�(6^Mv�1���#�鋲������/�tf�L5�LM�҄��5���."�M��0�Y�~�Gz�S�1��,�[�Gr����U[�#��
��q����� q�]������L6f���a(!r��AX�Y%�>�-�7s�:,G��?*�븛P�xGK�O�=U�,4i�!E���<����h���kO�`��\�� /mֹ�B0ٯ��
-��kJ{q�ru�YtVSӨ](X cO(���$��`"�� (ZqЇ,�$1trk!�5H� ��C�=-�D���f�"<��V��u�}�(�y$F�=W���H,�td�.2�
���c�=��є��i�6Ϥ`fiuܲ��g8�p]z-f��O�w�k�Ay�a�V��F�0D��(Tϲk]{���(�����J��s��`kN��QS�W�d�c��%2��K�55?����J����#�tZ��[�V�����,Q��gd�9�N�ԡ�7���LV �o�sm�z�w`�;Q;���2wa���REɿ�9��>�"ӹ]��b� .�AE$������]�/E�s��km}b`�k�gI�l��Ac�Nk s)2�ټ��R}\��f��O�d���^�׊o��}�����7gPߩX���l`�=�k��F7TNd�L���tUi�ԩR�w���r��b5�B���h_��jj��E�
�~���B���Z~�_D��	����	~}�A�������m����;?z�S�&my���s�������4D�+ xa?����1�����V0�"��|Փ��}������~��b��v,R��}�訨�c���;��=�<�E�bl���ZA�5ͭ�F�b��d����j�z�(`�d����\5��wRT�nk�hfG.��B!����itE����v�r6�悇Z�v�ݐ:g�l��;��dp�F�4���I�#˗�����͠�
N�_��gq�o�0�Z��y��O�����;+ܴp|�`-[H���bjP��Y	�T�r�j��c������H¤��Z��V�u����>L�\S^7b6tvz�7m+�F[,>-��;���9� p�3���N*�$`[i�J`�D�n�v���`ohH�BB ���o���F(�`q���r�iz��?�����y���ﻪӫZ �2��$�4JJ�:��?�"�`e�4�����Ŷ���N^n�����2�񗵻�^���CशV-@�#T%��k�ܔ|�Fe�j�n��^���T�w� �R��Jl�fQIk�
�����~.� �}x~c�k������ي}���"�rMf�<�7����tӝ�g�%����uR�/"J����=�n,�k��/�,ⓡ3��b��K[��:��|��<���Dy��!�^����$�2.{k��YXk��V,:����-�O�8��+c� �7�^^۴IN�}J(��*�5��<�/�C��$o��I��Z`�8'�w&�s�+r�40�j�Lh�=$8eOϣ���:���̚`�E�W͐�v���ۅ��B_�T��.�Y2|#�p�E�y���?Ó �e()-
��e�g��X���z0;ڍ�W`�H`q�R;�=B6�⎅fӌ�_����wU���0ն�������|����.6��QS����|�c�)�= �GA}�g�5Xm7��F>@l#a0,���@�2.�A�qFj���6�I�m;�!�W�<�飭��u8=={�fB�2����zP��Z9�z+�z/����s����#&�o8�fH�����L% gd?\�3OB߸\�Z��R!#��Lj��b�
�t�&-�yw�ĆW�l�:z�����!�ǭ,�k���Ć�!���E���K��6��ƪ�ݧ��;,$e��$���r���N�%��F�DH��&�S{�XtJʄ�5l\$Uȥ��#��Ν�H3�M�>ooYyR�U�GT5��+�j�uPYd?&��d��@�������)�j�V���q�5|�Y���]�f>2Lg���:Z���t�a_\�U����E�9ʐVE��Q9t���S��
 �|k�p�rzV�>���j��5;�2ҝ�+���Nڸ�>�����i+�=qn�2�3|2H�qgiWW(�cj�w�R;V�'�8`W>�,�2I��y%!^���?��� ���qdCM�Jz�{��*�k��#r'DBO���CL�	v6QGo>׌0K���Q���i5����N���+Se�?���3ݓ�� e�A�J�`�
�}��c\w0=Zvh�m9����+i�Q�n���8�����f�$�P��W��@\�^B�i'`�Mb_�݆3f��T`�fڶ a7t˪�#����|���I��4���,r�h�{�JVߖ�`���^�-��j�KsT�g&�CK����3Ü���~��`�'`VOv ���V �����t���bQ'F���ө��� [�K�p'�(c�q��{��U����٤_����SD�h�5��4g4�5��`Υ,���:>����m���"X�.�|��J�w£9�=/YX�3n�Z&}9�ܭ���:$��:g̪%�"?�%1<�N�9,��N��z[�����C�qVb>i՝6f)Ş�3��"zC:Iŕ�F�2���Cz���	_��������/��)~H;@�����l ���`�U�\йFd!_d$t�3{����8ݛ��|����?l-֣�.��=B&���)Tӟ��]�4_�0�,��|�X��E�[�~C��QIo֎/:#ɫ8ti�v���#6�l�$�K&m���ȥ�lf3��� �
���N2���aҨ#�l�I]Pj�/n�B���)�5����J�i\��AJO��!1 R��I<F1𬷫��v�Ĥ)���mk"/?��ʟ�|zQ��2�	1ַL�y`�|����Z��l+9�m�ol�K�<��׈؏�3��Ђ?��| =- �������	���H@,���>f�)BJ�+�p0�I��4��~�5�景�ʙ.e���\�(�?�L�<~z�Ot\-�3�%��TB��xdI�O�v]@��w��v���MMvF��5u�̭��<۪ߟ�RE#�����s��Vy�d����ĵI���3HR�v1������X���B�w��fK�d��<A�����-�fa�� ���H:s6�>�:VΛL��: ���_֔�pfu�s���q�DR�Do0y㺱�Q�* i��T���4/�0��~�����k:|�_3G�fĉ��쒱�pm\��/
R�^{�#�D'����\���4���n裇�~��OCU.��V�����ܺ���+��w�^�f�kS�tB�k׽$q'���~�l�%�կ�sn�c0�Y0��2�((W�6ǣ(���e:�]n��/�����%1�sB�$��C��(��q m��Ѿ��u��).#z{ߞ���ρ�۴�"b�ּU��f��ǉ	�A�[N��y�v���=I"Q��Ɠ4�\���M���$_������)�R�_9�J����s�H��HB0�z���%�:����Z�߬%�P;I�m3��{i(�Z���9��`�|m�����g�Es�� ���b���X�+��>֩�ڥ���BT�3�(�Z&C��j}Xt �X��bG[�bg	8/���>5�}�`�V/�SW�RGy%i�<�u���� �Ha�R� �����դ���;��O?w�M�e�>*��D��נ:PsV?�Z�`ri1��ՔP���C^�B�t��˹y1(���{�h���۴n����f&x7���TX��_�V&�?Q��^�)���?�}�ÄJ�y��&B�b� ��B�?�n����m��ϋ�^
~j�:�$�,�am}w�?wڕH}t�]e��LA�	m횕��~��
��EKFx��Q�2F]q�kȁc����c����ߣPxs�r4�x��
�����7�+�d�B������Om�Jc__�8�����{袈*����'*�G	0
�P�e0�J�lO����N>�(��o'���C���4pWJg������7K+WWi�m��������ݼ�8� .�U�����Zo��b��~?�cy�c �W{�M���70�Pw���{zPz����[���M����2�L��_)/���`��I�Ө_I�+��*CSiyS���t�R���`�������6��>
Y�mmVd�����l,d鱘�q�=9n��b"�Q�SY6��3����u�J�x^S��|aZ�Bꝳ�FX�D�*�����I�y�ݮQN��u�$ͺ\]� ��u~�w��T�i�T�����l�o���پ~�����M��uu�-��UAB�a�Q�6ѥ��W���b3Z+^�.�4���*�o*�2O�\6zR�:a�1�u���ᄸ��oVrC]F@��*��C$Z�����-���U��J04��2<��E�  �:��M2|�_�ms��À�ݝ`Gǘ�����o�E�X��@A��lC~��=�.�(4��J;U������ �1J�>�=�ĚԂ5���#�'<��p��d�͛�.R˹�oo�
ÅG�ѡn�E�Q��QT>�ғ{Ʒӓ����Tx��t��9��&F~X�����I�	bI��G�8�Z+C�<R��V.�l� �Yh�=�/��{���NR~�Q9T ��g��S�V�1��8�+ i�$^�4���޿+���[ך]����Z !׹-��"�:�g��8�?e���E�Hybr�8����O&�2���ZvM��~���]jĠ�噜.AT��%D�*��J�ׇ߿����B�w�ЭSM��� 	ty���@[Z
��<���B0�s�B��=a��2@0��\7���Ȼd�[����_9	s����Ѓ��� �޽Mu=���R�}!_ʱ�<$ZxP|T۱�wh]�XhܒS ���θ��(�݃ MOې0$�K��=�hgf7P\9���2*C���)��g�f����o�1����\���
����a��Kgo������Z�<�ENo)�? �e�������!<S�7 #�BI@Ɔ\9�~b�iG���"�����ޝ���;aͣ�����!��M�y�6ǲ`5�7��W������(A�2쭙 �5{��!#x�o���d��B%0��F��U������N2��(E溱"��.r������P�J5�O���`�u�9��L<�eTߘ�F��BM���k5��x�z͍�Q��˂).JH__`�vG7w�ob��n��Xq��j�Q�(ƛ梭��Z��C?C�����|\s�a<��a���("~
� ;A���Ub_�Qaķ� �n0i��bq�b^�_��!p���ZGw0
��9_���e����=O�V8v_b��K Z!5�š=�y^X�;)���L�y ��9�?�R��*U��,�b��&���3F�&\\ӭ�
��HӦ<�T ~�Y�
�(�Pgӧ��>�_܎�%Ă�����I&=J�lD���H����S������c��0uQ�Y1�?�-��SM�	�Ԙ��N��)R1��fI!��Ve(=��I�F�s$�Y�ͻ��3D�d����B���v8}�W����	B�y��DnÅé�A:��m|(�۵�v���n��Y�j�OzѴ��l˔���w�0�N�f۔N1t��gÇݗ\#�e�5����>��T�I��9�}*9�>�3��.(ώ�\�R��/+{9(�g9#sn,�l�(e4
v�f9U�tQ���te�1�5;��3�����q��`v�uN�@q�[i�Y�b�6%2����r�H��i���� ���j��;�n��C��DU�f�O���s��Vr�ȣ��X�ד_�`юP����^��x��
����|z4����qf.�x�I�t>{���筕%,�D1���V��J�b[r�1)���9�h^���a��EB�w� ��y;��c����Ls�qd��o���x��e6���am>t4�����)�'���^.RT�v�����\���M4��o���&34DL�.">e�0XB��NB��S�`�7�I�vT�/C;���W�<p�R/yP�cj��\�dNH0Vs��:�Ħ�=F�FbV����udj�������0,W����C+��571I�	v��7p�p��'[���}O����ZW>,��Ӆ���(`�2��k7���3��}�0 f�����?�;��~;$m����n�P1�x�����L�_O�Z6�����L9Ҷ����2�r5Z�yz?�Ӷ���%�	��V�CӼ�@N��f�o�7�+@�0�(���5�Z�d�Nh��=��@�9��� �:�W$�y�qoo�o��+>�'��`�gL&�U `�~L7tP[�q��ݑh	��a2\��%B�^�������uy&�s����7ɠ�Vҧ�&� y|,�����:<m�e�l��_���NnP��]Jd����<��"���YB^�cn(n�3PW�/>>�'��C7	I�<X>PZ)we�,@KQ�N,� "C�B�?�������Cyj>y�WO ����2��~;��7�E<��CԋK�k~�~�߭�r'{��J���/%�>�Y�M�`�����skM�T|7� u`q���sԁWѿ`i�5�M�	ғ�R��+�L��d��ݯ_��j�r���x�����o>��g5��*�y�W� s��scӎ���7�����}kU]��C
2<�.�1"i�MiO�y>�����{��y7Z��!�/Z�߉�G\W���oz�U�p��hI,q3{����h��e"3IX�V�fh6�n�e2�Ex���
/�,?�gFK*�SK�jP` �N7rж+���"��W?��nD՛��$�c�����0As���C����K��.^�B�[[n�,��V����q��m��54�����r�ɑ��0��nF�6���u|ң�����JxAۯĹ��cl��`���˦W���ȩn�j^I�*KD���>3�~�X�T�؟�\��u�,���ct���y��r+8��L�b��� ����.�"������4�K-�p����}..:�Q���0����f��e܆�,Ԃ�~>:3+�&�f�n���P�)�kzT �a�i�z&cxˣxYoR9P/e�+9��� ��&H��[pՑ�n8w�@�Fj´fX��ȄV��(���X���ē�?���;�*Ns�z�e��%s�q�5�r��l�o��#!m�Ȉ	��<��`�_ֻ�b��Q�ދQ�]�.�*���k11b�Miw_��6mn��ۇ�� �z�E3�z�[�
]ioQ^��C	?;��C�Ԣw��lH�C�{����c+X�����YE�����ȯ<>ۦ��a�Ձbb�?Hv��U0X�}�Y��1M�g#=MT�+�oW���-'���5� ��:0�����0p�n�~�
Q����hq��,uk�d�D˱�;�w������������d�_��4q���[Â>��1�I������@�������qo��ɸB%��LJ��[g�=�� ^�y�ی]�/��d�jjs��j��jқ������6F��"��N�	����n����b�FQ�sYf���M�k�(G�����t�r(<|�ġ��%
�J~CWI���TVYwPǷ�jeg�mF��am=�n�$N�6�O�7�Ƚ��N/#����ɀv�QG��m+��u�-��i���K����T�M�Eԍ���b�WKP+/9�$��X��>7��	���,ę_�M��PlUYx���<P�D�M �U��-[�E����]r�@��_L�槊Ď��ue[���ū��81�TPBs�(�XL���.��ʬ_���?��M]�sH.H��E^�|�s+o��d�1�fO��v�r�h{AT�T��j���7&!7{){���<� b��*�K�3�-���I�p�n��Oua��c?�u�)H���C��pk3�f��̨dB����D7�ptt	��x�BCi0�E����[>�Fk|�����Ef,Pސ��ʔl�ۙ��Y�� �D��tQ��;���y��$W�>����im�JO��2LT��(�P*�ܣ�Q�h�"��r�]�ˑ�ɻf�u/�@M�A�ݿf�t<���
�@���L��n���gچUY���������7�@|�����ξ��a�VT�n��3�a����=0u{BK1I���-�x�e��=+��S S�Ou��5�%X�4� ވ�xG�A'���4��5[��?�ڣa���}�fy������5)%Õ��3��~Ӎ�����ܩ��tX���&c]�?��f<k���~��t�X]X6�1ʻWVӛ�=�({ Bԍ��`Y�?��v�ż��,��׬��a�g�z�7��QJ�rnG�-$ˡA��퀭�Gmpr^ʹ���gy"~��cgr�{~�0&	��8lT�hx|�ï�|Yn��0hT-��L?Mq��&��<�ZN͍��Z�G���d��h�8T�C�]�4nb��u�/o	H��5C6r�.	���aGqj�z1n�qkr�l�@loXŢ����ZQ�؂<t1+{��)ԙ]��� �B:�&ĭ�w� ,�%�̆�	�"�-��<���T4��s�[�X:�Tb�H�0uڸ�8;]|�&��G���T���P�0�7����s:eL��$[E
V�������e�� c�g&�8Z������w�TmLR����U���t��Q˖���3���_�4�ci�@�x�L�Y�O�����u�~���&M���_�^:��g	�]�W��5�����
��W(�Ş�Šk�h9��~��Pl��f���R*Z��o�x��8���(�P��7�����`|�tٜ�à`�T#�ś��y]��JY<�L����9�=�t_�˨&�<hQA�h��|���n�+�rl;����q��ȍ� ���R�J.G�{y��k���^@_�s�bu0S	���0�I��W`��V�~���� �Xs�
�0������*%%�I�\�����V�F�sj�Ζn�dtŏ�n:��W��2Z,-uq{�(p����Ge>���ݻ�EI|���X�����si�����:�+2?�:��;��ׄ<������7��Ut�q3x����rQ�Q�c����[.�_M�HQ7���`�đ���P�P:s{�n���8l�/5� �;�_*�\��_z�=�����묅1�c��ԝ�qx}�j�����4�e�5�{[�0qy�G@)!H�2��/���Kv��	 �J0,�k�����4��r���@��YN�n����_��\��'�K�z_��������"�1�������P�Ԯ��in	OG��"����T^�D��g?Mi1���6>��۩�B�,O/�?Q���:f�wO��BI�&ؘy\z�6P��Kcr?��/�6��$@�7��B��ps�m��H��>�鼄��+��H^��McoB���Bt{�	�U!0ƾ�c��g��2����1'Kj0�`3�n0��Sm��]�o�0�5+��R ��;Iw;�gZ.��1B��^��1?NxcC�(�A��1���T�;�$h6�+������Θ]�)0)t�M�n�5sie�؟�#՚��"R�˚p���7�z� ���&�#hg.��WeR�]������V��H��x�J+���i�HZ����'�x4q���{ǽJk��P���ju�mͅ�����@�`���*�8p�h��<�n��#%́<���x���>�����Tw��¤��惞�P�����u��Y��p]4
�)�s����LϜ�E����,�	��uۮ�{������Z�u���
�|�c�=��u�WH:\@�?RQ��dG�r������wX�N��wi��c..�:0�TD��O�^ZFYmVt{�Ƿ`���N�g\���*�n�┶�dBZu�3qa����. d`�:+&8�2)�ۡ�=2x=��vu�����68?�!lҡ�X@{�"qQo"��H�U���mL���g�M��x�g�&ݍ{�=��9E��AV�CM�2u��|%�@P�|�H���4p��k�1�[3�h���Y�����O���l@����m��)�S��IL��f\�K�Q��W�P6L��U����GP˔��e�����񧟒0�|+������ w�bH� ��� LF ��i@f#j/�o��
���y�C�6L�I��J�����a�wb-ߖ��A�AK�p�v�CB|�Sb��]�m�G��̙�
Ay�ـ��Ǣ���6�f�q\b�A)Ix�����=}v�U�E�G����>&�r
�/�f�Bڃ�O�ɷ2Ű�@q�Z�eO0�1.�Y��*���Ә[T�~)I� {�u�'I;fkCT��j`��V��7�2c�1�p�?�C?�`*��R?\|�.�57M,)0�K��aj��H�A�Qm�R����t�2D��M���m�Sv 8Gf�L�,i��sa�LdQG�V������R6��j�:9C��V���0�gL�ږl0�oƣv0��( !TdC٧ǴI<�#'~�ݫ��D�ŵK^$Ȉ\៷��8R���c�w�b,,��[lFP�\�3�)�C��2r�q��&b�^�����'��Be]6�°D��Jc9�;���5͸s����]R`�^�<���%�6`��۞{���O�Y+���j ���I����I.>�L�e���c�\��)ܘ1�3h_��R�<Y5����숰��[H���^k囆��>m���%��6�� F�>���P ��I�4��{���{FD�.�G����|q����ҥ�;��&��(/���NVi���"���Y�.J��T*eV��#N#�W�px%�WX�@;3hu�W�:�}!'A�l��)�Ч��S���Ծ������Q`�G�>1H���{���/��������<a��}{)�'�c�<�|v�D.��mu�z����G�"����n���dt�0��k����_��Y�#��KoC���%(��OKW�����lF�#?�,��XH�Q�B��J� �J��i�?���c�Y[]�����X'2�Q����XU~6G�0�m�5����ǰ&�����Nu�#� �%,ƎjB�QӴ��<GGR��עY�a^���cO<dm�v���9�*��%�52ᄜkC-
)��>H��x�d�w�.=��k�����B%������]�O�zǁ<����/$�a�#0130Ϲ��r�T�f�lug�j0�G6�?E��hp�0�?��!�щ�k^p��֙��p"� �TT���'��6B�Ն�$N��j<a6>?L� or"i�H[���-��#Č��Y%�Ux�K?֭���<��Ks�n�-����<�F/�]�#�����&H�$f&��ӈ"CF��_�5��4�B��`�RF1q��^�&{�����5�Hˢ=���N�uiT�*��ې�����κ���E��6�=�w�ʽ�=t�?����e����#����u~��~�YJ]a�o։��x�z�x)�̡P�w�hdO�M�� v��SA��˕�aĜeN����N�h�	B�FF���>Ď�B��I��!�
b����b�>�س{�(�NJ�+�OI[��,;K�\X��N۹����uH9�p��jJq��������ՐA�A�KO�$��̤�W��Z��RӖ��R^.����'}L$!���������b��r'�raG�i|��-�<+�.@���%Oh`����&yH�a�	,�t�!�����8J��C�h*�v$�z�^{��i��&M��e����'e���X��5�H'-��]���tl)=w�H'�c�]��=f�����9���q�%���S���PaO�Ed�����L+Z|!�W!S4xr �Rdv�-�rw�y�G��H�j[h!U�1�9�C�)��C��� ȥ�2��9��|'�����g2��*-O{�r2cr.���|�2��ȞK�܃�I��]�U����"B��Q'���Q����Є���mx���{@��t\s�g����Q���Q������xyF3�+.�x��5$��"�4z�١s�O�O>J��w�VeWBA��p��{=N��_��+G����w�����,PMN����j����U����yê�A�Kg��J�����zXm�}$���7��T����7w��.���c��n����k&
�괜=yٺ�s��	���`����CI��j��v�9�ȹ�q΂�ۻq���	+)�9�t�@������(��>O���?|8'����D.��O-�Q�w4�����(Y���������K0�?���Ö�w<)� �_#�vT-t�z:��,tN�TMT�'n�3Г,����q���𼏴�)�IѬ$�@���y2���JØ�~o����p`�+M�l���,D�� \:�Ɏd{6�怃��fD�T����\���Ӹ��ӄ�e5mZ!����?X��ڂk@�F���6@��9m���Tm�d���a�Ɗ�-�i���Q�Caޣ.����Ƿq�BT�9}�-���r�?����)��z���jzw�����i�9�l��,����-�+�Ʈu�*E���lZ�r��j��jr�v���uQ��Xoȿ��p��a.Ҵ�� U�)��#�B�3a���-��0�h���t� Rq�-h�@A�JN9{z�{���=@�{ H.��
�R*�=ۻ��p�B��A�C8ͼ\�D��G��̳{g
:n�k�����gǝ%�u��p�'b�?��QMp ���B�8��}��	�C������n�01�v�����<�j�^�4�ʝS 釦��9��~�ܖX�Q�+�0��ܖu#���*������0�'{�F�:)�����7\��kd��N�jic�`�>W&��:xZ�FuUV���B�i��.�(�u;o֊3�=�-uƘL���jk߿),y�R%Ʊ�ed��#�������wtV��t���8i������$E�c�Uqd]d�"�D�3z�<�ԩI�y�>_�)ڨ���=�]�2Mt�i��K\�A���r����'��r�Ә&�͉!G��@>�.��~o��v�چ<����^:�ˊ�(n���q�/�Ӑ���B��mk��%[[��Z��9�������GiA(�E��B��W6��K����H~��?��w�����!Ǔ"bx��2�ŷ��9Bf��AG�O�7�c�I����U<|�������RC~R7���PD�DS���Sܛ�Ʈ,��1��Л�RP�j$�!��y����� 'A���
E��.��3��BQ����_����V��?O�K�D��J)�у�������C�; }�R��!bG{��ouOh���(�-a5��5�����X��-�~�K٧*���h<*�=j�i�4\x6F@��B/L<��>�;(&&�����Z��ֶ�����.�V���3	E��m*����n���n*�H�m���h��C0O���)�WKX{d|�����;���n�W`l�Q�'�PLROҊ%�Y�y��<6�b��l��|�x��ψ/�MޚnU͌I+�R�NφMߌ�wY��
�x����%����"���j,��ӆ�#7� �:�(p�8�ȷ�y�b������:!Qm��f�����T'���9����㯜xF1ZKl��O��J�u���{@�ǰ�gP� �c�$JDe��f~`_`Q ټ�\�La)���vNk�@���GA�e���q�<����d�,�(��'7���\N��ΌS{K��?i?3.����"��[v0�����%a�T��c`�<���]Y��a���J��O&M~�~S�����t�����6og�Q����0m�x|B,V��ҷC?�[�+wt�ך� (&��lV�9	!�o�qqR ZLͷ�)�S6����>���F�z:�� 3%�e��yA�k�������4&�#�`�+��XW�B��#J[��)̠f�����9�/o����|�ƴ�8>���:]p�n�c��ű�8v:\?&�A� bWk�1��G�urUT��$d�r�̚���9���,	ы �)���8V���* sؑG�h�J�84�+O�Iv'�$�գ���#�����`���$��t  �Y,�	}��\5�6��܎LY��nn"�ĭ:�}?v�dUG�6A�8���|�1�7�����'&c�{��\mK�`�8��BnŮ^lk����`��~�5g��hU"g$�r.lηQ�h3�"�N��!��-BD���V+�	�~� �Ir��X慎(�s�Ќ�2��$�%0���^%I��z�6�ܾ�l� Ȍq���'0ݎW�\ma�.��`�H�3
�Z�\�0D{�D����R�G��������Q������\�������?KM�Z��qE�01�e�jdč6�4C6,U1���u[�%�}��뺌w1�2;�Ŀ�x[���?\]��8M1O�e�C��SZ
�uI�5M�p�J;��J��6�P�L�CF�We�qb�8L.�mC�Kmi��PY�����ubb¡�Kk�b���Q]��d�{��u�uր�i��
�4e���Ɣ���e�Dg�6�)�ۅ��5�Y�c�'ҵ "��p�8j#�)и9���8=�w�u��ޠ��|�zK�k���-����=�%錹��r_j�K;Ά"��Yʒ��=ưBnA�g��0�����[ڝA�D�����W�B�k��
�X��0���#x����)�2G�~~�"�B��g����F��\VQ�q�BDz5�~�Y�LY�w'�p��g�{U&�Qx���b�A���A��p�Cr�Ag��3����O$U_���x����տ�{�Jc����N':������-�{L���l�������q�ڑ�G��`�U2�K�.LO��!{���H-\��r��JKY�����L�r���?�������Pm�w�E�SvKa"�j{�����[��������hN�h���.n�y�nf�r���_5%�n�|�y�H*C�^�T��T~j�L�Q�i��+�h�/9�B �!&n��n��H"PM-���a��B�q�������$4��7(�JT�`���BxM>xg��s���ꐀk��X��O���ni-F��̸.�T�l���h�ZH�5ܹM�����ry^���*`�n�?�/0���4�|j��#}d���oV��M�Z(�����W�z�%νbU|sΜ�`8 .u���0�7�������G�qE���7�(d�FvX�[]$�������
�P�W�{�f�T���&3Dlv��|Z�t��D�J	��`�w�ݷl�������=T��*q�T+i��������{h�|���z١��"үƷ��C��4[��UA�uq�H�!��I	}�PX1B&�i���Dy)g�j��n�:�ˍF�E�L.k�c����>�M-kbN+��9��vI�+�e^�m���\OD���L;�,�Tθ(
b}	[�&#��	���|Ϙ��R?5`|���<�k��I�J� YI$1u���i��I��欺�0� �3Kn���8��� �΄O4�DNj_��H^ùH� =ACu����*��]���d���d�,�m��#Z�Jkc	�z��PC?y��m��y�e�Gx�$�Ѥ|j|�0!ff�4� ^�|:�)��D�{d�%�ė���b8rw����](�>L���G��:���TϨ�D_Ssi�H��F�$��Gi�k
��3��W:��!{l�t��P���\�cLfF���✩`�z��pA���#�(�����w��b����Ԣ��GH�=1�}I����W������2�qgc���b(7y%F˭��|۞���9�"-�a�"�'L9�Ja<���
�l�ې#�b��2i�݀���W�[��gO[RK7��n�����N�gC�I���T:)�e	�%d"ǉ�P@Ewx<����@��k���}B�0���W㫩�zA��cQ�n�V��9�f�������©��4�y�4'} �Ȅ( �(#�y9�[��F����0��Z$����:uPעT���Z<+�1����%�� ;��*�bi3������>���~[aM�+���/Us�wq����5S��-��I��N_35���%7g��t6ݿ.^l�"�0��=��u;���AyP�՝vWw7�L����ҁ�G� ��F�y��9A2�/і��23(AU"5�"A[�*��0�p#B)n!!H,�Fl[�����@�uXj8}�d�$c�=#�TcZ�)٘��MZ�lS܈ _��PT�AO�xa|�t��Z^�}��0��W[X/]���s��}Cc��7�$�[�VD}F����䜸ۖ��5|n*Mҏj�])��r�m+pgR��rߪ����q��u�+z�u�_s��Ms�F��C��X�j)Ce�갎�M�fY≱Ka���:����^���$���b/�����J�"�7\��@A�R�?� L3��u��X�a���cC�7 ���i����=��uȑ�
�o���\�)������ΐ�el+Ryj���/�T�*����	������=#���E*%�k��V뚓l�;����j����U��һ��(��`�_"���Ǹ`���p����ZôRlgh���firzo�s���A�\��ьVk�������r�ᗃT`�����<.��G�R�G�i�j,���h�Z?�y���.��A\ħ�����	�%;fh�N�6=<�K�1%�ރ)no%_CR�#]�X�6��e�P�����{����Qf�򻤵�1�`��)Ж\���I��� `W���J�2J�� �6��LT��yN�F��t���x4�ǇP}>��S�������~�4�4�)c>��d0����Zo�9���1��FD��7D���mğ#I��poH�֡������iV��u�n��0�O�Њ\}��aq�=5~NJ������cD��8�HG���������K���OP����xkd�+Jː��M�����s�7�~<Jz�M�zT�6Z��p	mͲ-��B�>��gՋE������:NLם�[ �X}���P�\Z�U��C�`��M� �w{u$T�e��AYF�/�/�M0��1�l�v�@��h�	�a<m�d5Ͳlq�O�z�g�u
�RQ����À`-����!l��RlE� �+�S$��|x�O2�!cy�1~���*���BN�﵎��*�Cƶ��"�W��h�����_�Ǎt��E���̻�,>�`�[�<���	,>R2�vr������i1�=P4����Ff���9l�99_�����-����V~�"x��4�Ŷ�K��k�E&7*�T���U����=d�Ƀw���G�䖞���Hk�1�� H�����	��&���ȂP��ϱ���y\�F���C$BUro�?���t\�F�I1$5�n�1�~��/���`l���"6��ɢp]�g^�O��x��h�CCLL���9�R|����zǇ�X�t�`'��Vo5�-��F�ߒ�H뵉x-͈�%�̴xbA���i5�����z����P��߷y_7�'UTT�7>��%m:SJ�IB4��%�Y��W��J��z����s���ܺ��ޚKF7	Q�������vV�ts��o�p�>�3d���820f��@~��������$�k�
 ��L��L%�kr�	ȵ�L�y2�5jJ�P�AjW�q�)W����i�CY:V.�O��i���}y���W��˂?;y��\/� s*P��z����{@�.��08`Nd��"V��9n��B)[��'/��_6?X+��K|�'��0{��J�Y��΍{h~y� qsh^�Q7�8fT�D��Y��)L���i7�A��u������&��l��}��0��O;kP磶�b�j�w�^�i)�5�P!�1Ʊ��S��[�B���!S�7���8��p^8Ўa�x0H!d���S�ͺ6r�cP���> 7�L��g&��G~��	�{�����V�Ġ9X3O���{�ͻiO�Z��hԴ���**Y�,����+U�[��z�O�C�aڷR�HhF���_n�'j���T;����/B�+�$mOwB��8+K�'�Mo�6���.�̹nT���2'�,8��𩤶�\a��-�F"�z�t�_������P�P� ��9�Y�J0�\���/���U��ͦ��s�Z���Q��hR ϓ�#�^eQ��0�
���	c��,�x�`�����4UqD]�n�g(�dd�:����z�l>�9�O	���qq���g)�7G[�dE�c�a% 
�2�	#^b@b���'�X��=�Y��C)|u�ϗ�+��JB���6��­d�T�]��'b5hԘ,��3����93*4���&vM\�3�C�]�te�.-�d��6FS&��~�>"i����]mJ���վ�$�����R�MR���D:��@ր�1��|���c�}�@��rP�=�*�/��߮5˷e�􀣇ĒNr���� )��}��U���9Y�"�$��	-S��6����q��W�N���=�}t' �w�%&۔]�H�rӹ�6�4'����'a;�3�dIG!	6':�9�|�F��ǭ����Y��MA2��7d�a������
�bEi�Z���~K�A�W�<\haLxT��7���q��G��z;)����qFK �3l�3@�ܰ�*�B5^\������|"��?bb�f��m��Β���|fό�5�bM��aW2:q,SH�ݒ��sմ��^!"�2\%B]�ĥO����BC:�z ���/cK���S�Xt^�M@	d�s��[�z�W垊d6q���PIe��u�:DT��X�m�F_Y���>�J����{����cH"��y�� [|E�hA�M% "&��u��zZ�Uy�	��E�g��o����*�Ã#�7S%k�Ң
>T�w��ws�}��6��U.o�������L��]�c�\,�	13ھ����B���$�}�d�(��궱��{F�7%� 3�H�]�}�h�J��&ɵҙ�U=�u�KF�?�E�b����G���L�q�g2o�f�+J�:�^��?���f|U��N����׸���m��FG���ִ���P)��8��B>Cd�)�|}�]b�����o|�	���Arټ8�W݀�u��\� �eR}�Zz��GE@>�m~#k;<�����PJO�{��o�A�����:���G�= �'�/���$ ��E]�%^m���*)KAxE�<��S�ι� 2v�,e:�\;��j����r:�
@�}�8=5F8-5�j�'iǳ�x~���{kuAU�-K9����SG\�,��IU����U%�^��N ��ڟ�����{�7�B�u�A���A�ʀ�
Ǔ�<M`Ou��m�̹��9F�@o�����,P�/я�_
:��Έ��q��c�|��hh�Md:�,Q�(�+20��b�@�,>	�BQlz�nf�s�e��d���{�ǳ��S�_�F2�a�ꬵ1=��MLJ�9�m�j���^���y~N)usut�H��\(o�ĎT��u@�cHa�����N���vwQ�d�{ӌ����W{��T%T3�s/[H>�0����ܑ�L�L�7�nMY�Dsiδ�+)�)�)1�Z�=p��<ӓϥ�.������?��c��b��w�Y���w�I�	����'�/J�1��<����o��/��xX�?�*�Ne
u�۔�Қh���ҙ�W�_��0V���Z��� �;U{�mx�^�b^�L%�*�����oX�l�MF"�a�a�ym�y ��'�`s���艿Y�m`���oWW��9����r��a�� �m�$'�҇�H�-�A�l�Z����H�V'%2�ph�n��m����':����c�+��v08}DV��B&�ܗ\���B��w\?E5�<�fY�j4���BcvQ�cI���q��qS�Ќ�3=l�p�ή}�}: _w��ʼ�!���Q���@������d�n}$kSU��������>E)U�F��G�#�ˣ2�Kji�����)t&��c�.�3`�MJe��4��������(��W��R���[���al�M��փs�#^�'D����U�P�)�s
��+>�x���@Z�Z�wu�y�m?8��0fG	�s�.R.:Fz*#�O[B���u �3Z��'�Mo�Wt�~���B�n)��4��T������iw�����"nl� |eP�a����M��G�����i�IlUR������UI.��I_kÁ����i@�ج��s����r���`��5��aΩ3i
��Z�F�^J~ui��A�T/0����2H�(Q��t�+������B����&v\`z㓃;qdB��c��Fշ��ej�o*x�>]�
-)��H�n#���U��$�O%�r�c@��鏗��c�W.�׷c�V��^�����Zd��f�}�v�^��#��So�������t�M�@�bV�0�ՊQ�*6��Yf?7���LLb)�h�f�N�?~���]x��O�ff��+�\K!�	^J�i�	/#����u���	f~Ū���A���Ӗ �[�X��,�pCK><�@��_�>`��s��a��>�8h�`#����Aϡ��@��9����ͩ�K0�=�$�\x�����Ṷ�(�D�z�&Q��Y���K?��S�+B���ȽPn�	�L��^�N`��Z*~y���ԥkR���Ī����bNt����S�j��䋴�a�(������ڿze����4}��kAe�n�A�PX
j�f^h�!T�Uɏ�뷋������p�����2 ���粆ja�@جq�̖DЫ̤�*1DW�ھ���;���_��<~l�-��+�U�h�.�����d�j&��0�ם�j-��N"e�&y!�B}�ă�H��1�x�.�7���`��qx���X�y��ble�ID�x3|�'��T��	*i�U�Z�K(O_�o>t�f�9P��.�M�::Yhw#\��>����/
����y�j;jY>���B��'��J��M����s���`�OZ&;��-Y�'���됝uӟD��L��eMkPzh˴'��q qL!�us�����EC����'�]�q��`){3<96�����4�����;�_�K�f�m:#�v��i�PLS�J��%���m���UL,	�h�Q��}qP��G��'�4�W,����;�[`k�R���V��@(N.���T���X���c�DWFR#q@}�����E:Mbθ}|�C�'n;�*�����_8&���e��4@g�d}K�/l6�R�aG=ɛϜSp�g`�4�ۓh��T��_w7uȎ��G��%� ��H����z�U\��-b������o�m�А]��=*�[k�1��������F'���.� ��5t�����e�]�\pu�z��P��x<�hy�) I���NZnD�[�@	�;�qRx��8i=/�ڔ!�3�m�����#	�Ey)��s�)�Z������� �Z�Q������=o:μ�y^W�ϬE꩹t̻��ٶ�O�[����;X�y~�>���կ>�\��Ј)>L!L!惯��_~Ơa�R��"�$Nc���b75;��J'�����(���7��XA�a��g@��M�x�Id+Ԗ��g@'f�-L=3_�]}�3�����L���u�1.��@Z,�+�yK�ҙ[Zƕˑ���~���1�Z0;�.� ���� �H��X�qB&C�9F��Y�4B����ì�{����S���q������$�<��@U������͆"�0��-�!�5/9� Z�21���$�U���HL��f� ���ޏ��G�=� `��@��rAo2+7��p�Tq�������^��@��qN�"��6��
�m��1�`�ʻ �9u�-.Yb��Җ�N$�D�Bj�@�n�����T��R���{��*��H������؛�_�Zm�`J<;]�R����m֞�C;[Ɇ�S�9���6������K�W��嶈�S#N��_�9k�\�;u���F6�xh>-�x�<�O��,� $�6�*5Fצ�ҵƚ
�5�{�����`�54�1^���p����'qQ���`��K��z��l�
o�R~��v[U���×�R��K�5k����n�	+D1"��S˝8UhV�O��1����@���v,g���=*戩$|�1�< 2��7���Ny�ˢP����cO��A��zb��	��T\�����h �A�W��@đ��k�`�� ��V�JN��ԙ- i"���ϵA�c��^��a�D���B:Ca�C��_9T���:�������B�Jm?C3�����K�80�5���%n�d��BY��e3�[���з�|��$�Xi����N�h�k �!��(h�'�va��Wn��h�j���y1����Wi�*��/�P�!K�@���2[H�Ӑ"��"�m]�>�+=�A^;�0NB��T��b�Tо��U���WIn7�M�b�.�;��d��-�$=S�u����m�nRO�$����濩P�x�(�мkR{��Ī_�c��24�B"�>""A��%IJ{�׈�i�#4�@ɊJ4�6 o6�` ~�@�-�,�8���lvF�m]��������n>�B,)�6V_�&��A�N�g�S����-<
�Um��c�`���C�ˬ�'�,B�Y�u<����![��cW=�,U��i�y(��I0�'~S����`����^���~�[���~N��ʄ�z����.W:�3+�K7��Wv�a�Φ�{vd��x���N�������-��}�55�'��������irV�����=>�Z���{��^�L�)�1��^�,��U���s
	��� �.�z�`�b�)�ʶ ���~9j-_E��������p��80}��!�Ed���t7�u�oO)צ�Mu&����%vt��`��F 5U�xZ��U��� F�
JD鋸�5��#�jN����]�`V����/��� x��8�iF7�!*�cDB�w��1�%lL��%8��ʧ���٥��r^ͻ�x�]�|B�0 ���9~�&x��!�ҖMu9�ݢ3��1��8U}�ڊ@z���w#���=P��)�9�޾�fL�	��47���NK�8��E�����tT+=�~�paD�9|�����64C�Iq? �8�%��@^-�rq�b�t'a���@<��y(�i�u7��Ҩ	w��P����Un�Ê���zZ���0����I�|{�J�U�ޯ�+OZ��ۿ�`*=H��s�TA�PѮ�JT����΀w��"�e��=�Z*��ݏ26�{x������� ���h?^��b#˛5�ؠoٞk��2�Q�<Wngu�zu�ޚ� S?\��=�-�J���>�ګ�	���م�ٖ����/pN��h�jd�y	�*�\���/-�̾z�+���lEF���`�U��(�j߽<a��F��"�|���%p]��ga@2�O`D���hz��?�@�!�b�4Z��.�T��;��&\jg� r��&���\�QWI��܎�4�Ps#�,�
����0���Px�=�%|�<�4�<}ﹻ����h|�1�ׯTa���#:�2r)`�a��S���G�)k�����^�aÿz6 /R�^�T��Z*�҂��~J����t� �2�r�i$��������z	4��3f���9t�Ku�s2����yhl �J�%�ڪ����O�?� ��u��'��ҝ��Q.4f��g7�;���b9�q�E)#�;�T.�nQ�M���T��>������@�|4t�SU��`���d����F���B����k���v/�����%\�h �)���"�	��0O#�)�G�*$�;o�Pӂ������9�!\ҀԘ��sݶ 8^?Z�9β�bX�����& ڪ3#X��;7Y��8���:̜��1}�9�1լ;��1	Wz��Dmvɲ��N���j��HD��ۭ���C������Kl#���Kj���0������F*V<F}��؍D̫���6�@����~�	�ɏ_�1ⴵO�,�c$�gDr
�[�R4FV������Ҋ�J�#�]Z�\���
�	�~ʹ�l��/c]�gů�٬ d���9s�ZJV̋�eJ�Ad[wa�Z��>�uC����zl�_'�LA��.l��p�uH,�����w���]��m��8k]658��Z�g3�o[���ڴ����	*9��2��zyx�������8�@���T ��pv��Z ux%�Zp��1�1=��d\�A;J�@�$��R%t@�깧��� �����q`ni�陦�s���d�����-U�3�.,�N %�1�J>f� qͣN\���0�Y��u���r�ƘAeR��*'��묬�H��c��	����@�����fRly����r3�b��Y����\��1"5MPkt�����}3�SC�gS��V�va#����*E��1�ԝ:x�8���%���c����A[!`�u�w�d�w˦Q;XᲬΤ�xlŃ��0%a���@-��E<�q�����U�^���w҆�ح����v�ƁOo���2&g6�j�3T&k!k��KH.�7]�u�Q�I�I;�Czł�-ύ�$_�g��T�te��8Db�E����~-���¡�-��5��V�! �g��������"fҙ!�:�� --�"�[�[���a5T].�`��ȫ}���M�U��U�q��N2�I�P5�W����������S+u8-o�~r9���V��+��D�����	�pP�<̘�!.��yi�S��!H�K�{��G唗Y,+�(k���`���s�7��Zn�ǲ?W��HJ�$]N�Z�!���AS@|$��?��$��Y��Z�c�&zb؆#���|��o�^vhJ��U���Bp�8��y�j�5��7��G�m�������~��HF:�fmV>�O/���A�6�rE���n�C��B�Գȶ��[)�K"�#��b���q�i<D ��-N\7�B���v���<i Ix1��\�.]�:՚4g�O���UN����M>���5|��vZ���	w�kP���c�x.����}�E[�j�1}=Pe�5\@Vd������WU�z/�)])�x�yW9cvx5��b��D&�����W��/4nL9�ĻG��و��UT��ܕD�H��gay6ֈ���!�E������ּ�8)Sq�r'��0g\�;�2�M��)�6�j!�`�����s��
��s^��i��������*whY�� M{y����#eP �f������t|�(-�X�������U���)|a��qDy������]o\y�G��Q�;�z�֎�f��-��ŵ�U����.!��8�m��e-��ln�s6�����;*��dcD��Ոm0G6I�O�h�0�F��tQ
�s�w|7�)2���)�U�E�Y�r�̉$�|l}W�80�nQ5qf�~�ࢃ��$�:'�H��j�a0)�	���E����Z	�/��$|'�N��Jǖ��$��L����S���m!LF��,����.5ag^��\����q%p�'(��G�ngr�� �ng�m�`"�ճ�c���6a=��c��+uh�qǔ�>Z�Ci�P���vz�@��cD��'���Dk�d�wx
�Ǐ$�h�S��t����4�'��a��N��T`�N��0�g�$�I2����pÄ����3�2Ͻm���VG�d%�z�?��+�E�� pLXADc�v��
�&j���8w����N�Tp�-aϹ����h	�.�"Z%^��G5S�x�3Db�ނ=�ja�B������4vk����P�}"�`bI�j�����v�D9_�?�2K�9 ��jc����@��<'�9����Vթ����U̱VYx��(��=�h!  �񫘖�t:�F�����������$�w�(d[�o�u���o{�n��$����i�����~�HOw?kE=�x>5��<\�i�߰\^RM�(:ǡ��F�m5����
�v��jbqmufu�`�\�x�T��:�I�$G#�q�Gɢ���v<�-}Q`��xOL���-���"�,�����,_$�0�ޞ]z#t�%(��<���a�m@7�<E�	�{Hvm��#l>:{�8��+Et#'>�5�(����Xȶ�M�Z���9dH�<ϥ�8!u��Ũ�is�p|NM���z�^Bv<[St�N���j�Bvq� ң���ml�W�+Rz֎s�*d��f�Ƈ�c簧o�D�Z#o����F�v7�3uB�8\}��0��I�����k'q��O@M�?N�e���Yʖ3�������uA�s�@Ѥ�����ãے��G{,-�s��L��1R͓F�����:h��9���u�&�EoU�����:�<������a�����8/���-�n�aq����ĢZg�t)��Ei���V���k�}�R!{y��$�L�(����3U;���b��VB��-#v�-�(�iUյ�t��a��VW{���T���cC����������0=K���ITcFp[Oܷ��U쟌wU��׋>�Nrae*$����[v(M@��UOǞ9v #\�"���v]ǁ�B���j��O�T�%l���Jv�U���֍��<���p�4����^�s�.�]hO6L�I��8�AZawh��![d��D7�ȶ�5��ˈ���@�<��A;������9���,ہʌPWJV3�f6��(�:�U�E�I�|�ݘ��Ѹ�i���(�<@�`��Q!/F��$v@M
m3�fL�S~���Ҷ��[φ+f�!<'�B�af�q��q2����~
��]ۈRC��ۧa���j��0[����$h�l��?|����Љ2���^-�8��,��g�h�����A�^T^W��:��3<��Ou)Y��+�[%#3�,��	/�p�9�))$��}	��������4��Q/�lc�!u�$��c֛�>�g���b'>L��n�&q�w9�
^��c�(�{��� ��3Ӵ>(�����J.3��u�;����D���%	!١|o�R';N~w
�?��.��L�N}E~��ޠ�1B����L�>ֵ�&��.�f�v����z\�h���0>��]wn�-Ҩ鞼���T��L�1}��a'��Î��g�la�qG��n���<隗GYXf(��LZ̝��h9�p��z�%݅6mt�2��_N�[y�N���u����t�&(�=�p�7��7kL1�+K�F��=�se>��B�l��'��^Bq�MLОX�`I��2�����Z@E�.��j�����k�J�s��`�+��~�S�������E�:	�fP?�l�^[���O� ֙\��g|I�^B�P�a�����xG8�Q�yw��Zy{C��<�*��8�v�ݳ�����kr�	�i�N13>�k�;�
�'��$ �z4|�=�p;9�ʔ��採��G�S�MIX~>TЫF�"I��Z�y~P�2E��ǹ��"Ry������g��AK1�	E4
�
��5~].ON�\
���&-d�9Ή�]+4���ʨA,ō'|�O9��C��╅<��N�?��mͤ�rz=�m����+{2��ܽRw>dZD�,l5�D-����j?7��g�ݘ���@��usg�D�;�]�c�rf��&�.����*�se�-�9	�����u1\�g�Rf��J��a���"6�mYbƼ&L���g����k�<Z`��c`���k��T���tn�{4{wC_@֞/?�0�b��kH�5U�$�qx�j�3�r�D�<��m5�n�ji�F�h�fJTSf:kSȎ��@���`���p�~TW&3�t����L����������]���!#�<��Is3�����PsW��O��w]�od��3���"���z����4PR�6��'N�"
I�Ø�����h�fe�f	������W[`P|\�PzDJ<bc��$C`�.���Y��(O��KgT�m�Qgy%E�yU�C��dWϕÄh`�6��b�b�z�&`���]&����+�|��L|
��MLmߍ��T�&�+�>�E#l��N�[*��{�S|�={�Snq���;��"Ԫ���[5^V�6Q�����K���-�G��˥�����޷b��^}X.8�T����ט�<o"�{�L�wY6�gq��"��,
%��@�w�0V$s����AH0Ժ)�5�	~�~$�AJ�����;�?;�
��o���y�tM�ٞn#�S[-���0n"�-�-�����>�&�S~�#A��)�[�t8�[| �z�-%��?aگ`i��)��e��v��VR�A0r�C6>+��כ�f��P����8���-�p�E8w�Հ���0���(�ъ�꺳!\�� ���y�7�?)?��@����#w�t�E/>����Cy�b�Ѷa9w�X�u�aIۉ%;���3���z��{옆�$j�^r|?���ܰ��7}q!�̈v��� �
��vIp����n]A�����IU���>���Ü8L�+�s���&b�������(��������vET*��F��Ș��4���9� `�#�/��^�PU�ח�A�a ��{k���^�6W^K��⽮�Nm�">�3��}�M����z�CL�%�v ����u�ZvL~��D�ɭlz�Gd=���p�w�g�� 3�㝟AwA�o�ޖ��;%��>���Hl#�9��ĺ�B<�VKM�������:ƊU�`�Y��A�����˫xp"���?��k�?F!Kv�֘��OC
i�3قѪ��#q,s�>��#�z������Onp�c���&Re:�&��1t3c:�-�ms_�0R���Ϭ��@��W�ԇ���ß|�����h͋��L
PTG�����Z�	2��I����uI��%��zl��2�
���'Rz{.|\�9!���3�~2���*�xm��qhi��帽�8�p=�B&ݵL�}oX�ǺZ�+�cf�uj�y�j/�r|�+�S��m�	 �J���%�{a�aeD,�#�"�i9��RM2��[����mf��#mٳ	��5�0J.X�@	�J��'�'�R�}�^��V�ؖ�Nх��0��a89Go��[K�Ag�x�
��M"�Kb�4���{��e��.St���-��)Ce�?�?w����]�d/k�r�{��Oǉ���qRG�p��q�����e嫤!�E�%��E^��S=��\���������"��?h�:崌z2_|z���N4�`����FD0/�g�!�/rǵ[V;�.�S�K����Du`�2�M>��|4@�Pɗ�� 	�D���e�1��f�Z�٤�BF ZT�x��r����?����'X���#j�ܵ�4z����0׳1A���4B#�y^��|�zz�� xՂ#��� ��iH��I#b���K$v��V��]��A�����H������&���:��ax�e@�[�vg:�(���R�~a7|1a=1�CU�� H���r�	ݍ;��0��"��]B����?�29]�������{��Pb�a9s��5��c��֟M׷G�E�"D 	˒��mV�T�?Y��ZQ�Q�.ջ���e�/8T�	���L�_�im��s�����BC=�$���Ŝ���It�F�Ư�vxU����RRV�8�6�XηϱF�B9�-�������Y׾%�$�Ku ���=�l�W�-B�\`��%Y}h������UIe�A�@�Ĕ7��H�y�\+A�p3�k�x���q9��к"����Sb]�\�P1W�UGfH}{ �0^Z�<��W5��A���j����/ıK�?�'sZL�-4�.5�[2�w���H �����t�c
�[�
mi�<�>�]�f���DN�0mZY�W�J�5�-�n8�� ����K_4�ɵ���z)���e4�O$�ڟ,gq��nȷ�1�K��t�T�mG�cZ,�|4�5��^I<��y�.2��zxI_���m ��l5N�^D�R9�C� ��k���f�
�2�+%���� mS�����"�)�@��7��/]�#�R�m�	�&]�>�?J��	���ry�Kk��79��.m���CY��B�M���?�% M��#xF]�LK��Ne������)4���$S��~(�]1�P�"�V^��ۧ+��4G1`5���8�b�'����ͮ��6��?�\f�&�1�J"�'odi���y�X_'�A���Ph�-�!�8�1��Y%n=ۓƘF8b�'TYH���(]��5�-O��m����̛�?�K�8�.�[��^��u���k�����z�5�۩�)���m�k^Fn����m+�#4��oc~��y2�T��S�rx�|a��XkzS��;����u���FJ���j�4��mBUL2�V�s�P�@*J>YF�~���ʼ��&k�b�A L�H�T�E9[#~��}�E����m���a�N���)�x@��pf �wj.x&���?"K���E�cM�C���[�����<�V1>������~�CӶ��ϱ��3hq_XE�:*d5�H���0x��f�6S�,^IvB�\4~$7Tɜ���a|S���(�ԅ'�w��0�[�\ý5V�M��4���0pQ�����8�@���U!��c������ǻ��cL�ݐ_�
��,�������ۃ�Ȇ��7��d��8�	g)L""�S���h�-Uw���8��ǿ�y_i6���Ʉ� S�:Un9�x����w������4��/��A,��x��=&q6�0K����Ƅj�bt��N����;�G���i�=Qv!�xGJe*�5��<D��� �X�ks�p���o��9c$k�[���pM�Jy�z�2c����	��2ێ��(�Ol�
�����7�4���RLt�>�܎d�w��w`<�H��f|dz�:�(]��Ի��6imr#Ѓ9i�ąP�H��dNY�E�k�����E�F��JQCt�P��UU�ɪ��D�quf�I��$H��<e���P\���R�cw���o�ՠ}l�c���	�Ƞ���5��/��u�?c%�ф�<��G���iL������M"��?�d�eel���"J�n��@jhZ7���=���F�{'`t$�%N\6�`�h�S��o�Aަ��h
�Y.�z�I�eM�@�'�r�9'���3�׸��C�vB����A�G^��l�f),�C�u�ݒ�P��_�"��T�������W�Y}a)�bYk4�a�-s��c"|n�k����T���E;�󝦆���Ȼ�x�D����=�o��
��R_K8h}]��MI͑����5��y�E���N���5{$6�`�s>�@-�^-�v��4oE�@@T�gbB��e-��;�?,�;_4���p�c|�VZ���x��[��sXh�l+vy\���D�%���U����0T�#mӚ��llr#I'~�l��N���ۅ����*[d��3�� �����=MTM���!:c5{��C<��LL�'p��C���	��o~&�j����2+]���g�����B�I�r�D���i�Bw�/���:1+��2B�-h�7!��s3�j�4D�Kk�Y�YF������S|	�E
�5�D��FO��@�D�Gg���K95F�Z��ӯ*6 TAc�P~��"%]"*��\"�ȏ~��m}�j�D��*�~���L�J!�{P��*����(Z��'=ş,�]�7�O##ǝ����+��1~N��J�����#%6�d�~�D&����s���kTm߫}wm��X�Ȫ74eX��N�l1�^�-���=�b�W�^'�+z'�F�=b�a��Wk�Il��i��D�����NGٲ������*��Q)�4�QO�F0���O�Wv��l!۠Ȁ5&YG�����i4>ц����x�
8���6m���(VI<�]G�D��^��wO�"$[�n2`B6�
�Km���,�5�ƭ;G�S��<�c¹5+,,��o�UA��Ww�:� ��T��̒��)�l�}ڹn���kO�)7�'W�'�����9*o�E����)�#�~��'�j�z� ��5<!Z� ��A�: ,=L���ckGe�Ѐ��[j2� <*h`z�X���q*���pk̊��W��@���Evԕ�_ ��_�{��U���Y�&
��Y��;�rF��D�(7'(�W1�������#�nꡠ_����lEi��CnQ��	 %����n�}��[��L����H���6�$s���$�+�wjuW'U�SS���b j��f�3���Q�h3��h�t��:쫢F��ꆅ�q+�vW4a��\ܰ�z����PD"�}�S"����
�����Ĕr��]#�O|�+e� �4��BIO�s�cB��%^���1/gN��/u�x) �bW���,S�|��So�,����(�Ĳ2��C��`i.��Ɏ���8�>l�s��8�>:-�7�%� HU�u�?OB�.m1��f��w�Ã{iC��7�?��,�����������#��ȖBVQ͑�����uף�6X�<���;���g�ۆ�q���f_Ѫw�"�F\�)��۾禾���'��Q��ܜRiL�nlȝT�M6�{�!����ֵ�����͝B�7�5C��Lj��q �\l+&�%��+$ZA�<uL�k���R%�r�g𻐉
	�yV�����=�L+a����d�t-���'�i:����j����ߤϴ�W�S����'.�tF0j��++��.�U���j��� ����B.���U,��y8��hB+����j: �vg��}���5g�vQ���X���dӗ��u�����6��K��{��p������º-�b�@���g)*�+0t��NB
c"��S�}�K�N2�o;�T�ݛ��籓�l����PWd�Q��ƪN�}rT��5�h��zۀQ�J~����J��|�Qו|���G�Z����~����P�]X`�'M��5�H/~WP
����]R�B���"�.G;���b��H��̼�MI��}�h%ݿ��v:i���/��$��h^�}����˲x���ǽ�s���B6���kU��_�?�����x�������q
���t|�rK״�XT=��,#�p^�(OC�H��D_j�θ�&�s����F�
	�=�|!0]u{�¦*+�$J�Դ��M��n��ˣD+e>��.J�s�gRLGT����rS�!/�T ��q�]��`�g:�\�P~�3�a0��<������Z!ǝ���v��i�������#��8���B� _��_e�v���W�Ց� E���Bts�K�9е�nW^9(>e��4�oo�����~G���e��;5�z�m���ȋ0����}Y?A�`J�� �m9�1i�RC�a����^�l��'1�^e4d>K)vwéɣ dNuwP?�;)�[jr���Ul�"�	n��9:(Ǻ�q��ō�ϛ{DࡩR�=�0<p�+�����PΖ�яH�B�D�&r/�t\]~�(�������tp���dX�{�PNo�y}~Ƅ��VB`�k�q�x{|�v^R��e*yL�NΉir�ȣ�l�n��Ǭ^�.�E�:R��K����U	���qT�,g��r\=��c�%f��X��;��!�H�a��E��� F
n�T��f ��
��V�ۯGm�����g��������&?� �yn}O��
��yS1X��OP��~��
��Q��� k`}-Oϙixɜ/Ŗ.Wf�;���^e߄��_ �?!�,7Ȃ�ķR�h7:�H&N�O꺊N|��?vƉAC�;"z�K�P��d�^2'i�I�*�� P/��1�	��/�jֶd����hM�*U����n��v�yH<k3t1+���|�����dA�i�nN�]�ٽ�g�74(]w�K�$��	.�3͊�� ;~8����0���6�>����su8�3-�܄
h�-`J���/�r6_a)��ۜEA8�,$�7_���ǂ�����d�Ԍ.'ɏ������[Crۣ�N*F���"�{�;t��P6���W�*9�����k�U����V`h�d�++��=--���M-F<ׁ�z:�)�3�*�w��ޘ]�gC{K�a|��!~h���ׄ�oG3J�����2��bwYQ����d�M�,>�S��xL0/�����L��T'G����m�w���ȇ|h3|j}��M0*��bϻ��r��nça�>�r����<�!����x���Q�j���v��xg�]Wٻ� �ta��~E׽�֛5�fѼ��ɞk�U|�u�B�=�-A���/F��p
%|9����O`�apE�A �,X	T�p8ۼ\�|K�0*����#�[�$sߏ8�<��g�=�!gbR�Yn�UL��Tl\�$������:l��x��_7t����q���wa����&�K����a�}xq6NUR��2S�&�s�)���:X'R���Mzh��좖6̳
k����!o�,�AD#���H;F�����R���8�;��A1��[Ja#�;�7�� {R9A�+Sb��H�\^W�uc6fN�k�/��e}K5��c�=��"d�����C�%S-F{��R�ݼV%1�R�-�l\�W�]^��f?)=w$���꣯<�6�&�KDT��*�M�����4:�d�{^��������Ѯ��ЄS���Ũ�'P��[�y� z_�@8��'z�Ks]H���In�����ϐ��0�jA�<x�Œ��k7_�D˵wj��)z&�G��:}`$��_3�ΞX�GM����:��74j�Ԉ�
��#�m�d�xx,�1H\���"9x���{�=Tj�5HM��� [���[���m'v�<��/�����Ath�>
���.'�O5�{�F�i�ƈ<n�-�1,^����4?��l���<=�>޽�h[���:����I/�E;�K7�<�OB�XI7��@K�H|��t5�9�$��j�Ԟ��L�{Y�!{��W@	��Tg�YQ2W�ƥ���^��A���D\h3��c����
!;	^~���-*S_ۻ��I0���=~������JgC�T�pH�w�{)�^iA���[�I�|'�dE��:lU�t�OH����v8��jN�qc�<i��$��*�R!��d�4��$'Y����4�CMJ؅����w���$z�6K�
�M%r�O���,X�|]%�v�k���E�7�۲q�F6U=p�cԉ��W��,(*�B&���Pp��wR�پE��s��?FL�	������T�y���D��h�l9.����Y���|�A֮�����}')�4��2&&@~w�:�B�f���N ��)��p�Y�%��G��d'�M�˾R��R"���*E����s�k%���JD�O��#SJ�}��N���7��s�wЛ:u?��߇ȜX��p�-8S��uY\�w"�4�Ox6*V���bQx���*�ݳ>�&j�PN_/֟%���2xL	���9z�k! �U�QZ�F[?@�ۿ��v�.(�)��om����=8)N�!+�7l��t|0�b�o\�i���a�tJ�3��ZG5Y	�]a0�{`8��v^��Ncu]:��|6��U�p��]�̉x�
�B*@Z�P=�`�Uh�C]6��l�஘>��@�H�\(5����di^Y������^�8�M�C�bQ�����
B�o"�������{���Ew�پ圷�����1׃G� (Wk�9D��- ��Ѡ� �m�����JD��L�6]��"�H#L�~��C;��ob�]S$��<�/U�����F�bC�pZ�ֱ��'P^�D�07é��d��W��B�z��.ƪ3�H�j�̹K�@#�(�r~��uǖ?gU���27��Z[�<�L���죉-� o0����i���\ M�e]�hI8K��_�X�g%���h���!�Ι*8O��0\�����x�ю�Ҡc�;s���U(�9��H8�y���`|6@M�Y�ԫ�UZL^@�y�qӊ��{?7w%9�Ĩ��i̈S�(���fܠ�,?�t��('ĠYL�'5D���1j�;��(����|�FK�P���ɭ#r��۽������w����-��G�b��W�olN�lǘNG�h����1��W!I�c`{Tz��0�[8�8�&�EZ����6N(��\�����%J����щ,7���,f�Γ�7���0?V>#6r߷Kڌ~I8�e����sJZdQ�9Z�kG�=�pH�_�w�����Oy�7�R����S���#�<Ժ�ca:2��n�:��F�/O='��P<6l0�K�Fa���g�A,���,��<��| mTo��:b�O�i,9�8`�.�v���2辈*�z|e�!�t��5��!ѭ|�hcn�ٖzy�v��'W��u��ۦE�AN��cұ,^9�z�z�dq�)���y�=j=��������|J���?PKSVPf,��O��ѸKpP���$�P\C���G��b�X!�Bhw�(7��Ş���B%<BjB����JxCCxr��?>Կ�UAZj4�l��թڦk���r$�}��ɫ�@�ۉ��
}��K �C���]�X�PK٨��Ȗ7\@�XD��J�C��{-G��O�v�D�-מ�-P}S��
\��4��+�{�M��q	����Ɓ�
o�n]�K&���G@~ٝO�dRy���yZ�	�?���cS�g�S�J�s�y��<���0�#�*��n}R�?�>I�/���!:'��K�b��Gk��د����ߠ{y�\����q�a��EӋ�\Wx����$�� ����]�؛���.�YD�^�%�t���վ��l^�=@��jW�.-�5FQ�$��J,ϵ�B,�>�� �����
���	q����'VN��w�Ӑ��N#��`���-�Xc�	��@��e���d�����E�m�ܓP�VT:�6m��h~�e��I����"�h�ñ���|gF%K������O��u���D	w��;�$����DŲ ��sn�m�5&�L��l��B�ϝ����}��HU��>c�}	���
���x=%�͙ߣ�VG��ťc��J*�3��i����匧3 ���N�5{ի�����⽮�60s�5-ny'�UD'�@Nb��Y⺖���G7�r���j�^��=�����p��@<����^Ž��3�s�]%Zd��\��P�u��: >����5;%�v��̳%>[W-qIs��wK���޹�y5��[��ͼ8��p{:Y�m
,A,C�ܡ�?Y1�
�I �n!;�T$Dz�^jȱ��͟P�Ő*�DC���M�{^�<���qP���n7��A��*�;u�/L�Bw��iA`z�Sǃ�N�E��%���R|��f�H���A���H�2z�}��|a��Ƨ���k�c�
|*؅����w�b߂1�vA:�b�p��wX��TR��@3�	>/H!�	D��%�=�/��%m ��͹u:O�-��_���t��Iݳ�Gt�
�xXW;ݲ���!;�U?Ge���� �;֌=r�,�3����;���l�4Q�L�����ta�־J�\3��qJL&�9�LE,��j����хo/�p��JkmI�w��Xz�=�^j	(�����;i`C������7��%Sv�!ԭ.DH[%ہ�V<�4>�ǎ�?w�σmbZj-��6p�H��`?s\q��_u�BS�.�u]=þ��=A l�M���r ''�=���w�.�5Q��4�L�|�+�Q�l�$M�'16J�U��R�(�3�~��t2/����,B���ck����`]���n!T�z,�VS�ޟ����:�����5l�� �.߾�ؓ-���XF������������<�-kP�ʲᇰ��t�JZ>s�3ת4԰!�YL� ��u�7���io֖>�����8�F��~\#dk:� �O�d�m�Y�W "��d��2y���Zf��C�|��f��m"�M����M4t�p���h�%
l^RF~�m�I�~���L����n�ڦ&���Q��s4~-	�[���-ĞݣHCk���@IT��z���O�����yo�6��.��§n�d�1|�辁�!��"Z������=�S~9�!=`3=��j3E�фD=���V�Ε��:+�G�h'�NKW��O�����`�a�6Sg9���~���ƣ|����m>N���g��S]�2V�x=DYZ	�$��T:NU�	��F_Iz��y9�Kp��t�V�'���+3N����A�:���e��dV���e���E�ȇjK8�����6��s������9�)|R)�vWu�<��f/�,�,5�!���-�ʰO�������t�[4?�'��o���[PD��kb5P��_.5SP#gn?,e�c��B�BiR0r6w�=�i�!d0tT�ȫ��d��gz&���H�5���s�(���8���̔l5��zh�������<h��A��#�FhО*�@��*9��� ����|�8J��..��J��S��l�68K�B`[#.�}�&�������.������- 1��{��͞o.Qx�m���N��<��n���I�(�n�]!f�y['vi��_�'\wgr�.;q��=U�6V�%L�g�L������g k��%.���PBb�n��k���Q�ta�ݹs�w>ϕ��@�0��o�8���ۊ2l�x5����^�>G�,x��'���(��%���n�)���ʾ���B�!�9pA�T�&���G�UE~�J�-#��M�@Se���8�s;�Kt�y��ە(���^ڦC9_ K?�O:@�~S��W�0�)*���1ޯ��ɉ�Y�}�H�u<�������K��~�J�XI(�]����/v˦,[a���'��H���Kjʬ�����O��h��5;����a���8�����	tF#����;��cha�:�L Ă4e�wZy�
�@G@�.�|�A3�Vj2w"�e�9og ��H�-�{4�������2������N�~����,5�F�;��XP5n�:(i����sX�Q�r.u�{��@�q�ܛ�(�Ρ�����<a����")�9e!�2�U��3��l?+ �o�.���zB^�$`%T7���j����ro"�K)&�:�9 �9�]a�cֆ����#'��ӊ�@�y0�q���[k׌9	����Q?bs)g}$��O6?�}��mޏ��c�a����Ԟ�h��4ݪ�C��S��b]L����5�3�u��y���7`�{M
��/��p�	2:�/�Cqa���ĥ�gʜt?����5���t	mOr��A���� �C�{��2o���`sr�ҕ�+���C�B) u�|�Zq����6����=������<<��=�si��`�c=!�t"�-�$1d�XF.b�l��C7l�-�x6 'N�J�`�w����ޤm�� ������r�%<˓�-�U��\�q�[|����VX?PǳM3kJ��."�f��8F��EU�v��B����ƞ�Z�?�$�׋M�X��,8,�m��y��>޳QN��0�&�:�� �Bx��FZ��}��Q9ݱ�x�x=�$�Mbdn|�u
����C�m"�=�	u+`����,vs`�}�Qm�$c�6��K�1�5Ϝ,����B�cM<Uտ�6O���G�bGE:1�$:���%�7֤s�M,�>u�j��@6�,>���VK KW%�v��^�O�)�
 �n�,�#-��k~u��Z®_��OR�������S�~3��UR�ஸ�⚉��mKQ2�jK��G�I�vj"�������P�&G�<50e&��� @��D��CO��:�IH����n�e� �64e;�P)� ��H)bx���aƐ�^4Ԥ��Ǟy?��GH�U{�b��������A@��ƅ�����U^�.ޚ���;�w��������.6�|xܻ�'�v�q
]�C��x,��gݩ�--�D��9�Ңg�P��N6�K�jb��U�U!�J���=�@2�� �*q��G
�y����w|����F�r�Ȼ�أ���4�D=k�[ϐ��J�&��<h�@3-Exވ1O��;5��"����t���c���J�8��ƛ�:x�a�,qRŇ�y�%��Cc(vbk�c�P��S�Gel�'�幡bxU�$a�S�4��:X
�4�@I��4ܤ55�6�E>FY�~�`�u�:�-�G��{����|g���P&�C���ۻ]H=��|d+�$�ȫ����$:&	����=�b�x��;��.C�$RZI.����;@�|��$,�+@Ch���*�GY�?:�+��x��x��X�RS��]�K+E��c��_��q?[P��鶒���!�3���DX�YvwSk�P���AQ,M�0���֝�9�+���{�����f�} `۷\��R�x�@���4�V줨^W֢�uu�����Z�r��Nq�Ϣ<H'E�uu*�MH"~ۗ�:p�\�&P^���)���WO��p�~nAݲ3Jo
���;x_����G���)�b����>�(ϴ<�+]�J����e��_��CrU|E"+Q�$ �&��G�<ge1u���Q�dW�6�'�j���N�"u H�xV�pr�f����l���98x���ׄ󊈮�i/+λ�,��[.���[�I|�][�P]1�C� kS�К��!��:?�ٟsp��so0`�+1�by�ܩ��*�͝�ǜi� gh��B�F\&K�r.�DAW}k?'������yџ�����ҼQ�̔n�jRǃ00%*���1U�3Z�p�8#�7�K���HXU��O�2>�
�#�1߉	K�x
�4Q�+;P ���@-h�ÐS6p춷�"P�Z��u�ٜWƟ;�em�/X���3;��	L�ٟ.�A�7T���GV���zy?V��Oz��������F\�FѫD:q�ж4�Y�J���6G����3ٽj0���$o�3�`����E��!���(����b�c�I�+w��K������;{�x �5��vӝ�������S�
���·�������{�zG� j��׶M፵b�6�b��ac%�Ĝi{��A���m�u����Ѡ�}<,��Ǟ"�I�L��sQ��}�Έ-t'T��_:���m^�VfIK��9;��A���I�����j�	��Q^D�;��������㝚�����	�Nsm�S�C�l�ީ�!
Ii_���?�0�:$aɖ�Hk���3z��{�*�j��9�u�r���q�摛?��V�Ӫ�>�m�����,�\& %�Y�+�11�X^���i��X��PӴ�ST"0�j���^�����Y1��AH��t���������mw(��1�ad��8��k~W~=��G8s.��� Y��=G�y5�w��ߦ?�&��mK��$ A5��Յ�moj�z:);��tT�=p��UaW6*K�dz+��� �f[r �Y��L�P=v�b�ă�Yup�bz���ެ�b��w�)�AOS�3�w�f7Qvf�[
�}��glD��bG�:��G{0�>,z�����ȍ�����ڌ��v�jjO򹵚Ux�G~����F�e�9�!���a�O+�ʘ�>���R{\J�N�'�O	���� 3]���7���ѵ�-;7�sq�6:�/�_H�lQQv���qTKn�QM�4�D����2+R�'�z��C~?C�\�7W��s�8Ɖ�T/(�%�a0�!�"w�>*WotGl?q����̨x@7h<s��>e�Q~�������Q����d�g�v
�ו[2���"�+
v�*-jH�S���̫wĉ��f��;�mm�P-ې�3�g>"L"ZR��A&ڃ�+��fk{vZ�,dP�J5�#-p�X�����]��b�^�ؑd,J�U��:2I�;L�k^(�+Ap�=�Mj���'�_�E�,٩�3¥!��S����0��y�pmw�x�7�m��9R����KS�V�`�d�Ag�Ċ� �x��&>x�UBX���bQ]����kם����c��V�=�~�Y�����|6\�c\d?�J�$�f�i��@�lM�8��`%'�V�yŚq�:E*�v�4ګ��!f���L0�p��%��䎩9�dA�0�z�"���j�,�ϧ�^0�O����&�q������e9�
v�����Ǫ;.(����vӪ���? �CeQ�8M�L�&�A��9���������'���ψ���If~��ձWO�G�3�;�6,�Q�r���	�n��lѝj�1���=�dBk���0xo��8E��&j�%>�ZC�*� ڡ.�q�]��7���"T%9����9)a씞��{7�Z$��X� h�X��T���X��阋B~��p'����X�<Y�<��%;�����ߗ*aB�A���d�0����S��Cf�ܶҀj\�N��ɿ.�߬��(y�]�s-�N,E=rL�FMF��R�^;d�\P�
��z-�cԹw/�J���@UƬ>g6g�J������<��`9��9)t-V��Bc���T�!��o8	k�Ds�E�ަP�L�4�։a���[
�z`Y�{|�0Aux7���{�[���x�{�x��@��X�_��P&H�1���jP#�ԓ�����A|�C�.�,G�8O���(�[{`W	ʣ�Ϋʷ6M8!�
@��0⽕�g�^��:�L�Q�҇����хy�[v��a�Ռ�f��4~��v��/��u�����oC��<�7�\ұ�P���Kaf�.�dǿ+�N�����O'U���4l1���-`␝X���jZq+�3Y��6}2t�rT���eH|�c���!����2��
�'+n��lc���]wI����xF�O�s�Y����
dm�nV�E��k�syϑ�W�6o<m����u9׺O�DZo��?FL\��ߓ �Fi̿�*���S�a��vo�>�/�(�kw�X�m_.Q�Rٚ�/)?�v�~-����r9*�����T� e�YM	��e��a�j�<��y��S�1��00`�
6�u�%�D�̽����Y$q������V,TO������O�l�^�O�3���I2�%��h-���X�D��N�Ѱ��G�H����Ճ��(j�����Ֆ����Bo}8���޽���[��?
��,oU�۝�UA��"��q��D�D� 	;韪�Xq͏���,�D�Z�bn��g2֩y�Q��G��{����=y op4�X��,���V��aJ��T�����y�I�Ml��B{�+2�Pe
���棭��:���D놠Q�Zj�#|�����tDm���/�8�z�E,U��U�$��O�=Bt8�ޗ���x���t���'�(}q�ӘFaa��)SQ�;K�3ٳ��e���4^G��_Vm��w��
dD1��|�ԕ$}ڨ��4XUkXY���PKr ��525�ǎ��GH�_�@���j���_J2X�'y[:�E���*�ӯn��Vdܐ��%3���g���J��2�,nJ��B�S��/�cO�P?Lw��u�"#�Yp��2�~3�!��:��� �NV��k��]U����� ���v��),Mx3�t����EA���+�knЕ�fw1� ����rwӃZ�Ulž+�f���1�Ļ5� �z#�G�z9���jY4�9>��WW��TJ���r����X!��p +s�������U���kc���!^5��͢�c���C�MZH/ǍJ������>5n����8	T�>}2tȮ�TaY5��v�%~of6������?�SO�ۆ�8u�,t�7����x�R�}g���dZUf8����&(Nm�����I.t�<>(��yׯ<�ڭ�vQ<�3sk��-�p`���jW�&9�-��6�L+�|��>=:��S'o���!��r��b8�r庾)�vb���O�e��~s:�Q�4K❵���{��\�lj��f;�F�\J�~L�jMT�L��7�ܚ��ib?�5�fT�s
]d����?��DN�}K�Hʬ�*�
�0a�xlt8*����� ؝��mD7QEՠ	�U�eb�uʺ�c���v#lt�5b�6��ov��)!�4��������i��A-�m�aP�Ʉ��8~�g��������m�<3}*R���7���8= ���PU�>����~W:�1�Ij@�߽Y���D�[_�Eg�rٱ��nkY� N�	n��r=�]�Ī�V�j4��,)�#�_�ʌ�KI���t)�??��,��Wq��9fjv�e0���Ȅ�����L��S�ș���ߦ�F�N�A-5
_�R �N--ث����}�[�g��o���HL�fP��k�1�-�h���6б�k��������l��vK��湟�2�-,�p��&���w�'|d��M��uz>{�9����=���H��w*� �Y�l3t��I_2�D�0PZ�hj�d_��c�L��v*�|�zZ �v��O�EBu�b��Y�ɇ�����1��n���cd��r��5hvs!o�h��_I���4'u��\�� ���F8���hj~ �fM�I�kL��R��՝6�G��7j]�,v叀�����a����99t�1����l?�n�OE������P���'������n�a�;:Y��Z��V1h\j��B���>����b�s��=B���*��-=�ޫ�d�%?)�my]����ffo��'��<��|��v*�PZ�/"���aʟ~�҇����1j���!�N�즹�/���F*�65Y�����`ʕ�l��D���%�{���S慊���z̒�{Oc��R�Od�� '������4�$�N���upH���D�IJ��q9���)yW41|�X{k� b2Ė�Y�+N���]��((�pi�9ڇ���L��Ԡ�yz��JRIŔ��|�"��G���.*�����/j1�Q)�DF�68�	�͹��=FJ��9�A����(G'�#�It@g�	>w#�9��E:��% ���)$bg�&�nfD�:����6����D��FC����d��8$������Y:��E�V�~F&���O^7 \��&֩ݖq��܄e��>����R�*�h�N��k�pT+��Z���!Y-]������spy�Ҩ=,�,�
yl��������KЍ�½�Z��>;� ��`�:d5�k��?�ZѾ�:�׏��bb6+}���CN%4{qF�r�[���i���<n���Dxl�*i}6EM+�# #h\�ÇX�[C��,۾9���*���`e���pBŜlAL�,J.��R��p}d����n�RVC���Kuf�c7w��B=�v""M��6�͆�M�(�>�jh�����3탂:�H��h�"^�C��AR�tL74g(*2g>���N�m@=� 9���|������*���:5�EL2��=�R�o\�K��|K�SA�Wz�+IK�"t����D֬^��k4K֜��X�ܓ�u��p�2�k�u�v�7��SK8`�9�"�j�fE���������_@���_�f)�Q�b�+����S���L��8,H�n��.�R9\�U!7���Ŧ�G��WW4�ٰk��GFV��[��c�����<��K��s����;�K̘�}�"� 2��gz�(��m�3�Y!�ȬVQM����/��_����u�E͜�z��)��)�2g�Ty$��7�FC���mBU*�<�HU���ʺd*!$z�c𻋈��A��\ya}�M�+|+��mHb�t�$�Te�Lg����:R�z~M��}����4������⑍�2˗̖�:*�I��?5b����ɂ����n������R�k�@v}d�(��'�����˟-J�v`Y2����:�����D1��B���hA��_-#Ǭ�M	 X�t#%��Q�#��Ք�K�Gjx���`/i[�"�@��	}Q��Q�r�"`�z�f�50��~,�z֠(���_`�o�>+g ��$X<��F�c\����
�£!�$�!i3¯w.�����;Y��PҢ�X��
1!G*(#P��ڲ��|�C���w><o�Ir�5������S6Vi�r�-��h���9Q�Ԕ�η!�|��:�h������E\2W�d�5��jhMTe��P9���N��>_(�(}��C�f����L�����j[C��㟏�|��O,�퍦�M��(���צ����F"�V���_���3od����`8�z�y(��S��I� ��k�^eY�m�js��1�-	�Ȫ�I�vY����$�c���¯�_T/z�y2�����#��-�Ju ����w��N�O"���-���}SP���a`�9|}�C%�P�{��6�i�3��a�;�|����Z,�LU��5툋�w��Y��K�vm��n��;5�r:��CtB��\�&6����
\/�dfAV|aca��2��g��aDc" ܂���R�!���x�~�[��2��/�5�fyr�ȥ� ���eF��=��LkT}�aL ��Jݚ�V���^�C��T�BI�����s��i���/��ށ�T���.�Tij?L��F=��!�v)`�17:����g1��&�O��_��n����DGt�K9���Gxͻ�lx�ʉ�w)fx*_�g�8����^Ҩ!/��c�+y��ʿew��e�����iX"� zG�Փp%�R͇���5zKj!%T⺪�t�/NL�m>|���Ĝ�[�E���1�Y�.A�p����N:���'�����ibWtGM��Y��R���j	��
��I����$������=Bª8����e�y��z��D��l�w�/*��-Ӧ��%�=��Aۏ��i���(�����4F��g�-�Jf�㊂�9gt���I���N�\�U��u�.+�b��;�������I`-��r�\L�'����GFnMww��r !��4����q�ϲ?3�6�x�7B���BG�Z��9V�Em��ճQ��n\� Ȏ���R�
� ���q�u��'���V��2ϮsZ�F���p��:vG17[�ݕs�--��S�� Pd�&�w<V��m��`�5i3Aۈa;b7����G��H5���X5X3c�NK��&� ���W�'��8��f!`�t�N�/�����Lz���&�u�:?6�����D!h����ڬU`�/�Fq��ʺT����R�)��M��%G`��w��Ϗ��2>��ʳ���9�%F�M �;[��ۂ���w(9�eJ���!���^��)(F���T�H�J��1�3�k<�d=�P`��(�'֯����6X�r�����{��Qo)�Zy�!�/���!�W��5�9RM�x=���~��9��G	�);d!s�`�fD����*��N��8U����e,�^X^_>!�V*1�݇�e���;e�~'��f������2��ؚ��D���(\9�������C��+E6fW��i>I�2��nx@Ҫ�V���#��j˓�����"��R+��H�>�6���'��?���E�߯�c�W��P̱�beyf�'4��h�%��gGf�ڇ����_/,nG#�����r2
���pspy*����;ZݺR����������s�EČ��G���m@]�yHr��Ȟ��K�I��#�).62?�s����(+g��H�&�mU��A�a�3o�i%�W����FX˭���]%/�bm: ���J*����g��:H���F�Foy#��e�y%���{�f��=Y�瓜gA�@`��^�L�"C<-�R���|��أ_Y笮ES��Q�����~��Vy�k)� �y%E�D� qZ��z3GC�4
R����]�����5S�ϒl؂����fя��!r��|�������b���gm�	)!P�9���c	U\�Z6��6� p}qw��3�r"KI�C��Ұ�-j�h �{����\G �,@�JP>Fm�����N�P�.ԖX�B��~d�fC�'�/�~^������]���0��������W��yd��&���N�Z�Νq��5���_/���I���?;VHs ��S���+#�x��Q��\����k
n�w���t��o^iO3Aa����A�b��\�����ҫy����Je7Lna$+�F�g6�ل�T(߻CZ��0��X�~��رْgX֌q~㙃t_;��ʡ���HD�7��� ����vJ����_s5�x�PЅb[]��� �(�HX�4����ek]�V��+�z\༵�EP�j��|�>U�Fc����N�����s0.=p��m�ʸ~�x����t/b�C����~��9��8����lEјq�3F�=|�rs�8Cem���|&�&�"��_~���&n� LD�oGR�(`�a���8�ė�KY[*�GN�[��	�?wdzVy�a��m��F����ߟ�A9�'{������ߺQ:�.0j����G(�#��Y�HeT�J�z�U�q�-��D��x77M!�x-�;�kY^��v]g�NPM�����ʊ�N���������"����DÌ�� ]��@�?�����s����s�eb�a��"��G����o�f)
��j��P3�Hv��bȑV��q��*n�ſ���Y��.�z2��gK����X���sr�1��ųg)�)�px�u��:׌UWY㝧�XƵ����Q��Srp�K�(=�1�i�q�ao��i��[ę���|� wICd/ٜ�����J�YD�\��$��L�k��N�K4��GI�<jڧr)���삺��b%�����[W�
�V�����%q��|f�nt_|�Q�[��r�v�y�6F�����4ڣ�{jd��:����%`���V�/A�'I&Ӳ���Dف��1%��8A:R8�ǲ�FiҤ��;�b�F�
 ��#����җD��8n3�&�`^����bp%�~2�w�(>��/m�4u[�?�z�*�f�`0B�'��A�� HP?�X���m!Kն��!I�]�h#�ח�����N&�p���j�Fd����GbTJ��e�"�M�}�a�0Y��fmyv������,B��9�z��эzo�"�sc�YS�1�={32x]�DnY&���$����|ˌ)yIuT�_���_i�r�?l^�~���|��҄�S+��2�p7p���nnfJt����l���߳w�Jft���x�v��_�ԫΜ��xa��%��Ss�f��?��v���Csc�ODu�J{��eN-?��=��k��������Ϸ*%|ί�֫Ӏw�P������:�<�d/`�W\�i7m?��O��A��`�cX���i�6���~+���=�n�:�2�|��*�V8R�MK��v�R��pf��w�n��2Q:�.Y�6��%s��l���o.B���t�-,�"j8Ѯ�*ܷ2�y�z�	vzqS I�*woÀ�P)�Rǐ+a�Kc���hF��Tj�i�"S\��-�6')�8\�j�]�,���B�n���m�>*�ȵ �5�=�m]f��>#����t�FN����(�s��z'�V�	7	�pC��^^��/i_� ��N��5��
_��#( �R� Gcm~�o@n0���%Y���!���~�u�H@5��O��}P.�����`���j�TQ�ZG�Z'<�7����ڮth0q�@ gcW�{�W���jX[Y7���u	$��Ę�3"V!9�n����5�h�Kd8�G�F�/���60�S{8F�G���'�&Ó\�����"���\�4����-��_$ȧW��b�榞�`�͒ߏ��LP����S�S������+C��Et�nZm�,�'�zK��G���&;�RέEu�α�����A�
7�U-(��A/?]S����rŦ�Mb7=mV�U	�<�v8�qnvV�L��qE��-V�A�k��ۤ_W���;�dN(b��P5��jK&��8뛿&t�4�7K�'��:��c*���yo{!��.������.��!� ��l�?���	D'ڧ���9���V��@��zZP>�A!:n}�sOa�)D*��D\k�+F�Vc�?6E0�V�r��Bpn�nP�����%C!�bDV)N��]�z�Ng�e�(������N���=��mlTO���P���'�Y�q���1@�\�ϳY/��aΐ{�j�J4Ic��@nbr�5s��zSv�uM���A��Z�I�ɻ,��at#����5��W:�d����ȧ��D�M�/?p���{FYG)�
:�������1b�f�Y-�E�	S]��kY�a��[�P�=Z�P]��y[r���I3�5��B�Ϡ&W�K��孀VoD�}�aka��|Ҋ�25���>�s��"�i82�g��a�9n�AM}��9�d�H�-�'&�`�� �F��io�v��f<����y��6(�A
��H0�/��S_�P�Aӟuj�י� m�i�}\e�������.��uW�Se��++厹0�J��*����H�y]ɨ�Al�<��|�]W{���G� Oђ	z��(���7��f�?�h���������i8�v"�l��g���;�����]�YE�ߛwV��Jz�M�nNQg�ӓ_����J�q��v��v�A�t�0��K����"�T#aZ�+��;_΀&=#�y�6�&z�-r�t
X�C�)�Ce.��t36��h�:}�ڹ��������L��w���
c�DCڶ,:w��,ƹ��'��+�іm4��$_1 �îy�*	�=���e�*X��"v�A\����U[cp����p`��=U@9��6���m��4��(�{�A����D�^4)���U^W�����?W^��J�����G>��.����)�VJ��ik�=�U�R���&@ͯ?��g����:�= ��֥ܽ~�)�	��n�Ck�����Y���9�P��;qTs[h��Er�M�%B�S=.�Z�\�g�ҽ�Wbm��q�y@�C0��4�0�����d@�GOh�8��9r��q����_5�����VX�3l|
"�*�=8�S�K	X�U��TS_�f>?w�'b��vvkY���A�O���{+Gy����Y�jN5|�b�7�w"���9����k�h��T����^�[�|"!��)g�`0���@��]L�� j��/Í{
�$ƀcKVv�1�=.�bi| kc�@of� � �-.}�:ǻ������0$��;s����O��(̊K"[���G��  �*��0�rYx⹚� �d�:�\�4����?w�f>J�v��~���v<�P�_��r��m�y�*���.[Ul�'��lS�A�7 (�(�� @ί�n��Eq�Ƽ8�z���h��R|u�8H:�A��R��5:��w���1T�+��*S��r9�:�y��!d��ۃ�"%��� GS���+�[u9i��&�,S�͜%�����3��c���{���S�'h�g+-����uc�m���{7���I(/0?ZM�vڜ���~�}�|�&_� �5rF^��S?�J}]1�������F�U�����9��2}�Q\�+ܚrp���k\�N��P_�(��.���FPy츸��T1���ȣl$܍`��}�R(6�$�l[I�ø�4��^P:�Ȑ4y�H!�%L��3V�7W�ܲ�	9��S��g��@b�A�r<l�%:myad�s�M<Z f.���)����E��������`�] �+��d�!��K����
<�#Ji�<�םQ��s,)zl]��Qfԩ>�3%�!�������d�<.0��B�ʳ��/���ԮL��8j�A��8���5�:�	8K6�0:~�_�Ǫ�y<e����d���N���3���#~�LqV(>����0?�Q�wI
94����NU�QQ��ZeƩ:�a�y���k���-4xs���ض�w��4c��d|>�(l�m��V_l�n����)7�;�����l�/��遃���w����r���̈|��Z��N1lo�Hᗐ�.Q�C��1<�c[�.]J��?�qu��9������6DeKխ�hbFg���w���fsN�/�<�`��� Dʔ��]$r�`b��O��ԅ�و-H������������'$���˟����Xd7q�ʙ��M�s�h��z"�M@d����(�dP`�k�,i@�|��"ab�|:�,)���W��s��K�#%
��6��,6hR'�kմ��A^�>n~���3q�H�B� |	���JQ��,n0,� �*��d�AK�˔������fq���A��T\�)��J�֨6WN�P��T�b�c}е� dW�U�f���ǩ�<��C_�����`Tٟ-�d�;[oTR���� �=�d`B�A�>����W����8�6���S�S��R3֍5_�3Uk6U��UeBHCb(���.k��f���s��~��35�$�L|�9�1�����h�Ag-E-m��}f���<��� ��#;'<�@4Yp�7.;ǣ���m��9p���*{�׬ǆ�j@t�������Y$Gw_������8�n��7�ԝ��G;��B��|�?�J~�� ��ك��3��BZ�$Q,���`���Hw�UaO�6ڎ@���1��
�����k���#V���zB}{<PY�is��� w(�fEP	i"����2�gn*�^
���f4���ߙ�h�R��親�� �ahL�y�W�
�N��ճ��c�x=tZ^�v���l��C|v�}@nm�E��{�ȳ������;f{GC1~a k1<�Q�4$���i����}��0J�X��DU�~'�m&O/r����l���q��}Q������Km�"���{��5���!�u��ech�GԞ���lf8�;Ok<�u�X[�F�;r.���S��N��P�GŚ��7F#�����g�z�^VP�� �F��^U���a)�9hA}��Џ}+1Y5�0�̭jy������*��*B��V�m����:�a>D~m��o����=�IQ)3U�[�ϓ����}����c�KJޏ\�S�>T6z�8Xb��b�f&ev��>OC����tyy��=��u�3w���M1�g�5����.����'�V��Թ�w�{7�a������Q���7��1Êbj��"Ly�Y��/����?=�7���a6i1��f��h��K�zPZY����b�F��G��_�K�y&���iA<gX�EU�܁���1O�/�jI� F�TCKJ˻��>��Mj~!ݚXy�?�-���PN����b<���yB)���)]/�+��Ef��Y2��2')��p]�;x��#�>�b�}pH�`c)K�ڀkh�uB��m���ۗ��AK:���n��zUS��F��fW�C˜Ь.|gJ:s��A�2ޫ���%-���1�ơ�fg�&����qJ�W��j̈́t�瀋�:#����F��\�������\$,O�U���b�����~AF�}���na�H�mi8y*q� r�wH�Z�4�S�~�5/�T�_�<�v���Z�^�\î���B��uN;zlYv��[2 �;3pA�aHi�&q��#zzb��q%FZd=�l��#�f��/<k9�S�,T:��!��|\PZbc�9C(���	��'jx�!e�����,?�ue��þ;�1�CG��@h҄��p�`�������!̜���40�ތ�r2������9j��uz݇��- :���p� 늱��JN$� 5���R��m�Jٚ�Ȩ\��-�d�؄'��G���Q��aMG��&d����?P�����'�2��K:Q��@�<Y���s|�GsE)�\&�:V	��YI�������2i�wu|���� 8��/U�A�����
��JS- 7��a�Y�2�Vӆ���s���|F��{g%J[�`9��[�����Ub0����s4G�v;*���TM!*��,������!łݐ�_��]�fBe� |e�Yc��s��Z3/�'����M�M[Ko��#Us�;-�O�~�I���AC=A���23�c���=zNK�΍�Xq�!�f
SX�HF��A�r�Y���Ե�%3P�.�3}�]'S�js`��иĐo�\�K%�����<��L�I�giw��5�L��"�g�<��5�x7ߔP��:���is2�<��H���� �+K"Vql'l���*�.Q�3Y%���5s�����i�r�\\d�̌b��|&�W��[���G�2��&6���B�B���o���Uc��e=d���|>P���GAK��������>�d��ٓ���^D�j�o㣙?]�;�2m���Zm[m��oD���qX	a	(%	�7X���,̣�ߍz"�&��1�s��A�t�g�m���^��s�"#\a5|ͪ���B�[�չ��bo�����gl��60|���5������y�γ����op֛���U7�݀�����eH/8NH�&=��y�H�~:��d??4ZsF6� �3�,���n��o��E�j!��D�.�]�	��MßOP`={�!l(�HL2�I��$�A7�:���[Ir=��<�e.`1�8��s�{�UĻQ��|�B���b �
��� �=$a)5_c�����8��`ː P�UJ!�4��N�i�jM���Ň�e���16�3L���;�[jx	̛���ڝ�{J��4e�RDm�Օ\�h��B]m@V���--tRr5����Z�xz�(:��OY�]�n� ^N�ɲ���:��4���.������R�_��q����e�Pk���ÕK�{�?�O#�W�:1��HpF����^��eڛs�@�^�(f��W�B�����g˝��HT;G��S{����Ŧ$lz��7h���>�u\�FXm��UB�����$-g�	��h��j |�!\�$cfY&Hn��� �=�+4���>I�Q>�Aq"F��c�)Xh�(�M�<Q������׆~K�h�T�G�X*w��5���ԳV-��O����3�����x���T��<E�OLׁz���5�Hk��D`�����R�W�	����"T@`Zӱ�і}F����ca��dT� "���և���`H^�k��=؈Mp%�e�b-��� D�-+�17y �\dÏS�@��FV"Y0���������'�:�}a[�;�7��ՒW��0=�wĚ�S/�bH��b\α"�&7ђ+����8N�������'�����?4�Z\�R@�R1�΅��7�v?�(��,a
h�1�?AŒo����"j7q�0p���V>S��&�\[�W��Z�Ŗb�h>�}��_�,߃�Kx&:9������M�?��^���Ş����$��y��w$gwZfȾ�4grkA���^�3Q�8������i������ј�K�P	�'��2�������\��������p�WEI3��m�)hb�0g���0j%�R�o�׸���K�0�b�,j�n<є~+0쳄����>h�C��<���0���ޚD24�0�{�z����U�9+bK�3����h{Y[�3X�I�|:z�!e%��n��.��8Gih�/X����Z�����2�W�
,�E�pe�� -=L �W�`��#D�ᜣQ���B�W%�`��L�tg:Ťz8�FN/��o����^&Zt��΃�-}%���|�����SXb�JhĂO�hς(�e��ˋ��f$���=Մ����MD\7s:��?�
�s�L�<s>�ҟ�6� �7l0Y����@��ͪ���=�i[PX8�7[�<�=�ld_��^J�S��j�̈�:�^��,k�(��E^�kEo(�V�o�q��4��ZRO!��l�	�Q5�,?G_)N(�r�e�K5��hѶ
. ���8���������b����H��q���I�9;qL��}��8�?��z͚-|�`�(�e��WnO�
XťJ�`r#�Q=U����+$�ں
$_���EQ�pz&P��SaN�Ȱs���D������a(\�.�	Z��K�p��x��\�	��h�߷k�01���E��6̗	CR�QUNL�j<������W��8<��E:�Ιe��e_J��R~[=�/�L�ʪJ\�m�P�ǢD�]Mı�&�¹�	�l�@a�g�1� �.��	%����T��#�e��G֯O~�1z��N�I�$��	���6u/�S3�ɠ(0>��=[�@�q�f^�UL�M�Y�hK_&�4�r�M����C)S��?�u8�m:�����cU�WὣJ�mlq:�9��=@�t�k���Mu{����ܡ�|�&�_�G'��5	�wpi&�ទl�00`5K�[������'�	��l��c�k�\m&i�g��^G~A��p@��+�Wz�A�c��)����?��Y��˹�u;��I\�K@F���(0��G*�)V ���u�"B���
�L��eˤ('��4�C�#_GWn?������#}�9{@�(���Y^��AoI������V'� ��gН�Vj����4Y#SЙ�N��*�� ����2@�~eөg�N�s�6I�*/B'yNy�q�c�z̟/���yѦS���4|��R��y��P!x�^�=HG@Č��ߨ���{K��PƕJ\3�vQ�_����|��# ����Q7��3���{F+c� ?'�
�h�Ոa��I�s��e %����hYj���-0`�iA*��!�RM��<dVX3b��Yr�_v�}]��=KD���^Sf�hU�|i���~��ֈl_�����+��r�f�`�巐��:������ms��1M��Du`�q������O\@[��)�[.h�"Y}��������.�f���T|�E*�pss����&�]/�}9�jv����P���!�\h��=#r�]t��b��0�|�7�EK���׹O�-h�J:w�����j�Fh�(qp0�]R�Q�
���C��Ý�E-_q�;��-|�ܔ�+��^Iw��&8��SX�ȟ�7o˄]j��j��/`��~b�Y�t	���A#ޠ&`Q������k1��*|-����h���d�]c�c���v�n�χ<�摙@T6����o'�	R���s�և�s3���v(����Y5������:�m��I�?_�̲Ղ[��-,n�������d���.��$|Wך�E�P�]��x�� O"5�7�n�4Ѕ��tz@�	��3�C���R��C�#O���U�:�l��ɳ�A��r8Abcv/v8J-����� '9���v�L�HJ��t�,k���g�00��.��
���jưU��2�kLe5��J��s�C���qfB�EǸ�q��W��k)[�}�!'�G߂���E
���CI*��ʟM���v1��D/� C�C�#OC�fsI|��Jպ��U��'͜,��)?�e�x�r:�ح�h|Z�9��;���R�"����>>��|t�Gq�
O�S� �hq��*E�����/W�N�0Ͱ]�O�,���#rפ>�g��Z%8"����<u��e�Jޝ��
R��G/������S��o��zxX���lz��E�WD�?Ѡ3��"<ΒC��|�<�A����=�Q�c�g��̏��u��Ⱥ d���2�~"�c���3��z��lK�6�N�\���ic�Ȓ�{ץFc75Auh��V@���:��۟������޳X����Wm�;���f�� ��`�yoX��n�J���'�h��,eZ}��<y��� K�%�����@�cᘲ�3��)��$� �67���iGqrA���M�?0����@��/8����dh��J���:�Cp7H���Q��wd�J�k�Ɖ��\�cf
AP�ٗ�ш^��s
�G�F����-R_�
��������2���"!tw��"1�#[� fn��L������X�9���2�U-Y��Y2��m��pRMH���-Di�q�`��,���C�� .�a��y�]���\{���2s�U	aU.2��-����<dJ�6�)5���n�&���J��.㤼{Gg+g�2�[�u� ��z��dff�xyE[A��4�$/%�\��f/@0�i~9�	�������b�ߒ�����	u���X��G,m��H��%߆�v�%�u���r^�Z\��|C�BU�2����a��G6�	Z�tR����K"��|���X�F�az]�aZ�g�:���	%�v�4�?o>����Q�M��H%�=��9uT�٦m�$/�AFN��"�$4� _��
v炁���[�>zm�6�m��Cl;�����x��s���F@u�}~y�E?�ߡ���ѝ���O���5�D(�ÕV;�2���-7�sq�Y��W}��V6v��ֲ���d/�����_�����`�b�y���%��x�1����^���:�(Kg�#��A���@����d� �y��`n�����{�&��Nf��#��r�$�_\l���V��7ڎ�۽x�>5�
�oX�;#9�� �Ǚ�&Za�6P;t��S=�k �\�v�+��c֕oq���nL��T��aֱ��8��3��d�m(��%��v_�Eڛ�H���܍A�1��5��f���l�\4U���oo�6�4����F<� ������u1��P�V3��n^%yGKc�T�����^K�^�l&`�T:�*J�����U��Y��^�=���T!g�@�U�.����'��+>u�����]9U�|]cT�ǡ��@f|Rm��*���+�ӌQ�w/B�3�m�ߖ�v"
;��&1=�P��ę��V�S^��L����������4�����`پ[~@�0�
ڣ,�w���<��Y���Z�2�O����ge�@�s�ؗ�J嶛��\-�&���W*�:����m%y��G�9���԰	���oP��3#�H[�}l����v.D�F��_�M�"��;pS�l�N���H*nP���S��+��[Ѣh'�{��InQ�7����P݋���G�6�.NlX�֛4�6t�J�&T(���{��M]���O*��C�ZڹP�PO����O��M����ڜ;�}���|sgt�A.}_�	G�v���_mA i�d_��?��'��LQrJ�ⲵ���
�p~�3�
�J�x�O?sx�3�ðe����007�&3�\��%�矺�pV��;iV)���
�^��y���M���֟|x�7���ݲ�x�h�`��rs�i�v�c�۳H����,p���=�(u�o,�Pv ��d��x��\����(f�{����䨏Q2i��u���%O.�c��*�Ah�K�#Ѻ���_�2k�6����\�Չ�ܺ<g�����g�����`��6�!c_�ԅ}@�ʋdY������vM$z
j�N�wik�4�9�����A5__�%P�$`m[���������s�G��(����n����'�8��|����\#�x��#4E(���_� �����颓M��ORxA�LE4�E�p9��y@�"ÓJ��Y���\q�}V��[!K`�tt�3`�$��$�~�^�
r��0Ӎ������*h77'�[�T��g5}mܯ�����1j&�����m~�	�Y�Yj���u�L�2�R9=��;y�3�)~��@�c^p��TsR.thh�����8��]��sf2�lg��tp�4�,s�r��L�C+7뙊��<j�	�x�S�,�V��$�Ia���E�(0��y&�=a�d�$�`�m�i�扦�,�����9k���1t�����zi�)�h��U���o�+�V#���w��͜$^a���nM�G�Al��o��\v��~#��Yv����8 �>��2�*��C���jDWi^�S�کJz��:���S���j#���"+��/��ڄ¤��? ����԰�ۥ3�pq	ߜ����\��ٹ'ƅV�2}��ƨ�:݈5ҭ��~�j�4=΍V��,+WՏ,^�+-E)��',k=��\핉sW�ӅTY�$J������*�Zm����n�����$a)5"Ra�T�� P�%:F��)���e��:9 F$;�:�{�թ\�����	��g=��y>#�(��ҝ���\��񼂐!�{�]l(�E�ϫT�O�ԇ��A2n�}{2��ץ�m���U�p_$���j��߻yW�,�Z�>1�e)u�z��`����������Y�S�Y?�U\n�Tf�ֳh�h�iY� �y^S쳐��ۧ�	�"uCK ��Rz��������Y1("n�����r)�7�F���puD�jg v��G �ME֧�蟮^%–R�w�p���K��1�zb'��lN�l�&�����fh�|	oGk��K9.���~u�$�9��bσG)GQ�\F��qٔ�o"e&�dQ�֗�?Y�/�A�Თ�ֈG����9��^3Y���-���$1ay��(�X���QX�*K:�#�Β�AĽ7��w����X�Ɖ�vգ�P��N��пW��q��As\����r�r�D�^=����1%�I`{�S)��&��%������M�;��;���t�^�`�1C�a�S��wA>�,�̩�9��ya����\�G"z�V��r[	��0��h`P��{ş�b�ƺ��z�nΙ~m���C)x��/z��wl��֪='��ԇ�Aę����척O5�b��������ki�h�i��7[�;k8�p(����3f=����s,/D�]FpРN�`nFNKB�������m2$=�����S`Y��3�K-��X眯�M5�i!�3+�ݎnRW4��am����6-l��\,��x���u��:��K9��.��Y���r�rcxGlP�G0�Y�����j������G?��4�WN�9|�*�_Z��P�71��	�lU.��d^Y���%�{���Vt�����wQ?r�^�4 	�u���葬�&���Z2�pZ	5*����#D/+w��%�1��+�]�;=<�oi�}%l=��L�PLW,�Y��qC!Y�:�.��S>3��dO���Lz�T�,�z���4��H�.cGe�]9�i���O;��y�0r"�v.��L�Z+�����Lw�jx�B	
�y K^�g*�w<�)�����1�b���sa�"^��DT$&%�Q�|S��;��s�9���S�"�'7訏���(:5�3����Os0s�d��יEmR9L�tp�m���!���ERR��7C��w9I[�| ����	U%�z��L3�+��p%�#C:p�5T�+	H�s����u~쫎��Ǚ�А ���ٞ�[���E�*�e�v�Ub��W�������)�N>�0��#� �%[�>}���/)�aH��끤6�O`�F����h/�WM2��{ѐ?Z���5��2TNS���X̾����2�<3�HH��5�蜨�ՠ0Ҹ/z�j�-v�h�N��$��*>q�Q�&υ�d��5��uU�%9��A�}��:�����^<��%q':1�ǉEY�g�������B,�d9��g���{��b����D�#v5luq�o��p��j�zu���GQ 9��^���1N�P�R��
sM��8A_RNu���,
�O#g(�j�c٠a�%k����%n��Ս9�SOx��CTî=�V%��O������a�y���>��;!���8M�=��c�,����|m�IHO6�fP hdA�v0 �YUJ����Igk'x�Fy7Y0�v����#�����w�KGY��+�����L��j��_�������ITc�n�ग�i������g�ʗ�s�Q~O�j��˵��M�Ƨ�M�&�&�� �홶ڱ1�%��1�H��iF�H���+���O�W�ZV5����"�j:��91���G{��n����{E'�:�L9�Nv��t��o2�#���lQ�_l�,��d���5҇U��Dp��П֜��7�G��b��փR�OMO�	��>�໹��]|c�+���4Z�8V��2�S���t����t���)��-���M�]�ܭ�xr��Wݎ�Uqu�XN���GRf�"���qFE���˼��Q�u׿���s^�2��}"���G��`���M��ajH�"G'��j2�!vff�OYЫ	��/ƣ�Cb*��Z����q�<Rƾ��oƉ��q�<�gbY��?�k�e��~II�4�%U�QK8�D�:˳��<@Ҕ�4�[�~���x���Ƣٔ���^��C�'�����j�"�$_�P���Fh`����8_B2Yh����
$O!������E�Mz��n/Nbi5��.��	�P{��͌�	v �Kb�0�u��jVCЉ�]V�'� ��=�Q=��˕��m+nk����]�ҩaR�L��YVe``{D�^z�x���M�Rj�[�~� �z��#$Y	�ڰ�-`(B�i��� ��
l���lZ���ڍ:7��r� �:�l�P�C�`r����N��,��V��u��(z�kJT���8��=5�8���ȏ:������[�c0�5�A��"dJL/��k�Nt�y��?�m�ad<nJ�V��2It�@���<g��'�<lD��Q���%1{��Ȩ?p'r�t������6��̅��X�yd�bw�W�2d����[�5���klI�M������˰8�V4��Zeg��*?�ibK!o�y����[c�X� 	ZΓ �
2PJ�ӹ�I�-�|KE�Az�<�;�t��6O����c?@�W�"{�7�U��@�S�D��%
@���X"q���ix���u��Xש����P����º�}�ӵ�46_�i�X��h�/��輠�%t�m#���_�F�)	���k��17ҥ���*�X.R��V c�t�QӸ�b�i�H�\ydQ��y�yv�����$��%k��:D�Æ^U8(	�HMKp�O���Թ����w{�aNMP[��	՝����EV�m�t3�c3�p��3oJ���UZ��M�̀�����X�͵�a��:�mFxe���oDhX"T���&GF���������C�����ա)���l�фK�l�_���"^�n�Uie(�ne�!�.�O�@�@���n�8(���*[Ǡ��=���n=����n��h�IYE�$�b�
�p����dEԄ�).�^�h��-n�Tn�ָ���ڵ�@���a>G�xBR�5��,H1�p�P3K{�0qt����;���/��W��	y4or����@��p�l	�	S��)dm2k;������`!����p<����o�$`�S�����jZ�h�h\�:�;�7�����~%,=��q9F�
-����7����zq [�]�76��O���b�3�3f���wC&?S_(ؗ��X��kw/	���S���A�l��p��ė�u1���2.�qUZ;���brO�G��� ��������!7&�;��_�>IAA��2a5�c�g�x��[�T�tts k�h���
	�Z�tXP�<$�ϋ�`�˚�ŗĻ���'~  ц�iHV���U�Baj�o��C��Fbm������^pf���2l8�����j����5D���lK�����d�Y�C6 ��g����Dڨ_��1���3�,j������ؕ6�G��ݒGށ(��k%j#L��?�|�+3��]C�-�=���O�*t@���Mp\3�H �^Ӷ�K���E#D�����M���%=���j�WM�O(��%����>ze�ϕ�/ �+Ln���^07�ZRg�\4��ɾx�j�P:�l�YG����d�aj.>� �4� 6�K{Kc��d��
c�~z�~�-2�?�g�2r7�`�R�d.�[�*A0!�M{�9���O�o^-�鐾����y�b�x��8�%�fl��1M��i��㛭��$jO��ɚ��~�*8�8Vs���.m�y�s�&6�jM�j\=JJ2���N�:��l���j��#cڊ�} c���������?ų��JE)���c|R*j��leyH��)������:�h������
B���G����g�Öo�\U9OE��}��ƻ���u�����"���V�1�&�9]@��z?2a�AI���f96�2�*)o�b�����[oFҢ�Uom�0�9f;�Ҧ����<�G�Ѡ`��M]�[ �s��rW��C�q��J�D����1y7ݰ��1�Z���x�>�t�Āj�-���m��vֽ�����)gؿ6����K���{j��	J�0���$�s�e�&ے :�����IQ���a�L�
iO?��d9�E��Ul�ܺ�N��9h/G+.ɜ&,����s
z��ɛ�'?Ba��e�_�+�@�˝t�-�w�o���v��h�O��N�[��'��؏Q��0lu�}3�$(������s6W��j���XɽN*B2*=����ա�I�?�wNA���4�5EE�4�1~��j0P�TV(즕=�@���:8(�.Y7�@-Z���D4=�+�W��V�G_P�2C]�r?}q�gѽ��(��b�~`X�qq��?Be�\������h�����FL�\��%��{�`d����f�&�^��K���;�fVj�wö��3�"<9���=A���ucٲ����&����ld`����0$��ןm7�9�w�8��殇����6P���9�����L[��N
D�;��qV�]�&��	}y��Z�.���3g��9!��u<%��]�~HSů��g�[��l� ���)��i���C��ͻg�����	$G��������G�2^]�7i���x�\�!�"7['�-$�������쫌��d:�(��e���_�d�$�o���0@��7k�R^�[�Q�ei��qBg<g+#�����\��4+�M7��ڃ�VWV0��Sp��'�M[�;
C*�PcUp2�#�n�7���Í��4͗��V���ky�1S����)�T�+p{[S��N�'*?9x�¢��1�(�liO��q��*����u�k�/���j���ʚ�plkEwąp}a�PD���}�Z���a� �X� v���"�P� �Tr�ơ@N�#�1��]�;e�*��˲��0�?�I�DZ`���b� :�Z�?:l;7<��6���d)��M����@<WM�����{'�"J |�6z�P
(�?�n�=8�^L��݀;`Q�r�՘�ƈr�a�����;�6��ٍɻ�`�)�J���1���8y
q��F�)�P�T�tG»n����q{��u�3jb�jy�nчb(���?
|F�����dx��˧��2�iF6��Q>Vϴ L!��`fc��o;iA4 yۮEЦ�<sa����)��񋩴�B�� 1ibçù�t�~��T}{���t���j6&��sR?w��%;F��
���7ۋ�F2�_x�7Neg[i_-�_���I��1�@�����y��ڸk<����&k��Y�\8Y��.�������a�^/a'X+�!�+�|q{�I�� �f$��*�h`�� 7Y	T#m%�/PLW��R�d������$�� ��oK?P��K�k<�L��Mi�i-�7 ��L���P�柬�~��+(�t/���#��%R��R����I��$�=���S��Ϭ�"���彮�Ǎ��Ǜ�N;_�L+���͛&��|�\��䳒d>��.n�H��vtUI����`x��њ�M}ԃγ���G����=@�ز�-�'R�]�U�p`4��Tz٘�`;Pî����FB��&5*8Z���[k�D��(�Ju$��u�I{�mM�^�C��x9s,���H����9�x���G��Y6�®�i��
Q�~�1�->��=\��6��!f���2
r�jM��X{�:rX����)1Pԡ2�<:6�+|\��)��vJ��;zSC6��v��&Z��s�;=a��ZGR�pz�A�_;l�R�<C�æ��}d6T�N�'�gi�W3R@Ȓ��3���		��2�]� �K�@�~�Z} ��xſhz�n���&%cD��,� �׀���0X�LPX�CvQ�\E��gfM�M樰� +G
�t�^��l�O�ޓ+�w�E�Q���J�<��鿠� (�&�����cB�N��偡qrC�� �tHh�έ�.��S:%��-9w� �h��Q��Z��ƾ�!/�n	�ѫ>#�J���E�q�L�T�b�Xc�N�$:A�xG�p��	T�m�<h׶�LÁ�������=�b/�S��n�(�Δ4� ��2��`=?�������p�����J���Dؚ�a��b�aW&����Yęlk�%Y�=ʂv��~MD=@�'�͠���y)�@;J�޷�Ǒm���#������H����Ձ:C��r.��=L�L٥��	���� ��=,^��W���+r�c��s�����6ɉ��<��D+RW��V�w�Y�_��	��zZdP����/I.��BiaɃ?��G��).�o�%o\������a�n�p��#\&�G^�m'zQA���:��Cn�������!2ka��#�8�\�X���R���Q��%$��FO�HF�X��l>ck�����������a<�m�q�'Ah<H��0�U�N��MTX��9g6f�o�IV�c�fP��dx�9{q9A�7:��S*{&x�8��[�Bb>%�[Ϗo���J���I�+�d�WM�5�8��?D߱|��B�v$7_���>iq:H���s\�{�*8�}�o_��r�,�sn�g}:�gѓ�:Rh�����QH�����>k�TW��fN2�2_=���x<�{��q�y��d��j!��W&K�-��
�{�m!L�,p2kg�åJ��3S�m�[�2��9�:����U"��3Cɗ�?��i;_̖�^�t����s�E[�A7B�H���(\}�l\��\vZZ[:.?_M�O�d����E�6�_qܴF��u*�iags�LPs���p�U[��K�nL?;|���q@���u��um,�#|�(9�ݻN��Do	,y��{#q�����R���P�X�K���C;�����L��<�.��p�(E�P\t��\��/z ��!����%{4!�/C��]��t�yWl%$�| M�K��?	#������SM׃GZ�Z:����(r��5]Z�i����6���� � o�����:?�|����D�<\��p�H�.�4�u8�^��'��渏�@ZBF�;V�y��q3�<���c<4x��4��o.�6�m6m�K�@)B�� �mgU� ZC�P�`ͦ��捫[Ɣ�Yi^U��l
g�x�ۥ����\!�H�+EI5���<��!4|���ORv����c��)+�~K��63{�*� �0՚K�n�52��Y���:%%�;ơi�.��cyw+��>4��������)"N��� m��p}���׬�:���n��7A�j���@2(��Acs3�M1k^�L!�n����n���Y`b�D{3BuҺA�Q#��r'&Cs�G{R�K.�z�s������~73�OB��8|�� q2�F��|8b�K���;��B�E��;�FExńQ$�Mԗ7a�7O�,FC!f���Ɲ"�Rn@�6��LMZ���T��D���\O)�Ɵ0�C�<�u���΍�kwG3-�=�H �]硇������7��4����<.����ښ3��O�ESr�t�M��`�"m��H��e¬�4�ql�5�y��,�:g��_�-�=�	���*n�^#��z{�BEޡQ�5T�%@-9�k�}�<mS�.*w�!��g��!+UP�ק�:�m��g7,O@W^|Z��8��?��u�9��O�IW��k����lu�q?�����	Q��hU��Z�e֢��~�~�:�h�t��ٽ;����d#k�|�'v��T��
�YpP���Y�(���êC�s!��y���
�,�S#].���g��[ �����o�e+�)���$/��Nn��-U�U���xeQ�'�WL���4����Y	�|Hm샄Y��UI�6�!F��{l��f/����ɋL�e������(#~������)����]�8��X�Ć��3�6���Y�����4��U�D+ڵ�˝+
�]�N�wR��/h�`R�u?Ul�jh<�����#�A��K {�� ��@�K\����gz.Q\j� ��{�:�-)y��v��j0q�HW�i�D�#�h�C�/��U'@ٷ�h�s]N�a9�l'�3E�y.�}�E �I��~��Yd\��N�TJ6-{]�Q��w��*������Mʀ՘O&�l�N�*A��/e�t�����cG��Z�*#7i:�����j4�  �?[�� ���рq�"��z����6 �(vD'K1��n|�,Ra�sJ�I�l�b�0�L�K���R�7��������@���3����R4�9i�*[h��
��L.�M<� u���.@c�uH[JAJ��/r�"E!(=YdH�a�2SF�_�t�w�K��0��)��6E���8�<�fӴ�$ �H�������8����b��RBD�M����(�r:��e�9��5���t	��y��+&��3b��Oxm[0[O�׽{�"�si1������r�������b�
��&a��T�EZ��s�L�0�k8�#��B�~���v�ܟ}��i�ՑqD�u�2Z1�VCk�.�S{�x9wep.%ι�"�ʞ�w&ڤ��;���&�-(n��z�G%뒕���15�O횰���=�d��ߡ	I�⪺>�.�	��Qg���=����M�x��3���M=���p��
S@>�W�C�?�S��F�btpS1�M�F���=��fzsS�������k�#+3
%�ҕȏJ�KqQ:_�S�E(�gS���L}�6�"H̗}�!�W
8]���n"�,~�<N�e��ް;�u��}S4�]2�e�rS��x4ϴ"80rQ��|�$�E��qw��M��ʿ�����Q����D���� k�ů�7r��Pv�:�Q��y36�뮡�,i�j���(K��=�?%o�*5Ç�B�e��tf�5y69��q�N��O���7p�BF���Y�@Sj��nD�4�[��ݚ҇}|�:�
ɌK�O,|��A��ou}nřD^�� �ܜ�ɰ���'T���������LS�F�a��c� �]�0&VL��(~�f�Wi�h�t2�)��s���-�j�zV�d��*��K�1����	��rk��:E��c�TZܻR�3%�}��s��,�������8�xc{	c�$����n_P[�8��Uƛ���lNnD���y�9���F#�D��(TeZ���H��q+ip��������
pU)��J�T~�����>A���Ŵ !TY^��J�1������B`^�F@}n�Ԓ��H�a�k�㲑jFm���с4��K��'��$��4��!G����qg�XX��H:(������pj���;��@<�]2ܾ(q�3>V�����`�1_��3���^�4Q��0�Y��j��o	�V�֫3r�9��hαJ�v��h��\j����_��.���� �$@���F�}�9��S��F:�2�U�6v�"��!,��+�������PE�� /7�D�.��8_A��ߨ��G���5]7� -e`."�ۮY�ݱ��X,��r���%ǼU���խ{q��9��Ʈ���Ф9�����ˡ��bB�/�R�=O]��@6#�s�¢A}`��BR����'��b���f�t5l���K�9`�s'A0.j������,��f��&(�;������5Ʋ>L�d�bb���R�L�Ψl�	'� �O������z5K�`��BҀ,�a,2p�@(��kC��:#["��Mļ�g�����B�l��Rq[����F��52MW�9<�"Hv��T�C�7.���_��Wh���g幨�0lxu����b�^jb;^�ك�-8��&��M�SǎI�������;KB�MqЦ))Ĝ��9=h��%��C�Ş]>�W�6.ӫ�%M�U8��i{.<���乑yv��㕷$X� ��Ԗ��-�I��W�p�9�TUDo)t�Jp�$�^������n�.n��nB+Ԧ��a�<U��e����T�6y՛;]&bp��������<C��ؔ��BnO�E�7�w�$��1��7�D�9�X���� �2v#�W� i�Ҽ�ޱr��ݗ�{�)��ƅ8���AhI�<J�%�f�����$&m��6n�#[A~"�Hb!�4p��Rc
R$�! �j�^B���������)�lr�'ڬ�\w���vrSڲ��/��QG�iM��à]>R�;b@$\���{�˟~��mɹQ��O�6S���Pc�Z���2G)����Op��z�YЪ�D����Q�z1[���k�k�Ӿ�썂�}q/j��5v�Z����oS�p�3cä����`��+A>��q��
9�9�no> ��5)oY�s,�=Su1��6����ļ�����U��c�y�Ё�LSr�.�B�=��ƅ�5�CYa	�^-���9���f�[�}T'�|�-<���i7�-��|��`1����Ul�	��^�gz�P��t2Dt���UO\�U�K��(��IR]��a��竮<�?5�6�j�0P�%��Z���Ϙ���=���pz_:ZhC9�����kyZ��ꁀ��de�{!��tI�t�
�Ǌ��(�2�s�"L�5�����փ��Ҋ�����?�݅$N��5h  ��)��1K�e|\j���#T�d�m�6a6��usBf�(������01W.Vz��a�����ƥ������U����;G>����98EdN�ӗ\����e�'�``�n3׭�0�uj�9~��ۈN�f<u�(F���O�l��
�! T狉pO��2G8��2��ÏoR����z�KC�Ag���?��ϵ�]W�N4�Q��h�����<"G&�s�w�4�鉶���]	2�"���3?�i��p7��A�mCC����=Q.��M��*6�3<�%���ͣn�sO6�e���EV��&Vr=��x����=K#���Xl�n_@Ѵ�_˾���`|@�(��AR61�r�(�pxv��^�Y(He=\�8�:��cl�7'��19؎���k��r��%)�)�(�����(���rP��id<��֕���'w��N�P�|����DTr�?��k+�e��C���dU��#����xah���Jm���~Iz'>��w�+7�i˅*8����'^���v��4�Nz��Y�Xo0������{q�uʖPnUϤ�E�����&���_�С���;�º[&��?MF��΄��;�=9k���k��2~�އ�?BƎ�V�2_G�'(��~�G=��a,Z+�?��Pg.�/�ݙI�Y!�`�� ����T�J�F����U�{ߵD	���m�6�_�����잦l�C���d,I������#�ud��0��K[gF�h&�+H�>��|
 i�v�cs�U��3�T�p��хt��'�P�eIs��:�#ŬI�u�n
�F��~nf�ä�i��H8U/�z�)�y���j8�/Nlx��J.(y�>i?��g�9�֪\�����A.�u����!q��1mf�'բ.}�?��5<AbG��`���{vy��ƚ�K�g��-$�]iU�e�8��(p��&�dV����mYMϴ�9��?�@��T�?��Q���켯y�%vE���Y�~?Q�q�*���z�$�q�Tb�> }��K�>��6�	%8�D�5'��$~�ae�;*���t�y*�z����W=�WK6�ZK��W����\o9���<��J)R�v΁F?DD����r���`�#�K`J��*����`k�ц�>��%��L	D��_�KD�e�|�V��;���l�ڏ������m6��3���={���͎1N��	�#��D�q�- c"6pt���%�!}��y��=z}Pڗk,�:�נ�ih����pn�f�����ř�t�qJ!��[�)�w���O�V��ޣ/����񛸷p�o��Ӡ��O[�`'A�6b2}L#�0���[�j���s3�_
�}�\����j���kT��5�a�;�� ���x�`ay_QD}����u���J����DmA-"9 ��Z���*:{��O���[��̈fB�J�x���Wg�)��,�>3̀�[��[����[o���u��3]����f�omn,ǿ����XT&~�9���<��=^��J((����3G�5I7fn6[}[�I��-,'_u��Yх���Ϫ�,_�wRj����U��]>��u�ٶ���� e- �N�M�)�ɡ�6Z�>6�G�]w���oE)_c��n��UbX����|u��hK�kT��f�:x��z�8��Q,��))��q=��R�^�	�qϞM��R��>eZ�p�1��aR�������vT��t��U�#�m�R��H�I�!~��)�*=���`�gE��}"��I	�1O?%-��G|�9���-BB���4�s9(�YAq�BJ3��H)�B7S$��4D���
�ة�Sn#������ERk�a"�u���n:lӨ�֌lLk a���%�aC�>x�������S~��s�|�z���9w���;[�Jf�q��F���P[/ɘ��=��~�4^�R?NOHƆ��YQ�tI��Կ�е/�Ma���[�e�9�H��In�I�֦hw�e0 ��SO,9as$h�g$t�� ��{�;��4|,�k�j��Gz�N9z�!����I���� �X�P5��#O���}d)0]���d���k�̐���Z��며8��e���ΰt��2��&/����� Y���ڳ�t'�z�6c?��2h9}+�Jw���h��}0 JA�whLe�����^��p���ΊmM�N���Z�$�1gE.���I��8���?��zy,�u86����F����7�E��T�Z4t�r�X���-K�p��O`h�� ��#��]C�]��PV!���,+*)��A運Q���7�N����!�b���4s&���~O�$oD�a�s̎FO/��g4i�n=I+�|x;	{����x׏')�c5��9������uLMh��B��j��:'-ţƣYA��r��`wj�����"��z=sKIk�CU�V�i�?�*=�5��"k�'k%Hq�N��]܀�(��[��K�w�A���i���!v�0܂�C�O�j��*���T�2��Y�o��3E��(� �p��4���FA��c�vw�0R�����E㏏/�e��ml��5
���1��@���iu	bR(�6I�`Jq���^��^��X�VR��D�5I�Y�P���t�)c��O*r�>�ηo���6E���yP�{��9g��@�⌇�M	�
i���68xa��PaL�τ�73�_s���3/c.Mvh�M0}��'�3< ���
�]�)2�zxe��� F������=�Y|9��ۤf�����7�U�f���g�bx`$/5~K|nG�o��Ț�C��8*T��*ɏ�վ��.t�v��7G zq�3�	��Ť� lbPy�	���'n��_�R[!B�'�;�r@U�ж/�~�h�]e1����1�u�V/ʂ~q��Hi�r�FF6MK=��v��R�5�� 'QJ�#�#�����Wy�%����79���g:�X�vk� {Tevq��������y¼|x1K�ꂜ}����
ի՟=�<��bv�d�D�틔[y̷�|�G��&�Z
	��u�
�������/k���^"��k�0w=��*K�E~ʮ��e�?�͊��d�cuy���ƽ��8�Ӥ����3�{h�꣢f���,q"�u��m.����i����ۏ�^����e�a$X �]�Ц��!��M��v�@���Ju�M[_�Fn?l%Y�D�"
u��q=��x+����Ǖ׫�V^)������_/�i)�#����us�(���C�'Y%�<'���XO���d���!�5d�چ�����	� �~c^��)��-�v�:���Sd�=5�@��L�ܫ����G��p|7/[��;��,���?vxD���|����kv����ƍa}�v�9J��W�h��j|�NX���y�z���?�Z	��7E�����\�:����G]�(R���"�x�,yɨ��c|�	9�V3��h7T����6Dz�0D
5*R?��3փ����lC�Z��o�u��&e��J�N3�{Mn���~E�ɨ�!Tj�9x0y��.�N��~L�Ȯ��d�X{�p 
h�|�	^���$����� (�u1bd���b%٫��Tu��!�9�q�1��)-|����C��� �(|-	�����$�= ���f���W�g�$Md�U��h"Ţ���=��,ժ�a&J���ͼ����yF�|r(b�ҷhn8�gH�LXR-�ê�<�/{�b�|Z���6ﶻ}�\��p3R��l�}eVG��4:�~`Қ]��Q���iI��'f�����	M���8$�]��dK�Տ��@��$�O)^��wO1����U��=�A=�`�\O�c&5WN{	���=M� 2�G�J�%���P��� �K�� ��@o�%�V�C���f)���4��>-l#E�[,�p��S���YS�'*���P�Q����Y��N{բ����,�y��aR'$;�T��z̦�@�Ц��yZ�;���e�xl'�huI�zЫ��&�^CLh�/Y]e��Zb����rF5�8�Vi��"Fڞ��1 #�0����Gߣg{H��6�Uz�h4i��Qs�9������?�Y���"G�8wDH�7re�����.�L������)G�j�1Sr��J�7rzJ�¹�[ɰ�^̾pQ4�6s�a.�ςd��޸,J�g�5O��/c�3�6[6l���A��]J���3P�O�6z�^&�4Eg���:���{Y�̯ŝ�K��Nr|�8)���Ώְ����i:rN ����2��_���6�:���/�I2�!r�����zѤo��R�3�+?Xk���u��Ffk��-'1ރ({�%� �w����*�˖�����'��r�'��mV�s5ӏG�F�I ;V,7����E�G�lb\��*���}��9C�{\4Y}9��t�L�r]�R��FzZ";�h���1�/<�=Wh�����*���Aa�@T���b�e���+����&�P/����A�U����󞭊g;�Q��I�A�����upk��L����gSަ���2#�`��~�}� ��k>kó9�����E�d���di�Z|��T,���@w���^�U���P2�� Q�7��oZ�6��%���8��| c�;�Pv�Sg yP�e{�k���GBS�n�jlp������<A�-Y` �q�[;~�bsHD;�jQ+V&:n���	����Њ�F�V�e�������2�H2#x#���������Y93轥.�-�F�4R��؟H>s-a�`Uk^��/�x��5��7���@������)9�&jV��ǄY�t�~I"H����q��r`���L���k�'Dj����c<:����O1�вGބd�쇏D��l�>�Uq]���
�Q���d��舠�v�:Dv�8�b�W݆���!�Ŭ�����Zx��/������R2��$�`�G�i�7z�r�繀8ʯ�#�$3��vS�µm	���>k��O�ߠG�'��%�/Lnj�� 4�,Y7w� ��{��^�T1��	M��=��P�
��'*_2	�! [�lp�Êѧ�O��kV �z�	l�N�.Wq%<ɑ�;)�i{�D@�L�ߩF�?�)?�R�8#���q�<|�pL姥�����qn���G1��ak<8�����߰�z���W����En�.��Ⱥ���6{�ǿނGyg�-*����K��F�=Ūq�B�S�9;��oO�e�N�Ј-ȏ#��@DQ�67e[��8�#߿FV���ez;	�??,��2��%�EYc����*���V* ɴ<٦��S{�>n�ygz��H�c=����aβ�03V�������D�Anh�D�
���������pO��X$է���!�>��l-�f1\0j���~>�!ol�\5�I|t����)B��� l��cu�D�;B�+�<�	�Ҁ��ł��d�t3��Z���q�XW�?/A?G�)>�����W�%�u��R�P�kգ��/e�51���V�kB͏7:�cC[��]�K�|s�i�n8kh�2�bҀ&B�걤���ެH~L��h���h ��Z�ꗔc�yS��?�O�䵸kF�����w��t}�
�riKv段����1a�T��Qya�¼ޑ�4ڃ��o��;s-�I�p��YDb=;ԍ3�:��#���cT¢�V?/��|Wr;��p��zm�
��h�T.
7��NrDV +o��7 ��ƒY~�My�����V}�t|�Q��]���(�=�1��~f�I�q3@eb�HH��UӘԎ	ˈ.t���?*�D�Dn�]�aL���--hJ	2P�I��!,#�h;��A��� �N>5�l_���g�%��v��0�;���@1v�	㍘��Bg���T���ʀs;�bx� �}��3f� +�@�yrB�~�9`�B��vB�!�� oH��8Y-����!��ɿ�:�|d�6$��{��h_�i�0A�m����]�t�
0���j�Cd������N�.��0�z��` ,b'���1�G#*��WB�~^ys!5�se#�0�p޼�*��
=���#,5��B�O+?��p�G�-���o:�K�����m�w_e�B��G�g�:4}�s$]O�gM�j�v+�n������3�n����LjQ�J�N鵺n(��u����Ǆ�8���b��
�	_Z�%�:��u}\��p�Cj��G�te��k'����f]��B���a�~vń�e�Q-ɵ��wՠ�����I���+�C5���n;<��*��}ʺL\�dj�y[H�N�A�C�UMu-�9S��͸�lO!��NDH�.$i#��nb�t���}�oq�'Mx>��,.C>/�ihdBG����A<�v��ҁx��F��§�\݈;G�}��`�KJ�-��\R>ga��?:S�A�r3�Ѡ)lѠ}M@z�@!,L�����%���a�h�
#!~C������1�-�م��xz̤����\q`èh�j��-�{�^�9@.KY�X����\ `EO$�V2OP�0�Ce};`�k��*+5=0�Ls��D/�XQ�{6����@��)�dS�+�ۀ&���N"���]}%Yu�NΑ�H���ˆ՝��������àH������A�<[��C۩�*��ٻ`1��I�m��9�GǙ���vf~��e������U����?0EA|���C]��C�s�m��L�lu�_U�� ꟳg�ܪ�^��������E�6m�ޙ���3�1��LV�aw��j��%����,�|e@d�j�����N����d*���pֆh$ğ�����qa�%�O���pZ�:}7�8Dt#��C�\1�(3��w�#�*֟��5F�kU��iV�r=�R{-Ć�2�ׯ����^�gs]�kf��7�&�*~ۍ�Z�T8Z@����c2���q-�ǔg@�fgY�j7�)��V�h!N��S�\\�t�~�r4����ᵯdv��dօp���	<Z��(c�пw��/�v��߽@+ы�
F��˵�-�Nś�Y˪�&7U[��;�����n{��7L��Q�^K �Ӓ�=�-׵8�>*e�Ƶp���H@�&�	ോ��J�_xcTe'�!V��j�X�f��5�������rz1�ܭ+*���H�E��䳛w�@��T9��[,b�͗v�L#�$EW�9-�!9����{���p6��^قG6���mQdQ��yG:]�Y~��K���p�-! �Ǻ=�D�nd��� ����:�N�zAl6f��f� �̂Hjg��sta!DЉ���@+K�&�n}z�kB&��a.�~vݽm7 �V��c���w��@)���$��ہ��8����7���,�в6����f�R�V-��6�}s��k��!����A:-4�%�o`)�*]HV���r\�U:VL6�<�
��x�-��"�il��������9n�X�J[S��i�A���M]ؘs�o"aH��r�����J��\�
{��]ms�Z��e&��t�p��1�ǀcd��[�����&�H������tn����mfʂ��1��j��?(�=���1�lb�,F��θP�W��ޫ�V��dj��"�֪q� �6�"���#I�X6�E��@��9gi�{��w&�a���~�~}[$n�������@<]�N��?�M%iHV=! 
�^�wJ��:B��)�^��˫��s��`?U��\�=te������[^4��{��${��T��q�qn )i��	7 ��.I\��R��F��s�h�;6����^mނ�U5#�h��P�75�Mt/u"�$�+�ێ��]�d�I���z�QN�%��$�+	����E��J���G9~��mH�VQ��[�2�f!�K���&�V*s�#Zq�5�(9�����������$�h'ȗ�32���Ql4V��4M���;m����[ȱ�H3I�~�#$��<���&��&1Z��u7��@�v��{^WP^	��M<dZ�qWY�r~�};���
�M�Iy����4�`o{>؂� �d�5|�<͸"�:{�~2�� N��2j���Q>�K��mQl+��N`��ԁ�Þ��y<Γڍ|�se� '�7����>�.+�v�����ĺrLܷ�T�=L�w����M�1@nyRvY|BO5X^Yo��{��ntt@_��vu�z?e��q@&b����P=�\�2H ٣��B�5��tȷ?�������(%}KX�-;8�.��{Ԓ)җ<�WB��l4i�8kz�!4����*wM�}�y��C;ʭ9>T�p]�v����a�X#���W��j�7%�`B��j�YX�`D�0d�X?�c���G$e�}�t�"��9F�})��ȴ�]�M�}Z ��Z���>�6]Dt����z�?��c ��0 �IKaU���e�`)�\ �G_�=i�����à��س�3��m���L�ΐ��ʇ'�v�Ξ�D�nN�>4wA"�|2
$\"P/�N�vxe�Ĝ_ͮ�D���v�n�[��	}H�����Oi���ߒd7� �����������.DG.W,��!�Ƿf������� �:b�x@�k�O�FMhI;�a�j�4�cL!��N��m�5����FwLO��~�5a����"�&4h��0�,`(�Tb=�� �.��Y��34�
[�CxD�d�`wO7�����,��N�����u8R����W�.�- �{������vʘےv9����lV)(�i�O�ą�.���#F?����I���fv�H}�ub�P�}Y�S�>���e&��9ƾk�wϮ6��[��"��}��f�x�����!�!Y�9����_�P"�W����P_n�e�pL����F��q곜Qd<PF���6����bHܢ��8�|�+#��{�����H�(/(��ZF��H��c���ѩ��G�s�ZɎ�R7�k��<qk�M]���Su���Դ�� ����P�e�Y�-u�[��9���|Ά��l�1]u��;=�~��Tq�7����8���*�,/}CqBy�絈Ŭ� ����2����L#mj8� ���ƈ2}�GpQ�Z��Hp��H�����>�(%��\��O��ʛ�(a��3;�^�w�6)uQ�X�6�-N�c\Ͻv�|;/u��r����u0��M����������>3��acK�$����d�E咪#�i�(�͖�#��ޕ�N�A���jux�	ƨd�7U�w�;IQ1tg<���ʦ��v�K�semΑzT�7��sD���H�>9��m���w�G�~v�jC�v5�]Z�U��d6�ܾ�N�$�eB������4��|��<�A�m�Y�I�c�0�L��p�40��AE��'H)��4Ϥ�@���ԫn!����$(`�0�T�L^��j�������y�AzR����s�,�H�����^+���~[��݉�Q�0�����Üm�1*�|cձ%鼻�#�ΘQQ�[C�,�����{�Z�.lU'MF�"d� ���-H�UT�ܥP�}H#�`�W|5d�҂	��V�y�m-��ǋM��O����A��*��L���rJr�o_�s�S2oF�T^PFb#��i{�}bM�2�R*��P	:[��oܱtɦ:Q"l���QaRK	�{�h>���e���b@��U�tZf~&y�vͬ��s!ԣ%9�&��ZJ:��gp��8�q��N�OW��SBU���L���@]�	�o�jG# �m�oɝ�Nǭ0�b_�\��)e1]��7ᤉ�/�^�MVe���SO+�ܦy�x��,b�͹�#��v:�TJ�E4e�h��[(�����`)��M�����W���9�@r���A9s��J�G�Q��|�B��7�=l����i�^(�	�*�� �/9����g蠗VP�1�$�1��b�G���{W�ɫl�g����Ia䦡_��T6��G��u%����0�JS{W��#�!q̞�r���M>�H�<n57���O�{_(��!��x�X���*�e*`q��2���/䷾�Fs��p8T؆M*>��?�tس�W�`�!� O8 	��w����}�m���ѡ�����rШ�fN(��9�g[���U��wG8
�����\�TڭwJG����=;&}���e�U�hp�[̣&B�55�����s����yr=P��CS]n��)�����Mz�$�{B���o$����?�$w-,�]y�XMe��`�I��\]u�I��m>�Rt((g��A�A����b/�]��3Y��}�]'�8�C]��cf6:ly*��`4yN�fƨG�kn����
�0¤A��1TV��K
��!�Q)G���M��(I:��G1x�E�Pu���7]�x>�{=���(?�F�u�ka��h��G�-H5����R�Lߧd�;�!�̍E|���7s����s��To��P�+iH�s�f%��E�;f�E�e��}^r�cP���acy^�d�Yp�~JM��|��I��pR��	,ĊN[h�>1UR�[�^�st�x�8� B�)�ʢ��*L\v﷕�����4��,�5��栵�	DǏW���Ou8̋�њ�,����0��5�ZN�$
�n�*q/1�p��+:���Þ��x5�)#D P�O/���E4M��8�y�&p���&�17������p��׉ї@������Q�f�i��6�'IN���ZnuB�҃V�0˫B��'�p=e�����"�-��|��K�\�0X��RG-&Kߓ�����E2.��c;�8q���q(jbI��o ��i;�E�1��e�k|ڤV��{��A��hA���/[��DD�>��>j�\)���65�s�|^,΢@�=��H�w/C��/���Xrj�e��{��{����bE	��~\�A7�%[?uj'���歮���D����쮅U��Zx����@�+W9�H�g�C}���͙X�����=�D�9g	1�1��M�<qa,����:�G6��jU�J�y��9p4�5�� ��&?����i>�#y�M�I�XU[�|Oh�66�.��P�Rr/}n�V������<Ϻ'BN/�Я�To�僦��cUK���K.�-6Jj�{
'e|�$ �N�DV�5�'�_�@�Q�L����k�^��m��~�a�6+�=�^�:����ʧ8u�i��`fk�KQ9��4�N�q]��Z���(,(&u��}��"�ne���LO|X�@lrs>ήʳ_�b(K99�6=;wxJv���1�:���TA�|^� Z�4m�;1*�Q��3��&7��(��e���aR�}��\e�ܔ�:O�vK��0,�q:�%�ÿ���OR[4-��u���Ҍ��̟�`v�v�3R�^j�p	a�n����1�_P��+�]-YWƼ����I X�Ə�5���{78�%���;��s�@4ڄ`�T�c���/�Z�6�N���7��1#���e���t$� QQ,�iL/�H�㨎�I���Z �)���=Z��4�t��|��7�~�]��3-퉗K���c�b��cW�X�D�:�����f�|���_7x�=��`��U��y���钪���x��(逐����!��b�W�>z�&�О�,'�u6O@�������iҧ_̿�Q,/o�y�|?����V�P�Z�Z��T"���/-Dq���C��eC���3�:{|�ht��\G>@�K:�Ҩ�9����s@>�.���2z1�c����2ȼ_g��X�&ED�_X��[�.�˱���q��m>+��_t��CD�X�$��n��H���c��8�l�TX{�gcJdЀ7��$�KHm<1���S@��2���ޡ�����gi�l*���u���G&F��	����UZ����p�{n�R�j���9�J��S�W�6�Q�?l�����\եۆ�����6Eb(L�x9\�Y.�J����ݕ�/��,)�k��>�Yr:�T$ѦU&���\Ģ�z�17�4�;��������4��4���~��t�q���H6n�m_��'���#:\E�8r�;�"��M;L3����K�J��<t�3�ʅ�kX�}���BfD6�|��2Lz�m�:v߹_ps��zj�C%��)�_10Sd3�ac�"3�����Z�XV^�q�Lk���֎q}�L$�^�����߳��|�����"*�
a��d}ᰯ�	��fH����@ʩ9j��==QB<����=ykav��^�Th����8��j4�$І��mu)�"réB�q�h�I�M�+ �[���iå���'���<M���7�Z�K�)Z�n�⿓�h<ʥ���'�����nn?R���.�g������T��V~��p�b<��U"�PDm� ��֕{�ȡ:���cA(�\����ۮI4]4���
Z;��ރ;�̔Y���۱L�ߍ��Y�k\��:c��'o����%���d��fr�g�2��;�����H�����������#{r����ǜ�M@B)4x�?`/�AmO�$��^x²�Y\�#��g����?��-6 �*�����1�}}8��aM�!
j���sh%��Hyb��aA�z����ȩ��,o6s�ĐK�k�����5`oƷ%O��lݿ0������?V�̎s~�/FަED���̟���Q� >=���j�Yu<AvhC�!�y���HNm8��+���%�ґ>4�=�����>����n�蜾�����ǓFN��c6@W\/wg�_������6��ˤ'������x&[
u�|�XN_I�����������^�k�U84E;o�~>�S�	e�)&�O����T��pk����ɱAi����g@�b�E�p �ff�׭(^`!9��������P�a -/9��a7äU���l�*]_p]ߍ���|ظ�ħ�5�i9僬1x���hP����� �FD�{p؜I�:iBG�Y �����K�?���#�=��^���S0��2N_������4PR+�̶�a���55Q��EjOLAW�+�+�뙤0K��B�<��9���Xφ۽�JJ��D�Pe
o��?aI�Y@F|�諯���7L>E��E�� ���─�B�0g�x���$����ǅ:�����@���o`���s���}`��js���Aa���ƈK�bL��a�JF��ws�B��7\��� R��fI�"?1d�.rv;�v� �8��8�)�גE���qf��Y)����4	����@[�(l�O[9� �1����A2W@�}�7P9	��ryUm�ώ|�du�AxŔ]��d�wD�������?�CW��`���D�f��X3 3sf��2��.��&��A��:��x��J��O
�)i\�x$�)����S��^8�o�e����Kڭ��܍�F��f}ةKη��ϨIpY�z���z(G��\��i��!G�~��ynJ����E�w9������Ps�~~Q:5|����&]�%>��!;^'�t�1��/����7X�T��Ȱ��}�F�?L�;�����)n�C��=9�i��8ܶyG�'��<��)��tG}g�	\4yRq�L֏+#�_=��d��8�0���Z��H��X���}��
�k�9���"1.</��{ީ+߻�0��W`o���q�_��EÝ5`	�b.���тg%F�j"�z�ꆪ3�e�+Ȣ���n�BG�0p��ѣ��9���M�-~7rxR�/v��m+�6��pfb��t^d�Maϸ�uS�$r�p��|�@��S�<����GI�M-��|��#�w��e�ֱNH@�+L;6l�桄B��HfC�$z1k�L���EOM8?��~��1g?o]>�%�(.k��c%H�عP>�����/��h^���p��ˢ��x�E��ɋ��d�g��g-}W��-��W.Us�5�E�f!�z4V\��,��vH�9�3��b�ٳ��8�
��䤮!ո�բ��8_�}��ec���[lZs/�ck�O[� :cw��ѕ[��1���ϫ�T�7��ḣ+;�g���I���+��@hU>���H��%~���XW��J^H�Q�$3{�ѵ�����e>�)К�L��n�������KJ^N3*_�"ڨt�ۜz��7��A�W��z�j��*"�ӥ ���0nS��N���ڊE�ف�����	ኁպ+~�@�j!�a�=�3�e��g�UX���Y�q	%�Yk���b�$��Ǳ�+ԕ����Z����(̹��E=�X�Ŕ��.w1)��5���Q% ��|�a���轜ԓ��)I�