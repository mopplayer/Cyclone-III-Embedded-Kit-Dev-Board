��/  S����3�c�ub��_NЀP���t�,ï�!U;�P{�g��Oj*�x �*�'|�N�Q]/]l$�W�]@	�r��GT[���)O-�y��1E�����p+�b%Wq�d�MPFQ�����ty�>�WW��5�5�����5 ��؂��E5l֩+�.d�f�&c����/5�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�PM��1�,=�f��.bG� O������y
e��&�F#U��OWU-ܜ���-��~��]=�Q�q�� �'�'�[��[~^$g�3p�
�=r��lO����#��� J|h�(��PM;oΞ��EQ����G�� ���)�y������&<.�o�L��D�m������F���d��:`��Qj�A;w�XiO�F,���9S�͜���ȥx]����j��S,��4��|5�)�
Rw)���U7���e�-5���TQ� �d3�Kr?'�q
�95����I��,(v�V'h����Q�IG��Y$�v��|��������� �+�o��+6v.�s�=L�}x�h4�3����5�uP1�%3��y��׷�G�1�f=%M���Mɋ�s���c�F�I�J� _	y����"4�������/�`n�"X���K�r��	p���Qs[�>��!�54H!���v.CwN_zu����TXsi�W�c���{C^�_�X���P�t�@���j�����R�Yp��(�N���ytx���x#ݞ$ʡ�����	+�(��,��`"�M?KԪ%�2��"�df�b���
�G����a�ʔ ��cv���9U����)���_�!^�]��ҷ:�æ�1F���L��0��׆:��%�/��lU�̠�|�z�-��vm�檚�T����P!4�v�TTG�&�g�0�������6-�"��_l[L�����B�4�]$�s����i1G�C�M|��lIR���sv���	]�9u�/*�5ʵ $G�^���R����lx`��Pk��՘R�B��E`w��?Kj����u�{����͊���kI���n�S۫�	�:��6߅����V @�6�wöqu�[w���_�H�&�'AT��-R(�Q�I[*�9�a�lh�o���Z�L����,�d�B�E�r�`���7�	u١��׉�T�8]���	)���fR9��khz�wR����줲r���۩.�D�m�Fx�����)�M/$$��ag	Ei+�,��zX������F-J�y2�X�+�	��= ������b4#�������:������|av��Y<`�m�!�س��JI�0s�����J`Tϙ-S2 |�oHP$��������5�� �)�pDv���q�t�H�_*�=������[>j^k�H�	�(!�b��}���~�<R��޺JC׍����vr��&$�fՊ�U�@a�d�V
�`���S�p�L��6xB`�G��|(&�6��Ό~�Z�)̧aE=eGk�]0=��q���O��1Z��8xH��"�g���?�����y�k��K�Ջ��5L�w�q[-�#��t}�;���J x5�����Yȍ��~^=�iT��w�=fn�&�j���8;SC��
�>������BB��������l�8�JR�u�>;�C{'�;Ew��D`�	n �jS\Vz�\خ�خ����г��B�I���5/{����3����o�#O��3Ӊ$��iu��8�=���z��3T�I��-{���U�5���CKs�~Vy9�d2}�8ChK� Fg_����s�O�Li�9���CȺ����pF��5&[_0��!�����澃��a	���3^=!1NjX[f�v@�X�Y�eņ��G�Y{u�?��o����?�TIQ��B��{�u��Ƃ��<E�D����2y�&<Bí>�S�"e�v{�����d�Y�'��)��jàt��h£n]�#]���`��'�,륾��r�A���;�\G���Y�N���F�)Ə,��2Nm�D��\���)RB"Ǭ�=$H���N���$� a�1AU��6��'9=x"Q|�`~&�WL9���
�UL��=SL�0�j���ث����V��?=��M�wqTw�������P�\T���8��\��	.c8P�Z�ByIf�5a�o������p4ǜ�qa��;aH&�t����>>)ܳ���]F������G&M��&�s��tL�����=7��+�'�U�gjm�MIť3��W7�d�m[j��g����'ŖB�9>ihP�s�u�%��r΅�ӏYzB�j���S�h���-�P���r[�T[��$�E��oe�s�z���l7�xPf��+y�G�Ͱ�,�>� 7/4!o-Mo�U�>���d!�%h1k-�>ox�����uǃ�0oyI?�9�43ԑ��>Od��.Zt%*R[��]�4kO63��s��D�d���S[`P��W]o��-�\�v
N+��]�\f�Tp��W�=vjf�n�{���J���怨�{�3U#R�^�����>��;K�����%]�Q���+�p���sVS��'Әq��s�ڋB��8wg|C��M�K8P���"� |�}�"m��fB�}��[	4{��A�B�J��[�R&K|���3���K)v�`%���.݇����]%�i�'�.��,�m�N�mA<8�d(�9���DH�`ɦ���hr]� MJ���H�Jf/���7��^[g��mk�Ѝl��Je�x#�6�M�#�X�ȷx ��~r�rC1��T���*���Os��N�m���U�!�
C(�_3��m�Km?��I{�ꗅɪ0	kva��|]>-���� c,��^��d�dM���s�XDS�=����{�FX]ZZ9�u�N鈖
c7���DQ��?���N�[ԓ�-	����|�	z
}⇤>����n:ijb�FwĖA���@��1u��Oc��@|��3�)3Ez�(����������Rmk������/_��Hȃ�-�F�4#tK��sFDߠ��-��N� |���-&�\�����[_�p1���;b��^�]��m�&�A�X�}��9C���Z]�M��r�l�@�Q��=}��a�*���f������Ѱ|ߣ�Αȫ�HZw�^��Q�6SV7I���#|ypN�uEnc?(w��r��;��Um|��(o��^ɒ��Wv"v0+��@\D�����6��%r������s�Q���и����i������k�a=��&{�d]�TE��,�T�� �y '����a(�� dY�Y�ό��Z��m_���y%j��?y~�ufL~��6���F�b�B�����P�s��p!|�<������n��g�nZrs��!.�}�،������+z�dG�6�be�nC����ǷY�B`�@��$#�;n$C��=�$r�d8ٴt� �[	��ر���/�����ջ��2���������/2�{���r��bA U����s �S��?�N�H���(2�d��~K����#��m�0������t���ͯ1F�S,5�la����"�
J��	�7>�:teF���Ln���n:H���������x�p}Q��򚼥���7@���G�����8�7��լ������O-AΎ��]Gv��#�,r�栈�t�L���8�$G퇨���oYr=�f��C�,�<�׀.�i��-�sS��Dw;����Ӱ0fJJ�i�1�����0ā/�}5b|�Dn���0v���Y������]�������#�7�/#)%�������
�.ԃ�H[�9�� hn�YV��Z�T��,J���#EGr��X���{��ƁJR��O�Վ6Ι�����������3������u�;��d�ۉ��e��Y�{/����*uP�pn���3,�b=�@ՂRz��-T��h*:�%���NI�qJ/��%�A5��_E]�k�.�	�w�9�ŴKN�>��mD�wS���Oc��5�ԦˈE߲�ڣ�S	�������KRW��� �}{�*ಲ�)��Z^�M�c��Ǐ28
��>a����V�#Ձۦ��U����Ϯ����o�Q�8hE8Ȇ�$�<[��9˲�@�1m��KZF֠�C՟x�nH�y�Ӭf2����\5��G
bf���7���y��mou�!O�0f0-�C����P��@��k�ȡ����R��k�Fh�aT��j݆T?b�t����:B	;|e��-¨5RR� ~1_�����=Z�<t ���,=f�?��S	⏾(��}�bXCv�ޤ���u�x8BA�����@*�9|��4�A�����~˲�p��a�ˊC"�G��s���'�������D�ǐ�Rt
������
�n���CGV�g�=��e!� ���{��.�Prv[o�.H��ӟ_����ɧ���(G�QlEu)q*�@'uM�1�1�>`��� ��?�ne����
�
��p�2d@����O��"(=H�8�:2���a�8\���@�M�Eۖ)a���̎d���\j�'�C��G�(S��%�ʟ���3~1�곂�S%�8��9��m�u�Z\6e��EGm`
Ah��Ux���ɰT���m��!;6��ݣ�{"���`��yz�(�~�~�R�k�Hgh$�5>0W����J[��o�}	4���@�b�0pܞѷ��\~R���ܔ��HB �R�?F�Imæu���yכ;�!��N�$�?�_��l���.����w�(�~��i���uex@oyx@�U�F���p��O]t3�A�v&�녷Olb��B�D��<�\�D��s齆j$�D���.u���3���uX)K�N����PU�0��k�)�S�5�Lʪ�F�D�u\�1�G�U���y�kta� ;�����>���(FK-`\+x�|�vw���~�������x�F_��]���&�)o�|O����c�䷧eԘHfQ5҆_C�O�D�e�J�X��&��X��8��P�����##UQSZ}D����ɀ�V���<϶�L�Ő�)>���#���3L�%Ę*�%�j; 4��	���S���Y��q^-Y37��C���f���R�nP`�F��������.���g[,�N#�2����c�}�L�Vg������I2�v�Y�m�B�C��E6M��=p/h�-9ݟ�x6����0#�L|1%Um#"�﵇߅�N�l�e��g=K�M�����Jj�]\i�4#�%*w��8��%5�or�����{�������w�î�qP�&[*��HP{�'�0�`;<a>�Lj��a)�&�������OU���q�\j|+|
_R�����M�������32�jR�2w����[Q��Z�D�#H3s?ِG�2�:����)�)���#�f��xh� IJ�Y8_�}@��\��A}���������d�:=�sӮ*Fݞ�����&��Y޲����cz�����xs�Kޥ�K@�Pn�B�&�MW�.̲jZ�A���g�N`��U��x^��GS�q�ø�m��'{�)%M�\�<�Ԋ�/�=K��B���~>2���7	p_����%n������iV��\#&^���Kz�n�c�-�؝y�����F�{4Cz��*���\���	�@�i4�NсW�[��"�c�ZI�0���j�L��B�N�lM�~�K�8nl�(�(���,A�JY�r��3O���Gc�8���eSj�+�h;��q�*�Ї Z�O����m���U�j�}�j˝"�S���7�?,Sא�g�F�ߗ���u����ş"�!���4K�x%��un���J5'�.�A�&$/Ɋ��Bf��mjC�m��#��z��ˍE�5����_o�>#WmXǚ'��Nt�<Իo㥹0�^T�j�)-���jð��~�Jl�1��	���N�}R��߱�HL�D��<��$�c4�2��Hy���l��z[�h�����4�E'6��C��6���j#9�h���C�V��������%ʑ�:�-ѻ`.T��N����1�;WN���Bʽ�J�(5�*2�����k8��Z�r����X*kS�9a�"��z��l%5�s�̓���o�Vת��p�
����lBeN#'ś�U�/3W�5�A.u|r�OGո�Y�A����6l�f�!����1@ot~V�b�Ho�Ɉ�(-��k�L���-ݿg�3��\�օ	
5���Am���l��L����=0���r�%�V�֑��Z�I�L�d��d�BbO	��!6����`|��p)���~y&�v`ڜƕ��qvQ�a�D;3�5ȗ�-3���` N�3����u�\k�h��j��LG`��nz'Û9�L=3@x��s������Y���7v5�������(�+��N�� �_�g2*h��� @"\�g���ލѾ:}v�d������Yzjt�|�Ұ&���D_N��$su-[�V���f�td-`A��t�N]:�t�?7S�RC�j%��<ԭq�L<���˰u0@�[x��QQ)mM1�U١c���ml��C�>��u���p��~oda<?�T��O�?0�6��g�K� Og%��@{@�PN�k��! �x��XQ��gP�j����7�-�-�<*�9>$Vlp�8e��L5*
�"�`ϡ
�}�-�O�U#e@����U%��bZ`嬗)Nc�mL�b��H�BR��A��0�p=B�c��r��E�����/��"O0��1r�1������˹a�����}tĝ
H���'`���I��E�=�)�iL����P�4h#W{���xDMH,rT-�ĜgW/��b�F�w�?���6�8����k׽��Ms}��ĸ
��y��X�����y:���h��(|V#8��^�)2����{N�r|b�<��כ4]�
�Ѫ�C��4�X�m��d�{��� ����+�TxBX���W�:t���Q�ʬ\bpӥ���X���Ж�R$��/��%�X!��J�Z�:C	���RIΌ���]aL� ����0�YQ���L�Լ�����E��Zi\ �dC[�$��sө�:��P�	�;u�G�GÎ�
ۆ|sbt{L���jȦ�Ŝ1�l:�_��a-.�7o��+	����չ�i��4��\�h���3�Y(�S�v����:%OxY�gz?����e*���W���M�לCu��ۀ���j�=�fN�%��%㝎hq�TU���²Z.%J�
���'krIYۯ����&y6��fV����^���-اc�Z{1Tw!��4�Ήظ_��I/ \���Z��Z��l�JXV}�G�~������Ό�����q����Q�8�r-��-�����=
�GG;\?�-.*�=^��ϟs��FkX�[�V�!�"Ӛ�Z'Ǝ�&�(U�la�n᛭��3�iiP�����[�.�N� � �hC%Z��0}�}�~J��s_�wy=_4 ~U�j!B���~L�
o�@M���a^+�|��
Waqö�K��>��vN��g�d����ﮠM��^��B���pO�Yo�~�$�0��((��,�6P�/XD�8m��"�����R�VX@k+p��p�2�~:�
��դ߅#�@8$�L���4kp��ޛ�OҖS���~3/ؼ��PM�B-=�xZD�_��
��\*T�8����r�q�%�r�9��<��ߝ�[�Rk����DLG��uU�j��-��h��>(���B�y\e��L1�Rzb|-S��m�a��e�����nk�NJ P�{��̏��1M�M7����7��(�� ���S�Ot�@�Z��e�.f�����-��x��x������=�D�΂���Y_:[4�&�RGSby=�5w���Ƣe�� �%�X�����,#|*��P=q_UB���U)a�U�$����9�C�w�w��|�B�1H��}���}��(�Mo�� �Q"kY�{U��6=�g z:J�ئdJ'��b��y��n%��wT���S�t_��k*�,(2B(;%	n�Fm�)`��9�\���"{�� @�����Fǿ�ҁ�묳��k8/��8b��p�T-ǥ;���������"�)�L�}?���@��S��M$�g��<7��X���i��"y����0�GNd_e��J��ɟ�MSW
c��	G�w��jJ���;;3K]uwX�U9Ó��eֆ�5^�7&z�4�Q�xm�+mJ56���I	�\���_�����$��ҥv� �N"�'~w>��k���V��r?3j��ai�����?U��z$+A��\����y�%�kȍ��kW�Bk~f�{4߶D�S!(�v��'�@R0������VԨ��5�zT�9٥�̎�V;V�.]���
�2��i	�EH@sN;��5w�&�K1����i�`Me�G�rM����I궭�{���}�"7���@�Hc�c����8�|���Ap�@A5p�ޕ����9ˌ�m���M���V�N��C�u�{�dK��&J��AВ��W�������9�.���iΒ��e��,��s��? ӑ�-��z(Q�ҹ�.�oH���)Κ��ͅ=��`2΅�`(\E�ԡ��|�k���J6Nx����k�=�~08����z@[�����ڞ��v���Uz�?{w�r�/���!%��՝�]���i^�p�)?�w��F�g��55�:� �r���	 ����m���J�������<se?�c+;�R�_<\��_]���1JR��#��vݑ��/��:XvyD�{D��Մ�K��m�W��LM��dLo�UA����)W��.Py�f#s;VT����U�-k�VYǵ^�A2�#n��Ss(���ҙ���~.�]Wz�x�p����	2�2�~�i����������Y
�N���-F�!+���k���Ơﺪq�����Ks�"�b�q�E��]�%~�?����'�=����S[�+��
�y��Hh%',���ߧ}�:�$��w���X��j~��_c�s����0�s��\V]�o��`~-�(���3��b�I�������$�M� ��dE�dT�F���^	�&R��|�4�Tݻy�~�pq�`脼S��}��Ya1�/R3�ӊ)�&�ފ_( ��������)�$(q�8z֠���CŨ{U)|8���]XQ�Υ$ܲ�NT�k��3�	AX�t���ie2zNY[��{O^�&\X8�^�L�"�&	A���(�Og�l�ݚ@� �l�S����k\��/h���{k���!�j���S�'8@"&�=�gpMB�|Y��QNE�Ξ�S�!5�����!_'�2�s�@FB ��х��T~�;��cL��m��?uLܢ��Hn���G�zy��4�nƴ��F>5��D�a,O�լI��R�B��~�-s$�]kM��-��`!�Y��H���qxm�j��6K���z��4�����~��D���i���<�t��4)�:�:�����T�[b���Zx~�O	CP��$����Il$?�N��ָ@�u�_2+��$�ǥ@��ko��^�t�LǄ᥽C7�xܫҟMp���^�-����j�����!��K�3�:�#1�?�	���5���	A�Oֵ�t�Hq��yX���w2� d��_�����c��i���C����)E��3ܓt4��Zp�9�kс�t8��U������ָ�YN3�XG���3�<]�۫@.!�?�?��s��p��9I �.hS����N��iC�~h
k����:�#�%�Ud}/_����7-B��n���5�{,$���^:�2o>�ך��xt<RfF���^�;��ʟ
�_3��u�"v?�-�z4C,������`��a����H���.�&,I��T����v!#Tjx��dL��I�0��^m�1o��vYJm���o�z�ҽ烠�2~�wb0���zT�և��S��8��{	٨��EB�e �w��+ֈ�	͌_�O�,��i|�����9�����kR,��&>�+M���-$ɐA,r����9.���am`w�J���jh�mS��u_�E�Yz+%�SU�F#�4�5Ϫ�*�������bGM��@�~q�ed05_�2/:Κs1+ާ-ZrN1��pҾ׬�8�Ǔ�xa7�lG�M�����o����+�"�tV��ɇst��~��墓�:�>vK��>D��1���g��В����t#������cC�1�G-s�L^ ����<B7
1T�,�u~W����ڋ4ȅ⟅T��,��=ڶ_X���C�� ���V�$IZ�B�B����ȣ~W��Mn{������;]�u��Q���˼�S����G��,C)��k2�oP��q�����趑�aQ{��ޙ(d��B������吉��F[L5K�)8/M�M�a��5>"����:��b�a�|�3�8�QJ���fXi�/��sƍG6�x�kI�T�IS����8�&���	�:���)�ɕ>�	�</�k*����M�w�=.
��|Y�xO�4��̈9qu�߸^�|������U ������5�䕋��E�zL����BΙ���ө��xh��qǌ��暈�NL�=r[��������o����\n�T^g'`��3P 6d��7��DȜ�(�@��s1�9�ɡS|ü9b��i���Q{�Z�:)y�/��o��;F��������Ru���!W>�Vm%��#�r�I����(��>M��v�����`�I᎜����UѾ~��獾���	���zGs-�u~�c����$Ͷc;X�����#����g�u���/�Q�P3��n�>d��wԄ�j��%-�*|}��vҠ�x�k����P�D-J�O�Su��wD��H�V�t��%�r���JA��[��Kh�i��w9H�YZQ�G��"���n�^�[1b"L
^i+�O�76(�Y:5zsOm���\��#Ck��	v�(WdVh�Me��ē�Ӄ���mE��G�\ ��g�
1�B2���K��P4;}��2!�՜:b��|�\����n��S�Ou�[Z���mw�������K)���<3~�N���񑹈����Xx\��5�����>m��/�mم������\�x�ph�@-v}�5���������)�H�m�j���W���m�o���w��`Gh�	�e�
{
툯g���Z:�zuTw&���6�yn����P�ݣ�5n��֢jd�l?8���I���v�V)��!�a���ɖW2wz|r��V8*�+KO!�u�@��pg匨�9��/6;/H�5 �a�-qmU�|�S�N��''4�`%i���i����x��M}
3�M0������[��#��L�u�A�e�4l��O�Ƣ��1г ��{�z�ˢ�lc���^3Ȓ�ϝ<g.��цH*��BH.���|$�2�Hov�����d��=��r^ĵ��	�:7X�PFNa~׬d�
��܇Y���'/�r~����4m�iSt��c,�d�Ʒ�w����
��<��l��<ŌzZ�f�MY���� �pJ��ބ�|��asH�{�8��2���d6[W���}Dl�6Tj�`� И��%�r�]��p��` i��;��9%4����=E�ȃ��J�ݤ�d�`̋�Ԟ�꩕�7���nu`;�q}E�1�8��\bv�P?���-���=�eY8�:��i��q��P����YL5�CjGU?r���|';�rk��M���֔i�R���F��YF�Ik�"�H0�,��8`�CT�V���u����\oe��^��[~g�ҙ�0���~=��y�H�Du
�T9`���M���7E�&����P��ÂKu��%k�{3��^�H	x����kT,_iĶ�p�;6�`%�sD<�xiV{y�Q�[Aq�0���Y�%r��@�,��<!Gq�ƽ���Ar�w� 苬��UqAͅ�$F�=��ў���*�B-���z늖e�D6܉���N]���^܌����t7��P���f�P����h�ٮ�D^%�r�Fj��2��PS����^��v](di��b�.���]#�k�ᗷ񶏕"
�*ă�:���=i*��[=!���hת�/�"�w� ng�BY��l�W���o>�2Re��Ğ�~�`f�I��zÂ��������M��Y~\|���N�(e�H:�f��2����W��MyNJ9�f�C�������zyt�
~��Pm�Ə݅�Y���i,ov�`�k8�s��9���'�uA>yQ[б�@���t���	w�R����8mѷ�7ҙ���c�1J�s�NUs'�<�
er7hH�'� �"������<����!dS_�kD�;Bߩ%�jTa7^�\۽��&E��u����"�I��9��z���]�3B��b~.@���+��)�<X��c�v^�ش���sNA"��Y����P�}��O��)1�<#^	T�V%s\Pn�?�OQ�f�T��%�U��-��x�� []�c��淭k�OLZ��o��ƃ��R2�1~��ȝ��JQ�㽦nߗ����,p�!�\�H�֗跣�m5�w|�'�Ew�zLӟ�*'��)�_(F�#��&��*/Մ7���yԫ���j�S��� f���L$	�ȱ|���b��_��J8�[�rf��!�-z��v��ąc�H����=Yo�=�@J�o;:'�d!�\-�&*鹚�HV&E�ϻ*�6���"Z�ߞ<Z��t�I��RmI�Q�=w֕H5�'�i��p��]x�E8ؒ[Ü0�`;@��]i88��Tq����P�ǯO����{���-C[̷����>L΂wY8���F���R~�!f���Iͨ����8:n��hthf��p���1��?iL�dK8�S�k�5�q(4�-]h{F��>����@F��#x0�}G�5l"������$<�aN��i*ΡJ ���V������uv���bg��/">^xZ<qX���ءr(����1�#I�k�a�!�O��oK��sFŦX1������˘J�	�!O{��QB���x^���lˉ�7�"[�"�n ���4ZW�Ҁqm��bS���P���7?g.�Y��iM=�j'�軘%Y��F*�q��Y~�p�9<��/�M�vy�pm��>��}�è���m!��/(�q#Q��]�7�tB�0�/\z�b�_���Kbk܅B�vs�n۳�5��c|�h���C)W����0��2?�q�V<P5���0�؀���M�/���I}H�u
��f|Zs���ˣr>�?���!�(�ye�K��q��t��g"	�mb���^�e޵ jηɂl#�}
���:og���	5����#��X����g�N�0�c���1c�<Y�Vi�V�T���,i̟��xo������uW�\qB���.C��3�x�'$V:���$>��c�rv�T-�3ٕ�Uw�%��fǌ�;����"!��F�'����pye�ҳ�{����P&�M�|i����S;�W�3х�5|�ظX^����ΨaM�� ��_�S�k0����5"xg<��:T����G�9�߀��># ͙���Z�Xڿ�T��H�C�A��mm֖�]��׊�ɷc�����bo�q����yވ�y�{R�w��Aj��l�M^)~���{KN81b�)�T=��V�2�K;B�o�&���&�xh���)�$|�����LOoד}��I�b޳���}o�;�<��cC+�!;��!������0x�g��N�'7M���n��EpGU��q������G^�W˧�j!��2`3Q���I�� ��K�kW�<�KD�Fsdo��1��DŪ���א�HͲ�\;a���� w�(�a���4f�fZȊ�/�&�E[�aQ!�xVY��Q)��TV� gw�z2��������k6�aN��.E?7����]w�����y�GՂ�@,+�+X9��5h/L1�o������@���M��Y��_,��a͈�l�]l^���}�Ϳ�O�l7��ٴg
]���<\!���ޕ��B����x�\8m���158�i�N�#�zÛ�,��S����ک�x�"��}Ğϸi�@[��N��	��|����JD��ܗN^g��m1߃6������@���y�����b/;4�:F��:`�CA��16��v̃Ojj��ฎUˋ�Q0C��w�ӊ���W$�#�|�ϻ�DU�,(�P�b�M[�W�^���B���^��ڷɞ�t�z��P�����(���:2Q2�n��ov����qЌ��N�*�k��]�F5מ���z���$�7�OaU9�y�ٱpK�,gHVm*U�ͱ`��{�Q%��/�����5SzJ��&V4�v�=��r/\�4��f+���d MOQS��.;nL^bE,�X,&1\`�����(,(nW��y.��+:���9֛�ƪ������CSBT��V�)��S+N* g��,�ʪ���|ğ+����1���R%3�ъ�0"s%��6��.�F�U�|]s!�F�V�R�W�Ĥ]QD=RF#�q�:�����y��#����x1ɦ�D���B����v[S!6p�82Ci�Y���� ��q~^��\w��X�Y�9��!a��}�-��D��Q�/��E�r��^q�P1������RUt ]��r �����:kFd*!']Ł��ߨթa�g�Cς���ۥ��O{R�KZQ
����g�>��Od
_pEtī�D-����j2�������.v���O~l�!ޤ�H5�s��f��o�ORЏ�y2[��.��)��La�a�e��V��k�����8�d�Ƙ/K-E����%4$߿E����%���p��ĥI������������ד��#c��sޖ�qMsD"$��D��P���R���m���$�FE�+�gƫf�s��<0fIP��O"FL��+�R�y*������n���p�o��C⩥�S4<XkXn���)�����|6�i��@"}LO���� ��8��B�����hf=6�i�B�V���Ep]*���&4<�Gaf�>�ϊ۷_hA�s9���Gw˃�R��l?A�-c�9�4!�
g�C�A�u@�W0�t]uH2�l�����x���!zx�;Y4,
��ՀG���"9xv�*H��y�]�������#O�����*����+}��̇7�3�n
�K�`���~4��ṿ�H��Y�S~���Ρ�a��`G��(��D�`��1���Ow��Ox| �$�O�[J�����2ʍ���ѺW�gHh��~LE�����E4N�k<�>����t(!j�}�D��|���]�"�N4K���I�q���˽ʪ�1�Y&��.�p��o}�ZΟ:�wS����B�F��#�v~���,x*(GG΂�Q)�"���@�ԦF��Y\?3��<J�� Gl�3��$��z[,�/��P�F�B�r!Ѭ�	ر��Q�����lĝ�Y|;���`���˂�i`�Rh�/4�Qk�K)�-~g��0�9}LY�4X�p����q�l���e�ԣd�V)�,��n�2��w�Cʼ!ƣ(
ݓ�s<S
��j��Y@��^�I��9����U0�_�
]W ��"�S�b���j�B�j����T���/�R�a�[�v�Θ��V��8~��߮� �Z�-a��g����u������Z���L�;�P{N���k�MV�b�}��X���P$)9n�N-��,�P�m�#q������{U�I���s��{�F�&� �i׷�G>>��P9
&SJ�>�W�F�H�p_�����mK�5��!�H*�y�O3ܣ�6ԃ��&��BÄ�E4�ޝ9���$xY[*�����l��N�;�k�� ��iae�Y��#�=l���r7�b�7�#5��r�\�3�k gF\�`hV=m��*�k����5"
:�R����͂��vܠ5��j����R�t����ڄ�п��&m
���^ս<1̖B������9*�w#Z)��X� ����lm<�9��+�zK���9K��U�(\�Y0�`{�འ��s奄ڑ��C��R��&�/5h��� Zf���)$$�y=����0�5d��W�U�ҏ���7`�MJƟ��+��w��~���W��2�wP6��J��$�����v\J���E�C]��,��r��n��@�TT�	��}E��̑���9�y0�/��GNe�~���@G��D�?'��*��Iqv���5���t�z ����(5�o
M7�>dt|��p���b�$��7w�.� f�#6E��I������|���x_�6
�}*`�E�[����$�e׫Ū=�w6ɨ������>^
���j�fI���Y��s��@�e�d��O\k�Qr�n���Ȗs���K�ꫀ5Է5�ɹ�D���d����7�Z�;�u%PT�v�C����JOX\�̧V�Z>׋��(�4��O{�i|����Sh�T(����]&��>^^˳�c�\�9�et�@E��U hE��R���Fݔԧ����1�m��u������4<k3����zAqkv�@�幋3�Qp�]�W[^��{M}��O��±̦���dV�ש����%�9wʸY�P��
�}��7����P>j�(K,��ɂ>����˽�A�7+�Nx!:��HÖ�������
)@����V�lg�Z�YUx���)��D3���{��೅`�����Rۗ���hX�V�6����A��K�@�d�g���GP%��u1Iw�� ��x'���=$�l���l�%�C����$�,U?�||ᾼ��l#y؄��)����p@!F"҈�4���!��'/��fە+�Է
���>#���Iw�{�DutA��e�]O�!��W�U$�N���/��tY�Bo�6ܭ�v�)Ի @���j�f�Y�oo�V��ʍ��
������IH��7ک)>�
qS��4�7X��~���T�][|FWA�Ҋn�Ej(��=K�;�x���A�]���)L&=E>��X����ڂ ^�H{T�,��0���!���Y?}��x��v�B�+H�9Mc��jO`((�n'm1�d�Mm�(�Em����=��a��[��B|[H��aO?	X���ߤwu���K[�RS�rW{�w=3�^EfT��n�	����Q~��X�JIO�a��k}�ZP�v|��|*�|�����(��C �{oC��?o�4��\�G�ZB���C`� og��U�Т�|X\������tf7_���A����GD��a!g�MS�TL?0c��)Y�aJV�<�Fzu����'X���y;_��f\f�T���[���)������M�h	�Vֽ7˩���j���\,�D�a�X�Ժ��Xd$��4�2���Q��DN9H�$��<+��j����h��{P�/�RF@�t;O�W���X�A覣�-�|�z�7,w3��Bte\�*�ͽ[
�s��Wh~���'5
tbJs�en��1��PH��UY_���\����nu6v�G�˻�W���O������vh�a���4��r�[�<XX5|U6���U���D�Y���u�h��&�|� A�E�Ee�<��}w���U���K�$�p�ZHL�B���O�����/�:c�=�`��d�2�)o�M�`�]���!a��
d��9)�x�=V$�M\[#�[G�Cu���T�o�����A��x
 �x��*W�[�� 5�+���-G��n:5�W�A;��*���q^�V,l+z�2���)��@!��5�p�Ō��C�Bz ?�gR��z���k��t�-,��Hd�/��mm#=�c|��I����U �������'N��Ht�*G�dp��oa͟:�^�Գ��VT#ZY,��J5J8�֬�ZS�{��HN��c���e��u�Rm��s��:���j�����rJ '|�t�=�,=�b��7���ř��׭v:Ch� �c���jFS��qNө�q����@=�3!a�6qr���Ix�갗h[��\F��|�mbP��?M����Z��Y�F�K'Lg�a�h���H�ЭO���N(�|�cQ�p�/� �'��ml���@[U����l�V�o��yP=��g
zH4�cE����m�&��2bߔ�xi拺��v�^"�G����&q/���� 
Z�{~.�oK����X�tRHr*�V��O�J:��Q}1@��(�@3D{��#�/\������W���5Z�I�8au��e�X�N�چ�:� ��K�3F�����w�vԌ<%[�Q��������}�# ��:3���,����v�����<yH:�k��k�'�<k��^(^ �+ɗ���i��*�wĐ+�9��+��@�)1$L4}�&a��T5Zo��u�ƘE?��<�m��%�H�,�<z2Zc���H{�V�dՉ��n�-�nQ���2�*a����iEڀG(�S�a�al�7�<_��.�<͉^�g��&��	��A�v0::b�L(p/��H�� :lk s�s��kg��S�}X�����Z&�@עߦC�J{�%:襆��l��w�HDL?� �����Ɣ�)=)�s�K㮊�Aw�-��8�f.�[�l%��WPG���]c�������a_4�i��-��΂��.���v_:q��?l��ۑoI	��D��h_��c�Zc��ǢAu���{�^Bw�N��N�i\������V<A��*���6�e����Q�g��ihM����4�'��H��UW�3��䙛�}�.�>r��D�%���bSʉ>��
����8���'��t��2�ޙ�}@аҦ`	W�ssv�ª�䪽{M9�[��"r�ت�lmO���9�;cL��|�|�yk�J�Z�*���[�����~�=iO����(�Q�y����s
����ل�i�n:�U���S��]�҅� �`py�})�Q����/�O�w�2�����A����4ׄ�B��5J[.���l�$u�[ܟj"�g|��t��F-�ȳN��^�G��ȿe< (��|�$Y["e瓡&����N�x����7-#[�� ����O�F�,R/�P"Q6�?�����~�_�#{o0��8-v;)�TY�dG��+��YS�����#�(�����Y��O�C%�I�ܕߏ��GE"��݄`U�~b��]�Ǩ��H!�0^�U�� 9��-��>��n����]��0�w�����ТC�������]�V Kܴ"|���f�8���m�d�Q�{�LL�]v��G��$e*�����ZM�hx��u�����=��������Ò� G�p[njw��w�#�>�W����F���*U��������]�Q}�L�>�h2̋w_y��w?�@75s�c����_"߀�?�8S��1��{�_��Fkr�E��������"9�����v���5�U����]mߡ�,�n�R����~
ɾPG6R���)+�@��	���6��bAPA4(��)�T啅��rp�{]�%)�VDc��!�%�5��"OHG[���n+�MD�� �֫���8�/����	�g4{H��W���l���J\t'�7��U{R�֩/%M���A�B:�E��[Z��$0f4d�:&���t�n�Ų����eÇX�(�N�}#'�<��lr�c��h�ﲠ�z!m�K��-W}��?�`�ǌ���!P�H��I1X}e�z�9^��8=�%&��l�2���J�of�U�&o1b���O��]ۜSX�"�T�����:�ªgIj��H�?�6�������=i�dY������F2]�h��v������̸ՅP$�M��ɒ�-�c�������4���DQ��,ڇ��U+a6�7M�}9{Lpb��}��fxn!��1�ؼ:Wd%Z����g�q��8j���:���?żd�����C�4�	d@��$wzS�~�s-�N�Y��	�ɚN� �*�Ռ2l�b�w���״�

Y@���,��#b"\���>l��/��ce1�)ɶp++/����-��KD5�d~��L\��:�2��uF��\2�׺��li(5�*��Չ��!��/"\J�3�E�1���C�AMY��b��zxu�;PQJ�./-����1���Y �����D $�{��O%���6>w��$�ђ�hG3m����Ag}�ގ��l��RX�2��p[����P$|{���Δ5��P�:�U��LNt�Q�^o1�r�s5�9}ŧ�Uex{`q H�z��MgA��� !�E��R��ф���)�X�$��ҍ����C�j�PEU�T2;�Iq�!��^i���Y/�h$�5(2d������'��]\\݂t���ksn�P���D���v4>�f�����Ȏw�J�> �y(T� OE��fNq@lл����[�����&�78���h����6Jlخ�:Y6�z��F���hc�����#b�_2�(]/p�����9<����yS��޳���З�X��L���R=_^��ݟ�f�����m�����>*�ŨB�K��\KSq�g&�.;@�	�Z��P��Ԙ�=	������>5<1���iQ�!g��Y6<>����*��a�w�N�����1�C��V��c�r�S���ȅ;G��S�EZ*{LX�a���x��1fd�\6L����v�#A*�k�G���/�v�}ˁ�h�g�{A�c�{5깡�4��/��a����y��uf�F$ȷ:�u������<�^�9 ��`�G��u��tC2zb)���~1Y?ۤ���˛���̥��a~ɶ8B�	g&��O}1�.�����D�r�{ݦ�N�JNw�4��\��2�G,aQA����0���}���2���'�H����N��\x�#�&qL���n�z��H$Q�������nG���	�����*bxjC˦-��-B�"d�L�4X#�8�[�}+��k�V}(��
A��F��>�n����A�|�ah��E%^]��ė ξX�^�ğ[����$��Pz���l�P����̡�zq-���y?�<�j��i�;�`��l��{�xY%��9��"&�m��١0����C"L��賿{x�eKon��M�TM�ퟲ�I�n81B[���#��\�4�OTf��J�S�I}���yQ&f��],���`���e��s�e-_�遜�Vf�[^S^yY�F<R�X�i����ue<� �.�R!��ELr[�/�(r�ϮuLA)��S��5Jn ��a��x=h������N�,`�<��? &�Y^_�͊}��!�#x�B���§������Q����j񇧃��+M� ����
c����@ga#�=�}��	�����.lU;�.�����r!��,�V�6��󟀽�덠�8�j������y�I	,��"T�r�R�'�@���_:x>,� h��.�Q�ى���~f9�TI�U����k�4A��;D�
��%�D���S��1e���<k�ڤr�9càK�$�΁Ѱ]��_�j��t$�V�o0c�&��������	���Z#R�����T �$n��zX@��	����=�!$�V�����N9(��R���kQY+�5��5��v�ݬ��j%g�BNS:k�[�8+1.*XrT�g%΀p��d���-�7�:x|���&��&?�r�N&}~��|��Ӊ��QP`7��;�x:��m��gJ��~Q��]L���e�Z��"ܰScrE&B�����ô��θ�q��F��co��e�L�e*�ҏ�\HdԱC� ���a�e�[hKZܨ|N�'ojU���2!�Z��#�5���NE]�k5���,4�M%1���Z4�
���7(��2h�9{.�cC'y���f[��Xp�����N���
��2�\�n�=��I��7f>��w�P!0)Ӏ�n�1�tb��Ͱ��5�ƞn�V�|z[�K���T�I2g��dʗ�Q���K�w�J�TC�p�k����T�H�\��_aV�e���YO"Q�X��xS�hR*
V�v�n�}�<;ZT{Q�H?/��n�Eu�'\����3O���Sp�C�L7�u��ø,�V���v����;��#9��tFC��u�ڰb�LCI�Ҁbݰ=�[){|�\c�
W�H�%�/. !���Q�-	���� �vZ����J�Sx�/��9������p&e���TmE��}G��t̎]�0�ȷ���D3²���|���O��[��*��^t�"A|���M�ek���I�K�<��w)��sp������ӝ]�u"8� �3�I�	C�TKs�D<L�+"AI;ݕ��y�9p�A/�)�pL���"$��R xH�
�_�k���R�_�ϊM�]A�y���T�t�V&M�L�L�=2Z�))�K�kX�M�j]��p���	�D�?�uw^
��}��<��ʞ���Q�}�'�*Ϩf�/H�r�|Z���t�N�ph5���C�G3 ]�a�H�
 D�{�.ݧ� 1�Պ��X����t���b5�y3�A�^�	�:�"�m�������Yt�����ǂ-*�)T�4w1�׫����Lp��k}���E�a2�3�
�:������@0u:q�L�T[�$/����x��~J�Q�����&��G�bl�n�K1fޮ
��i�����5AH ���Da:Q�c�nq7�	��J7^:4��eY��d�Z�E�rj辮��ԉ�[�#V���x�3����6�`b�;$!�才E��G�p��D�*�����R�M��Kߜ�)��
��m��5�v��H֟,�=Ք��@�s`�au�kO��*p<��6~���R�@��K&>a�V�A����� �q�f!)�ͪ\ݫ���C'��X��5[�.�.�@>l�A�>�>�����c�"���TW#��C�7�� �]�t����QO.���R`ڮ��iY'c@���0:S��~�דڗH�ڎ��t/���"��=7,]E8�NQ;� �Rk���bDOv''BT���ۺᏭ_�68�ŵ9�ә%=A�5�ŝ�T(5M���F�'E4�1A�(hZ�l�<2�X�W��*�1� F���]�I"D^N|���*��7��(����!���Й�n�F�qDS�p4�d~�C�T�A�/T�P�,�n�KQ��v����ݥw�H��m�-2_���t�<��p�=���p#�d�mZ�<O9@x��5���4����ݳ/UƳ5.��7�<�<B�{Nd���M�����.�-��L	5(�~t�v���S�=r������8�7\d���:�9i9*��cؘ7���;��r%
�K���P�}���#;cʐ�jX�g~$Ŏ��ŉjdek�r���q6SN��Y�hd�*�f�)N�\sL��nϳ��E5��|*h
�s���T$X;�WU�|��Ț=���z�v��y^��U��"D����,���r���ި�w޻����}U���������ĉ�O�5t���?��z��e�\;��w�#E:�Z�ʥ$/��eh1 O�����9�����K���J�� U�&�-)�lJ�=�kAj?z��F!aȱ�aA�R�o.�(q���ǅ��<n�����Ǔ}��-�ri��gw����h���.`�\	v��W:Z��kb���1g4�A��-���u�<�w��lq�e7e�kV4��H��^����"P�M�>�%&�w��/�%�s
&��P�\;���}�h��N~ߍŭ6�ݴ+�$�&��$����؀���+趧�Q���?
��bc�P����V��L�s�LUJ��{yu�}�Ex�)SK�@�ڲ�㛼��������P�=��s\��$}k�ҁ���0���s<\�V�b57=���$�-b��5�n,�"*J��N��V�+Je��F�BY=w��7����r�D�T�vlF���BR��X��Q�V����4�}�S)UL��o<� 0��;�K���<ـ1_��^��d�-�칚@����F�"��Q�۝K]��p7���^V��A��4C�41n5b�pX�;ó�NP|[�(�#�V*+W��\:xDI���)|�|d��pQ�R<��yQ��P��IXf���:�� �vg"����9�f�l�s�I���ZP.5�� 3s��"�W�QVM<^��%��W ��^O�#�8=�C�RD����ջ;�~�7M����?Tqz&�w#D�ӧ�ݺ��Z߄`W�H=�V�i��2܍Y�g77}ϸy)gk�B[e�8U�^�Leg�@'"G&'I����������%�-m���)�U�W������W�����؃a0i+��=Iu��B�x��`�K��A��A}���g2m�A����Ny�xw��E��x�2g��~���Ü^�׉�$����I�OF$�_TeW��E�.�ł��
:c��O|$^���U/|[���=&.V���2���rZ�P�,ݵf۪���c�raƣ�gd(�#�_��D�$�"=�g��n��aVKM*�GzD�0}>�}�_���lI��P��/I����B�2�?��\�l_��H�����$#�j��0cfƗr�Ν�K��lxVY������O,�<[��-@(��W-��sCc;Rj��|k���j�9Lȏ����,�#���c�I'�n��m!�l6:80Id���(Q��E�ɏ�f�[Qv�{�C���KsbZC�E��4��c�;��[I�����V���,��"*LM�&�JK�����r�ԇe�:UJ ]�*��*ay`�����A���~sMY/u��t�A��܆�s�C乁����K]6L�mS r�i�n\�?)- 7}���﯌(į3L�&$�L9W�ȹ�Vn* :S���2��o��ق� Jh[1J�£��@�|��H	:g��]�צ	7x^�c��~a�g�Im²;U�����~���5D=/��IL���#6^�z���M�ns:�D�Q���|*+N�1�|[������1LR7� W��NK��t�n�=p2�%В���V�d[�0rp��ś>I�)9y�<OE��R��xWgA.1�,ز�d��ݔ������.Q�����G��eBVa��|����bVw2n�Ϙ�ֿ�=v������Rm�#k��X�6����͜x)���=%��vث�
K�bA�I���M�k�KO+��P�ſ����	�s�aF(�S5�\1��RH~&Uԉ�Y�B��
Ԝ������>���[���u7ڠ1%����ԲO`��Zn��*�I|�W�Ҏ��f� 
�����,|��p1�g8	uB�"��_I���1a�
�i#��m6&,D o�L��k�qn�ѷ��n���rz�=}m�}W�>&v�ǰ���a��6A�H��'�I/�
+�R�-�x#ӵ��L�a�i:D߃6Jt���!�u������S�]�͵��#��@��Ԧ�}��鱉����Qf�A�`��g�Y�����I� �8�/<�[�O�;���b��9E��+�ׄ'�Ye�n�|7A��2�**R���Q��[�d�`�B}I!N
��=�$H�w~ظiL-��ȕ���l��Hl�hu�c-���n!��� P�sC�&��&me�X�{]x�^�~��ϱ�sS?����WD�z5	��@F���ٴ�#�H0΢g�b��R_��u���P?��r0W������=�SW+�q Z�]W��/�)��mGښ��e�<��{�
I@��j�ٿ�����2�G�,@��,y��+�8��5�!l�G_�7���_���B�N  �Lr#��m���3�}3*U�P��2��m&`�<L��@�6M��YO�h½�2>�Ϛ%����2�(L5@p�O,��N��rF�k�)���c�3:���4{�r#JP.*.ή.�4"�1I��5����e���V^��)����n��SF��=E��J���.$�7�'�T�u�xЍ'�ք<�ńpp"'�}��]�V�D��"��Cچ������}�)(9����J�M�
��Oos:��T	9�;�gm�>�F�\���Iy
6�����S�}�����u�x��(�0s�����B�� $w��+�]����/�\OP�d�]k����GD*�[�~V~:� 2���k$�l�{�yvR���E�\W%���������vf�<�FH�s��&��-B_���J
D
@;�nL�rxdU��C�W��!}>)_��zկ�)�����G����6��1�[�`��Ƚ��� �F��,�e���2����I}6�%�\l�A#����f^�"?��W�o�"��d	z����l&�,��L�N�\�1b`97,�栍P$���d쮃����eZƗi��f�0��,`ۊ�%���ա�I�a<�Ҹ"Ŷ:��R��	�DrP�4�*�Y����a���{���d@{]�Ϻ�{B�x�Dq��[mߒ�K�/�`�1�������d��ߨ����l�?k8˘y6JIс^N�]r!��j���𓐭�W��ɋ�Z�U{�o@|��+['[�U�vZ��a.�4�Q�篶�M$c����O6���%IA��p(���K���9}�C�Y���G9+ݡ�,�v�4h��������P߽v-���:���/��o�E�pȂ�m���s>o�y6�N�ݞ�!����w��j��0@#�/C���6��ԑ2t����~z���ô��;8��s��4���<-�j���XA���ۉ �l�tu������[tҤ���r��ݏ���ޭ�����#�w-���f�X�v�Q�鿉�,�t�$�Y�t��4�	�'��\`>����&���S��0Q$�!�#3�Z�B(l��6��E��]�����3�ĉ4�0�a��Λ�͎�mb'�0�����[K��D��"�ň�HpPwG�������)ZRKT᱁�ѧ������\a���I�A���n
-ͯ�<1�V��6C1�4�*��m�R�� ���oZ�d��th��
#���E�&!5<Jwi������Q�!��a��{^�ˎ�},��'��VW��������NK��moT�c�����Q��W��0$`�xz�߫ܺl�z5
�(����_Y(�hB����O`��j4��6G5|K�Z��bԘ!V���	��x�m^���`�n��Q����	��i�
0��CƛD,��(���za�u3b����L{�%)��$�k��ob��F��dlOA)�%R�Idg�^2ݪ'Z8E�*��gx�DJ��1gp��s$V,�f�����0�(Q���gE׿:�SN�SE6�Ñ(����CQ��-��9U��݂s9��^,���Μ�Y6i1�`�-b�R�P˧@�!g��LE���T�ujBSG��'/6�%�֝�vw��O*�}��#l�˔��esx�a#�&����������܀�=�5�N��F��0+ބ*������k�J��Y&�/Y?Y˦L�G��X���;2Q��زpQk��؏�4B%���3uq��5�2���Z�d9�N6��{O{��M�-�� �\fB�r�lAu)A��T@��3��?�0��Y��h���Ň%��U�S �	�!ѽ�x��w�і�N��H�}��w��	��Ŋv����z��ZQT�����(T���2�	�:�8�@�u� �J������r��?��s��#nP�e��zqn�}�ؼ�='��!�T��h�(/�޹��Y��!�욥#[&6UȺ�
ә�!n����
��έN��-���Ө�dh�x�yDbQT���@�?���Mv��e+P��$����〳g%��)��M:\������S٨�[��O�8�1@F�,�mcx
��IH��}���J��x)�?Mꁢ5AI#�[�8�}߀oV,�ZW:�9_m�u�K��Hj��Ǖ����x�0͔Y�@�=١�@rXc��%$˦Ww�&��<�����U3H��T��:��]d(��2�G��Wη��`B_�4P��E*u5�v���w�+�gr'��qkW$s��+��Af. {6��\�:� c��|p��飃ږ�'b�#bw+�����TA�p���"牺�w���M=[m;@�JM�	�����q-Z�r%t�G���7S@�E�.��ս3,x�ׄ(�xP�V�x�����$Č�ǅ.oW:���Ś5�O��;�@��l9�\8?`gh������-Me3�FQ[m\�C���s�`���z&���u�"�p���l����~�N�/K�l��鱎��!�#��TO3 ������ �]*�G���{PY_������x1s��{uf��e0W��w��4�uE�6:�e����R�E�އ>n���Q+�K%�V��JOݽWʵ�^v�[ғ޸���G>:������i0°�#�p���&�����&�_�_`bcf����嶐NCJ3�G���r1�~�I8���'��ܶI�4-A4C��Kfn��lbt��7��U�%��hkK���x��gU�M�R�7!�������7��ie5��}�#q��qi��4�L�K^G�]�m8�-ͦ��'喋�V�R��	3Z�8ԙ���&�}m�4�P,*��v����N�b^��d٦:���k(�����ᗺ���8�(���٩.*fB�j�y:=��s��a��u�D�Ő?��Gf�^�f19a\'uMG*���1#=��zC����#��6�=8���ע�1D�cr[9E���1M|JU�,AnnSr�!1|�L�	yo)H�V#ϰ��+���k��\>��)K�-����{�	.�<K�z��0]����w���;3<��]SH�$O�Zn��F@ɞi׋ gR���x��F�.GM4�ٽF���ܴ��cY3'����m郐��v�:�q���U�ve�9�TQCu�~���"S�n:_��LL�K������j�&���t#ׯIvQ�	��O��\;����2!Sq~�Q���s�5�U�ؔM�'���T�É���/0U�Ҹ\}�._����Dc��l?q��я��#��?�3l�?��s��n�,v�Khu9Z��d%,�!R4�La�*hlୁ�ï*J���Hw��[Q]��]+�-A�|���A���a��.Q��u�	0��	��	��f��'������Q�\���	��7:ص�������=�z
����`!�Gsn�b��ر�ţ5��+���4�^,�
�Ĕ^B�]n�1�p�����9g7��)�	�x.�_��[D��dx
7|k3�To߼��t�1>��#~�g��*(K)��ģ�=XNƆ�:Kd��l蓴{�!yQ�C��+'�S�/k�Ƨh6��=�Y~�q2��;��~�?�g��θ�k�yR7`���*Ј�z���I1�M8���Ӻf�C,#[Pt������C�_�A������<w�!.Xl|�n� Ί�{^@�g�f4,C�4�CH` �oVk�z`_��[Y�iٗ6&i'j$|�NO��aڥ#�J��v��4}+�]{Z�m�S��ΪZR�o$�a xk�a
�+�V����؛���ۚ�M�^�Gf�S�J�<ƭ�����3� �'������nƞ1]a�ɖo�8�rת�h�bV�W�ʺ�<��+[-�LN�i���\�Ȁ�&Y��iP���ؓ��ٓ�D�
SQ
8f�!�P	�m�,�z��rS.5�sU$?�jn�:�#��e	�&�G��y��.�� �>l����IW���]� �pR�<�?�Y�?N�U �	�	ay%�/�Ņ���	S��m~�G�M��"�="E?	n�^���k��-�����x�3��v��~�k�to)NK�t�I ��|f3h� �J�b[��U�:~�Δqc���a%K*�����+�]�+�rh�����E_�xO��gV�~W�Q��5������)?��[~��d�u%;bȔ��ȕ��a<�Y���i\�M���FƮWr���ĕG
����}�����{��?4���+�?�� SO�F�x]#�횔n�[�I����]�{�׼+�;Vf����{�f�S�d
�e�@0Kx'�����5b��Ɉ�A����a�V�'��i�[_�C_*'ޝfsU�bĳ*�pa�޵�џ��<��>דz�I[�,3|#j4�$}Hj��X�� ��|:�D��y�tD���3�)�9@����L`	$�黾7:�M�Ǿ��]D��3ʶ�8�Ț^ӓ��:<s��(FG�����vTSu�>W/����|\@P�g�j+%ݽ>]M�#E�M���4�7-��^Vp��=U�y�pdX�snF�b�=�!P*k/ �D[���]�j���^�f�g
��CȚq�a	�=B�g�e1@�
���@�{S�I��U��_Mg�mq���`xL�B�z~�ܽͩ\��[�$�1{�{��y vhȕ���|����;*�\�d�Hݷy�s�x%/�2%iXڲ�9�2jIع���M��r]�]C`1jrH��%�'J&��rtEW�ZQ�n�+)7(F!'�?��?#�5f k��\dotw�T�Ѻ��iYC���BP8�A!�Ŗd�u+\C<7�;�Z f�y/S��ڜ)�X�UOTC}�6<r���J:���ӵ�m�Q60��_>R]�}�!k=	EO;n�l	5�E��G�4����8D�+�����% C㺍����|���,]R<�}�!�i����W��ޡS	�H��˲T���#��6V͵N#[�N�S��s�M�;�� �^&�m��`�
A�1�g�waC�`�[ͣ	_�Ĭ�R�a�n�}Phi�;ьu]�e���9�.��N`�����ꢱ����{�f�W�ٲi?&7�Fi����s�i��6J|D{T߮Jkw�f�Ĥ�b�44���B�t���c؜�s����(�:s�ҹf��l6�a8� ge�5��L���%�?;G}��4H���O����~�N/�?� �:s��0������?�(�.,��aŔ�Cu��z�}�Ѷ��{^s낖$ŷ-�:����8$���$t�������@�)�$��~�N�g�Y1/�vK5fH��<�=)�:��gL&h��c�9,�C�pǲ�T�zx�F�u�n�Т1�G�PU�?WN�� >_��]����'Uh�5}CAh(��B�{���a�[K��.�@��g5�̚���9w	�!M/�e4�Ӳ�)��*w�{���e*=���_�3!	/6��SN�6 ��-�lP�C|�C�!��V�N1��A��R���-�D����y f��uv����]�2Bkvz�f�	-"���Wq8k������������T�Ob���[��8�L�b�-�3����$����`VA(4�G"�D'^���VQi4�Ż�i�b_��v}r��۠���RI���~�'<D�^��>%�E��/�QA0;M(y�|*������_�W�]�0?�#�i��� y�S��1z[�ں�
dڐYcOg�G�_sLܱ&2�3Y��:��������	�8I�^ⶅ	���ਸ��vvB��L� �ɤ�}s6�����#_Z�����Y�����	!LPS��=��|	���/�s�����gq�_3��O��٦4�a~o&�+)���dq�R2bP��?���/ؿyTFz��io@Lxan��������Y���,���3'��Ŗ&cO~BH�^l�U��*�Z��K ��i���"���t�1,gi<��ȿ�m�zS��S���ǫV��(�	N��^�5���r�ŖPSQ�|��2k�gl���;�e�
��%��g�xBh�~S���k�b��#�Ⱥ�o�?)����������I����ᜅ�fVjٱ�s��E�dHr�9���v�k��Y��pGw��L3�D��0��R�7'w��:�ɒ�u��X�<j�pr��:O�>���[O�  ��EsS����F@��:o�u��?�aŊ`�X���(2��J��u����s��T]�
cOk	��d������YQ�+HNy�X�!�$�OP F�zn�2$�uD�R�*�oƄP:���ua)�!2|��"���&��L��u��Lc�Jn'ݍ�SՓ���q�?���8�ȓmK�n�@���P7;��1�ΰ��nJ^_د��Jf��lS(~ǭ+�e3����ƽW�LWh�N%�R�V�=�0,����`����49&�Xgo�}�&��6�G:��һ!r�R�3�h&8l��ӿ��9?ߪ���nĶ#�d��[j�͈G2���u��8DjJ�&����>�3l�j�e[�ѭ�RV2�]:�j�ڲ�C�$1�&�"�k�"kg��y�94�O���p��25����SV� ��U[��0�	����L�Z<^9�Q~�Id�\6������ԣ�������PV3���Y=(��ĭi�lJ�D�]i8E|���;{�}�L?��^� N������n������ e�<��e���.2xs�m��Q���؋���� S�i虂��c:̊����)_���Ryܦ8��g���ǵ�u7�G4)��h��&+j+�)Y�#W��ǽϙu�I� �wߎ���h�����b(�j� �4�| Bi��pP�y�|��A�&b�����B�R��M'�D�-l��e2*�����Ǆx�B����fg���-Vw����л#��9$�US�y�7�q�)���59����^Ĝ�֬Q���O�Wѽ����f�	y?�	��Y�5 �K|����T����r.��O[N#�z�u�}?�x�q�{��>��T$���.�����S�K� ��1�8�ρو6�K��T�)���y�5q%�������U�3�T�%JBCgQ<��Ob�0�v��ĥ|d�wCW �����s|��/�6 ���u��}R������h�"������J�*��{���ùrs.{B|:7�����tU+<4�S��mU�N��r_�`P���h�q6jLصb�9ͻR��
�Ş�dAc'��3= ���P�$��;fh�&nF�T��X�N"��~`p��8lzxf̻�z�'E������4�'�^$G8n�\�&nX�E�}^S���γE^�s�7�	��N��4��p�U��k��a���\w�C;!�K
�^��⨜��)����/߽3!��Γ� ��C�{�ߙ؛ՄZ1��"���چz+t�b��aw�2��6	~fF4����0�0Y�	�v32ψ�?G��X%��ۦ�������X�YB�z6}�s%ل}ȃ�|D��R?�7�#���z�#),� ��ƒ�b��j�p�� �7�k�3/���yq����j��`	a:e26�U�`���x������~ϡA��ȅ�L���'���$�� n���(:���\�@۫0��T��<�
MP,I�jon�H�M@��L��BH\��S7Xt�Ȁx���joh#a�-4�Ga�^��;Q��������ne�����:e5��4�zlP-���QH_*��pM(�e.��N� @�^�+2�T�Z♈cb��`V!�"���ۥ�	�A����Ί�gOU�cϘ	�t��AS��91�ٗZ��. ��R"�@�4����V�e�<��4��H.�`�bbl�g����N �����b��8���ߋ��i�W��m�D�>v>Pf��gt����D= �5$%�p�D��$-��&�sM�Yo�!9��$�H�fL�@/^
��bg�^r	!�E�!�V^��jԬF;�L��Fp#�;���� n!,�L�>����m�]�G%Q���4��<0��3���zǈ�g�r������/��z����Q��,?;�VE]<Պ�!6!����Eً�j}7��$�c�.cew�7dt͎��PD]!<>�W�r��Y>E���Q-v3��	���^HJ);o�u_�L�nnV�Q� >y�`�u�Ъ�T�	Y�4dpB�U�>��k�7��7��N\p��v� wC���o��Il=w� R3��ka.�d,�B����M�Xě?x�yG��yr1���h��^~x�{�*#l�*��4Nח��C�!K����������z��C:Y*���O� �ޢ�}'�OK�N�_ ͛=S	�Kz�����9�lŲ�[�r�a�ơ������
V5���Z{zIt�_���ii�0
�O������#7�^��]=�/�ni!��0(�8��C�}I0�1�L�n����mR1(��@۔|��/�x�o������.��7��O�ʙ�̦-��+�ǽw2�:������X�iX�;&؃�	���N$x9�ta.&�P�V�GM��S�4��Ծ �fc��[Pd5�����:���.�YUnު���0&�B������]��~u;����m�=*��:�4ܝ�U}A�H"�LO�\��;5�>�6~��c ЃgZ2Kx6���u�� R�K�޽�G��O�>[� i,I[D�"ѕ.�qw8�=[k�	�`�A��`�P�u㪺֖9Lv
7y�@��e �*N�ր�!*�r�pp2�'k��9�b�]��wV�o���i�}[{�m���}-��{����O�.�{WΡu&(�x)#��)X��@���]L��V��w⣉�j����.|t�z~���M�x���	������r�M"��� �8�6���+A�_�1�ɕ3��L���#�~ʥU��,���^d�<x5�%'����8ҕ$�~ot˾
�]���Y��W�H��Hp�}�p�s�Xprk�=����0��i��0���������-�>�X�5����:ŘVHt?.'QϞט���]Wّ�	;k�.V1{��T�gh���@��[��(d���94��״I�hh�{�L�s�N;ts�.d�o^�&�q{���*m�}��8�m8Z5Ӑ�fցX�3i��$��yq�j���ٿE �ji�M�a&�� �ӤP�4[	S�H�\ma6+�8X�+�d �jI��"���H���Vl�'c�� p4���l��T�tb���"�������7S�æ!�>)��_�����ަ�0��k$�韼<�3kc��]t�"z��4"�lb��ΫvATi��B�<H"��|��-�;k��<�ˡ���Hi{�(�L���a G�Gk�=uH�r�̻w�>���@]ЇL��w���V�5�����&�����R�Mt�h�v;s�E�+��	�n#ծ�R��+F�g6W��<ӝ���Rb���_@}����#��"�=��ڟ��a@�BT��2�a�W�p*[N�U��؂k>0\���n%�u�D���
��ս6�g��ŏ�Ap/C���a���Z�/������Λ�.�D�%ђA�H�8B��o.�a��jE��Sȳ�o3��_�Ny_�Q�J�[��4���qd`�"H�(~������]JWe�0?H�1����1�PR�Ӛ��
�EO�դ��l�6���	��C����>oG�(�\��\�Wo�h�b�z����+rw��?(BA�s��@at��� ��&�{,*�<?<�g-0x*5�}�#�;RB.�]����X�s*z�����C�% �J�IY��3oÕ����\9�h�s�,����]�<����⿞BĆ�LC����ġz*z"�����i\yT:Zᦤ?ka֬F<Q�9:�'E_-��|�i&'a���d������Y}ߗ���yz8�!�a�YY��(s�s�Pn��6�L��O��NB��tq�?���7��n��6^1�Tx��(�^��a��P*ф�O#��ۈ>g�#^&�ŗ��4�L���-c��8l�۲�e�6G�W*���V�Q�L���m��l���^�� ��������j�D����2��K�e��i�5��o'��m._n��yU���7/h�����Q�S��)R�K�9�����O���c�`�GI�v&�J�R���8PE�����a{j@���< �|��KVې�G�U��n�K��X����5,�yJS6�\�ib���k�>p����"����"^�g�|U?A�v��,2���X���_N�C����N�!��)���{]��"s�k�|I�Ӹ�1��u�C��Y�si-[I�&xs=51W��+̯��Z�Q
�� ��_Ț�c�Yׯ�
�S0�>���_��q�b�P�6��BN��G�@@�V��L"�{�yq��R.l�6�����]�2<6���}�-�3�@2��o$��Њ�|�����!z�2볖����bCje�;L5H����Q�;H��$��ȸh�e��^Z)�4b��{�B�!kR>�3A�ֆe�rAAJ�[�u$�y��I��	}�&���GKҜ����́�ż!nƙ<qJ�d�	�ь2m�8u�s =A��$��wn�h�I�� ��K(��7o���7��+DJ�:/��o��G���saF��k^@�35 ��yj��e��T]�o��&	�mD��|hK��a�܁��4�˫�UL N��������?�\�Cχ<?����"��F}#���)�E��sR���F�Ee�W0`Q͎�x.(p"m<�/W�
vb3*9��xŐl ����b�(&Y���������hVr�W%���Ǎ�1G�c ]}{c�?�O�9fC�CD�ޅ\�'ij�>�ӻ�H�lFnT�1S���3���A�T��|�Y��r��Ȳq�Q�/��`j���Um��+���V�yl��ѽ?K,�����b=�i|�2�2_ZN3-O�2/�|z�$���5�Ji� ")���&5�
3�!k�v��1���5�C���4b�J�9j��K7���Ul����,5�<F���W�d,1�d�Lo����a񙏋؝0��>	��쨣��]̉�w!���j��ఖy+�]���?����id�j���	�lT��ʪ�.v7M��U�4n��uힰ,IB}B�A��i(p=9�`W�y*a8�%%�1:߸�\�SWc����@�pf��, j���i.��LI�`N�w~H��X� ����7�Ӕ.��"�4���L�{|	*�����0�zv�S��-f�O֞�f��q�\t�K�>/%�Əbo�I�DP�\ح���nw�O
41�~,)5>uj��M`��p ��@sY�YE���ZX�������W��+Q%^�A��gJ�FP	��;o1��@Y��X�����^F�ǐ��������l��ײC����s��׫��v�*���Xb��t�2�����d���+����(Q�+*^�3���'�+e �2ݴ5�Y��^�ǪTfu���r|�h�?���X 9� +ܚ,�:m�ŵ3��Mf�Ȅcq�lCZbW1�B��?��:&�'˛#ސ���#�0�*�e�7u�N�E�C�+������A�\ ٢�.� �,~�j
��L�������ͧ��EG����;��EK/��p���]�{�k���c��{I��)j��<��a"U��A+��m��9$�yt��h�w1�jRk� 9˥���En	���Vz��}�|(�1ԍA��
?���`hE���ZUF�cwo��A�[�VH�-���eߣ�-�^s�ݓ���a�Wi�c5���[�w0����&�7'���.�H?q(�� I�\��u�V�����&�����Ƥ���$�e�k�U�cj�o�lqW�p�csI��$[��y"��ֆyЉ��g~8{�*ĒA�U�򼼈ځ�� 	r���I�*8G�4�Y��cy�#S��h^ Qn�-.��@�* HK�{��,c�By-�M]FZ� ��*0W��f�t.�V)�:��Uڗ\�R���cЈ>r�C�wu8=Ƥ#���t�w[��	T�?k�V�c�oH+i01ѣG��	���ˀ��lC{��1 X�ۢr�,�!�����	�}�P�fc�|Sk�P{�l������ԣXRl#Dy�k�(��4�tg�?�����6���,����T�I��	T%����g,eߕ@1�bD������V�
�sd���&���&p�╓��*��3j�{��C�d��I��3�� 54���B``z����Ϟ�d;.�	-�{����z�ym�	�������.VF%.E��*���Y��
�4�u ���sp��]��yz��NI�����0�G�2�_$�	��(%!��vh���"���}8[T0��c/�k��g�pLƬ��ϪB���N#˟��˹�}.�E�E����6n]3�8Ԭ	4E��(px>����m���h�t����}����(��O�4�r�0�gl\,r��vW������2�	z~!J�Z����N���,�W��Zv�$�����g��pth�VΕ���:ѱ�-��W&>ɗ�z���.�=�ˑKb}�2 ��)��<���u��f��oVd�f���5�����M
���*/�16g��ݽ9�x�-o��j�X풒�o�,��w�&UO��*}��ñ�(-L~�9���Av�  �ӵ_J�
�J�5p��He����7�hh��g�7Pa�N�S����ݥ\Іkd(�(�NtE${�G߱��F����	�
g&�&���I��d��"�^͙�����	��?TX9T~;�.x�4�rJOI"@Ŵ���ûi��#�Sܕ�R#���U� DmK�#x�b=����oH�;3��8Ƨq�t]��p���
,&K��ݕ�ٟב�(R+֪�9���%L�7���!�[����鳓a�}ݼ���T
���oa
���j3g�<J�4Ҫ�mؖp��O*J�Z��'Mݿ�97�ǡ�y�5�͗��te�R�-���tsR���\A�&Cey@���~�h��@�������X�حO�g����Ձ�} �Z����"��̓g�_z�ʾ,�٠r��؜*_I_$X��6�s�ahާ>��(R/,��ߊN���k�i<�Ry�9�η��X<�������E�Y��Ŵ���L����Vԥ_���ysoa'c���l�E	�aD�͉�3���}�������Z��&�]
���<�����?L4�����[�T:�U�Z�J������F�B�߁~�|-��)���R���ZN5}�>g�[;@3\�E�JI�MB"���E�N���|�7�;Y�9Ly���(rR��p�q��rL��� �x�.�9�e� (���j���)aP�*AӖ�Y�P�o��8Ͷ��T�m���[כq�na7d<r%����/�-u���T&���_�4nOL���(p��戆1�:�k�ӕ�ٯ7�E��s[�\ "�Wˉj+3��w�_D��ޮ=���cq�}i*��N�b�o>�HDG� 1��},���@\ېz���㴤���d��S�5�O��
�n�M�W+��0J����bx��$�X�)^b�Ƃ��;B����?��eHς|ä7�4���G�5 �����Tݶ�zk!�`���p��/��اĪX�aQTt&�����KT �{*�M��ۮ�����v$���d��?��ٳn���Y�=P�M���ݰ`-��ULvD�����U7��I�u�R��AH����'��ᚈ��!x�T�J���'���ZP�*� ��5���� �刘`.F���]�]5���G�Mj��5Ж�4s����	���?�A⧪4s�5T�
VOIA��P3S�(`^�>&�]�ML�uV��h��z�؝@{�=AJSO���{g�oii-��@����ghZ%R�;��/É�������F��$7X�G,慎�+M��(�+T��w�x0�d�s$WB'�d~f�Q|��w'��� ��TIƈJ!���)�f�1�~𗶴䟤�[�A��c2�E��}xw[W���M@| R����t��N���Yd����&=��OxHݓ�����t�X"�W* ����6��2Q����͸��Ay�ڱ�|�SE޻������݂?Ė�dm
��Eq���B�g�|� a�U`f�Ϋ���\�/=�E��X��)�3��(:��
ޣX��O��l�]JВ�at���&��2B�����������ye7?=�u�{�����n�38w� S��#�(p�@��-�T}	e���|P�`��eϨ����M�Q����us1��°\�T&�;�b_s1_F�LW�]v��,ˮLB����CD:��'���_j|�U�C�R��t��N�@H��QV3n����#��l��'\�s���J2_o��������u��(Y6 $�\��-$�w@ »�C+�uh(��[+��5�����G�Q07��F`�%�m0}��3�)/G���U,8�q?F�p*�jTV	W����В6��?B@s�e.��ttmU9E-�U@��1�q�߯>��X�3�6�K̬3��gʌ���0����(05:h��z|���ڨS�����}��'����Jn�Lv�yo�{�4���(�mB���7Z��3��w����K'�v�p��Xm8^w�����NPP�DPi�[�@���X�d�)״��y�N�֭�Q�^�D�]�DV�a~ң�!|dJ<oa/�z�۽�0?R�Ԧ|+���TǊ͇P�~ww�fҰ};"I��H?(��M�bB��1:��x� 	d����4�_����Ƙ[$��)����B���CI���z�%xh#�;��D�<֛�ǹe��n�G�ꃒ<|����� k���e=?%��0�隞Ƽ��o<�0�I��:����6�`6螞2�_c2$�4K6.1xVi��Y�hʈ��7'����9qǓԥ+��2����@2.��Q��}Þ�>�����۬8��\ۓ���рYl�+W�
|ZN?���b��K�/�fcy`MG:���t�Y�0%��2��Ņh�+$KG�N�=����M�3�~��5�qSjf�	�+�`$���Z�o��}��d�pgyn���p&^=n�H�2�oIԇ����{@H,,0�7vu��;iɉ���B@e�q�i�w�⻑�$뷣 kf�ҧB۬ ��(��Y:�s���"�HN�JP�{6m�wj�J5Ǉ�#��.�iy<���`��D�$�鼵��=˳"-ڹ-ɖ	a` �GavG�҂�K�x��j�}�	��L��2,8@��|Ç���#�O��A�2���D�5 Cr�<��/���@�*1�Sz�J>/���4�0z��y�'b5�a �����Ĭ��.g�;������ \HҎ�Qr�&3'
�3��]g��"�-��8'�4���)Ƕ|<��?�OW�'U�5v�����2SN��H %�����F��ows=���-`�)=)-�����%�"V=�����?WpY���h�(irYa�Km��1]J'�7G�{<�D>{��pS��Jlq�C� (ЊwuA7Q¼x���1@)�,�2ԝ&�
��B�m�3[�9��f*?Е.X�D���\p=������O:�p��`���|1W��&��A�=Eߑ@�l�!�v�KP���Ӱtn(��5��_�{$a�
B��H���,[���������(�[cIB8��
܁��J�k�Eu����Z�Yհ��!rr/Ph쓞�!���4ͥũwHv[�7v1�KE&�EM$���� c��B��]�5��u ��g���0Nӵ��F-4A�����#�':ou��_Ց˶��y:P�b�(���_�\܇y�����-4��S�=H"._����8)�#�*���̽���Q����dn�㘜��#����\�C�{�J��'rІ[�Eu�
�XH+�$בCH �,݃`��Yg�\v�c���F��n(Į�&לB<�K��x�
�4���S�%����GHB��t��r�'��~��#q�&���`�	��@(�~��G9a"�/8%�ja��=��C�I�D��=,����v����h�oD��U�&�A�Y뚿��x�e8����b0��:��I��D�#)�4�NKR���"�٭5�>?ޟ5;6�$�n��	�R��{zمV	�-)uh��\�����0���TXl�[$؊HE���М���~SU�,vi���f���[�?D���+ט����\�Q)�'��zKF�m#�.�+�B�)ץV� =��v�S�K�{��w4@,�nyYƁ�6�:�/�s������,8�.�0��ـ��>�IX�9���d������YV:;Wĳ�Ҧ����oI��ä����9l�Ke%2�WYէ ��p��yNI�ce<�NXwR�6<R�ý�� ����]�h.㿊������M�^R+���>1���?AW�����X'.t"4�1�z�mg�yX��
Nq�2�U=}�E#_k��RI,ɨ2
�K��M{x�>+GE�\�QH`�%|����`sq�J���;�&�Tlల�0K�1bj9;�i��O"5�6>g���?{]-���G���QE�� F[m�Q��P��`Z�������yC��"vUZ�x���=0�*+��́A�M���M��}��hڌ{��Qѱ���(�#GSR8�ZA[��{I�o(g��Q|��"?Qg��G�Ʌ$���\I�t�:F�̣�y�0QgurYeRc��Joo"@���e�$�����|ͪ1�x�i�>���>���Ųjr���������eް\�z�!ysF���������@0?q.pD��rYY��PL{�q9�d����/�3���C[��[��rQV���m,q�+d�dQ���uT���;۽��w�ȴ�+.6TWd��Ņ:��/iH�O@&���m٤����2��ޑ�;�`��.��^�۶��m�O_��ˍ\u�C_�C�!#��MB
��K-��OD �5�����|��k4����%���rDy��`�_@�Qg�c1��\����^�ȠQ�8��d����G|r$�O�v��D�c��#m�O�Ҏ���|��Dn%���B�u
�c�\���q���!0ϔi�z+�v!o��=�^󺑫)v�����YH��op.`d�6�G*{�%�-X_�$��Xy<�C�W[o�K��~4��H�,���+�u+@T���Al�^�W�N�t�-O��APef,�ik�>�.4�|vYrP�4�v��q�mmbb;� �Gk�5X��Qu��s�@=��H��u�2�j�ς~3M���Z���P5%,�S�MP
�+\(�D̘���ú�5ƣ*�t�;ڈ����%�]�7%o'�ɍS�p,"���B�ш },>w�~���y�%�*�6��sU\�7�4`[ 
b	��Tn����X��̾t'�wS!wa����}�˓� ��tL�8b�3k%��x\��Nt�i���^*L�s}�\�G�V�:vLd���z�/)罞 �[Q��3*G�Rz��a�|+~�z��I�bN�+X�J�x���K���n#��	��QʉA���Ѣ#����2rPuط��M��W�x�·P�_�p���ISq ���'TfB�bԢ�(�>5D'���r��GwHT�=[�b �o9�L�z�_�6=�Vd�����ݒ��9�4������{�|jP�v�LK#F1��sG�^~X�����Nҥ �l��'��x����Xe^�����Z�I7�T��Tر��iQ��0	�ݎ�aߞ[��1��6rS������Z�<�ʆ�(���MP��l��i�FY�I��Q��<g���(��٤#�������P�y��+n���Z�	2K
;%�{>��e�[�����ǩ���Ok��ms�t�\� �U� f򮮈=$�]"i9?9d�v�._m�Mn����r��/f&'����+�$������N�=���i�W�O�{?�T�J�����K΂��r~m��h/:��7���y'�.P�ʋ^ۖ���HFvڥt���C��uU����}��	s���ی<][+��/�0:�����d)��&�����ʝ����7�ةA�h�H=Jоv��N���gڙ�v� ��@�@��Ф��%*�ލk�E�/�/Ln��R�5�f"x�Xq�Ha��K�S!)�tuw&z �Ƈ-!i5���Gq�^�	5��������`ed׊Ïg�2v��9Z�1�3�:��>��U%�b���Q�Rm���}�M�Ut{%���>���&��ˏ�����h���+7g��Z�@z͈��z�+�Q(�ˡk�_.��;�A�r�te�3
!4����J~i�!���C�3V�Վ2#�\�6��1n(ZG�0
���K��g�Q#���%9� ߖ:�+�C���<J���ՄV
�����Q_{�bUj�;<	���>��\�����e���bl�#K�_F�R4�@�X�߆���c��K"�!@��*'� լ=]���B�� [�~ Q]`x��8ZE��J��{��<æ�N�Ks���E�ಝL�$2!�.�G|<0����ok"�~Rބ��!�9c6�e����7���7]�l�/�1+zﲠ�$�`}������@�L���,����C���aliȰ�:�@-F�)���N'c��,�����x�86�H�<9p�L��T�,O����E��`�i��^)'�PxW���=�0d~�z:R�E�L\K@�ą4�Y,�aʟ?��'l��/����a/e��oė,�G	�z�0��a�ߘ0���rA��6�\�|�������+���ԧ�_�}aKE��m�2͂{ދ��� ���?|���՝���Jg�ǣBnV���C��a���7�YDE�sj�P�7�g��OH�K�xx�?���S)��=X!���r�x�b�g��+Zʷ"������vk@ж8�mG�0�B��mIA�C����*KXIi�p���X4f$�5���X�8��{\����pF���� *KC��cN�5�i����E7i�Or]�tb��@��PT{��,0�|��ψ��B,�M�k�^�=$��*)��p�0=
+C�%ϋ��u��ʜBTJ�H�՞�J&-x��#�3�:uř�[c/9��QnZ310?�2��u�W+
)F�
(d �o���}C�x)�(c�+˥, 5�a�2�J��j,���e��+�F����]�W�a[��0,ݚkBKC4�G����V�>ͥE/���Y+߮UC(���ɰ�BYIhnc,�Q[�<DMw�k���Oǿ�ą��5��B��f��'2�.̣.�F~U�F���Ҿ`�x!�'ac������,=�!��ؐ/�]z?��*�^~����^6)l�j��g��,T���;��rߞ���	,���(�˓�C���=C�ا�űXG�ߞ���R�	N�I��^]`L�=�
������b�,�!!-(s���!�K�ɓMI@O=m��٪ذ��xA���Bȡ��p����9(,��B�<��A�,�a�n��<�x���C���!x�u��79�6�,arG{�>����Z��,a��XT��&u�X�V����6FTv �e_��6��F�����.���<_�CE�Fm17�(Q�=�#v;*��H��'��֏5Ƿi��u��ir��e�B�pw���*��+�Li�p��7�j�ҝ�p?�i�����rd���dXRh�"n�L���_��:��J]hߌs@e3	5ä�d׶HU��/|c)��*�J~�~�gw�����G��bSÑM��(˦v͏��DlXe
i
(�_�Nz�_&�@��7R*�o(��֑?�ɷnĆ��\zx�t��Lo�o��� ��caҡP����	P�,�0�u��&* u
��c_��K(8) Y=j�����t|}&�a���;v9O%~�в���� �w�N�=��>��2rļ�H~ -W�G����.��+��轨Rf������L�ї`y;F��ćFC����X������^��+��!ld$�;���$�G��B�ڵa� ���1By�-��һ���8o�$��E2�6�?e�Z���w悉�z�b�d�M\�+=�v���n�C���B��u�B~�#�ְZ�~3u9��em��,�#߁�ƹ�y3�B�K;��$�l!���Oq%����8{/c��ē��RTnQ<� �:h72D�¡odo�OP V7�����<&��M�A��گ�*��[�y���_j��Џ���tIh	;6d���k��-��z�|sX�	|�i#���37�0<�(i}�X�57eg
�CG�L~�j�ET1���Şl#2����?@�\����I�s����8F�3�%�����O��e3mq|EA#�������Թw�^d�se�����G���b��Q4����a(2[5d��ԓ�]aؙT��wZQ��(�x��йb�1Ff��`_N w�ů��&U?�c�O�-m�+���~���R�M���m&ɺ'��%�x�LP�'�s�����dA��%g���x�6"������Q�<�����7���I��r������-۞�G�����6�!!�֑�d�]����į! G`�/���Zo�������PLr$�ğˤ�Y�/��w�4A��O�i5�]g�귇�1oAN�`����8`��Z�K�e���|oڕ郙�
���zL��� �C*�n��{9���ǫ�$�`�M���p
s;S���C�{����`�a�ʹv�SQ�)�(]������}����`��4c��N��"�H_f���)��ⲅD�H��P�<�5`$�$��}�EW	= �1+���"�y Ă�TX�ͼԲ�\�f$����	�V�īl{b'�g���2�{Mp_�ѽ�+�*I�ߎy�X��0�Jco��Kظ'��@ ÓM'Zy�FJ!����f����x�*)��NA=����W�	r2o��
�Y˲��
��a�D�>���/���F�4��\Ue���@�ϲd�F�����"���9�ay6������П�����2#��@D�.-8i�Y�Q���q$V{.�S��*�4�݋�I�����m�XF�`�K�_�!
Eѳ6�)z�	���e.Ҳ'fp[��f���с;L�׶�"D�4�Lf���x�a�t"|]���W��g�|Z��"��G*�7���0ҁ���j�*=�*M0�j�GR	�c�c6#%[�"A6N�L��z��)�66)?��fǛ���	�M��0������ñnrnB�+RfkE�=�J��1_k�:o;�S�F��Or�#�Z���j�����@� ���E AY���Ea,��y��B`,9��:5i �^@h�d��g�ۀ0�Y[�e���'yKe*���p	b���`n5�� �kVD�I��u��� a��%F�aq�y(�hc/2���_l����v�(N`�N��P!$��pX�?
:H�="+.�������jB��T&�F>�ؑL�Wy��cB�i־J"��\�N<E!r��{��}'���,e�ِ*B.I�V�%o�lf��3����Q�\�b
���kI���1v�Ǐ�[����9��Ugj��*�I��@�CM�R<�����2�ҷ[�~7���Ϲ�(,�����4-@���A�^H� ��#�n{��p�S@^�T����КCF�*/�.�&�?71k��u��&�<o��\���J_��]�$�2��W��3x�xK"�I����$˺ͺ����3<Gc�5g��		��k�IS�>�!��T�c�o� X�Յ�l7"t���U9B���N'j�I����0g`���m&���g.+��_�70��I�������T0ʷ��v��ʊ�<��t;���]K�k��rt��%��(��:f�4K�}��c�`˾�����;�jFTv���X�^�����g8�5��;�>No����0㻶�z�[!��:$�ϣ�-�F����c��EK����k��RG����u�	���ţ��v�e'�=�G�����������ܧ���g*�'hx+>*�͕"�&H-3_bV]����U/o)a���ނ~�:�PJtLD�#��5��2���B�^�m�J�I�=�(�?X'�����ExD��op;���� �<.}ƭ��{f�eb_(/i�aƓ�y�������y�Mqt)�VDa���ۚ�� 3l�RM���M�,u���A���[0��#r��21^��@���X�.��"�O4�<�ޔ}����V�@�4�xoG�9�6Y�)4rV*��T�	���Љ��X���[D����h!�`\��4��v:�3l
�0�1ݷ�a�ެ��I�{ɡ������j�a��J=:��!\���A]��pj,�B���S&u�ɥ`�D���v�%��N�~^���lz��?�(������Ŝ�@�
�<J�jt��/z�PU�V�N��Ђ���V�BK�|v�W4���u"%&����9�+��%� �s��Bq�8E7oz���ي�6
r=0A��.P�h���D�s�%@5"�m&XYs�6�o���8R���o���G*���>�o;(�0�9�#j�t�o�Sm��"d��i���`�e�e��G�>r�`ѳ�\�I�?�?6�h�����n8�4��*��<�9�g��ݳj+h�XzG9nn2�C>�-6ώ�pwd�>����s�����$��-��mTm!�yH¿'i/K_L�'�����ܪ6��6��5_�U��,�.h��9Y��U-�"=t[9���v9��~�a�Y�3�#�5���6��s���ɫ?T����*�ً�p��B�x^�x���2bs�Z|���* ?1`[��dP�ű��ޤ)��7�x��t�F�<��Voż��G�5?2���f T��1�l�?��YD�}�ru�ʇEH�a�D_%f��J���5�`=�ΰİ�/7[>��j�5u2*�#
` A��:����#M�r� ��
��\��g���i�nPjO1<����]�|-S5=�	��\��sʵ��W�Ӆ�Y�<�/MY���X瘋͌vRxA�˫�z�0�K=�nڱ�о��T�P7�7�u����ޱG���'�X.�r�7���m�r���3N���ʮ�]����	!���U�D�)Pщ	�2�S��K$1�x����#��>�_�7l3����%�ѭ����PL�|�����]��-.�]<�Ǝ�IT+P���̶�x���W� M\�P9-�߁)�.�{�G-��Q�1��an�V�m�Ǽmm�D�hS�v�"jC���,�W&h�JWW�&*���`Rсb ����s�0!9�r(���1�0Ԟ��5ݑ��[���4��U���0�v2^�e�G�?�D�rY*��Yפ5]LN�H��M��qL~1T2:8��S@M�Q�W�s�h�-1)+��چ�qj��V���U{�K:Xn��T&�`�#�It�e ��bb`U?	ʊ/�Z	�F�Y����%.Q���B��x��nV�|t,��h��L���*�^�Ζ�z�W4��!���׳m0N��3&�*����e���[㴄ύ�X��5�ƻ��o�F�(�u�f/�
;�sIEy&r�Č�	4hd�$��@��4�3�p81��tZ�<��(�Q4W�v�2I*e������<M�|�b�qҧ9[t�� �I���0+���>8��!�o-��sx������Z�#�0#U��.a��t��9g���-����A�
�����=^q�D�ʹ��w: ����~���r)�Gp⑈��Q5���л�q�E2�(��4���~�<`G������#�I�KU3&~�xO�3��^;
A.(*��R�l�%��״��g�i�k8�SW*aA<���+5x��Hr����gQX�g��n��|T�3��R��7"]7���pu��a#\uF���a48�?z�;J�!Ab�g�f2�q�w	�"8ۤ�xF�X�,��B'�5�F���x�,)^�oC�R�s_y��4jH��e��u�m6���:(�3�	�m�u�o�����+?�%㦹���&�#T�i���T�i,৒�/DW%nWno<�c���E6:� �hd��L�-�u�Ҕ#YgA�J������O1ä%쳊�1�RϾ�V�0Fv߿:Ly�Yi��K�]�71�����K����ՅFjˊ������65�gl�����\/e�4gG��
�[8�/*M���7��٦�1��ణ�3�e�֟��#�7K�?/��[:C�fM�:c��@`{/�TL�jÚ�Y�ztg-	�����z#��ܥE.�n�`��p����22�����C��ot(�`$����jƾ)�b�R���
&1O�G�h��̕����s,��5��Խ�A�'�%a	Ӷ�Ҍ=Ɏ��%X	UC�9��1�/O�5oSf�K����!��Z�3�Z`ö;}ܨ��г�oԅ���J�z|��]?;`�F��)�{�����9��3g�,���>�R��[Z�J�~���bS�/U^�C�������X*�l˻rg&���54ܤ�m6
-���`�t����ɰ��[&�9�o�B���g�J��xA8Z��x��ך�R}�I��R�����\�*�.$�� +h����j�9�d��_�����n�B�c�Q���F�����ɕ+R/��p��\4 O��n�@?���7(5�E�Cϥ���i��l˲o��K�[=��Ӧ����m,�;��S� ydfd���x���Һ�5@}<�\���+����^'��!�,��:in���x��WT����\��S�{f�n{n�P����5��k��Ⱥ�,��pd�Z�*�Rz
��4=��t�X˹��)z{%3}MǤ��r4��7?\��[;0���_�ry��%��������S&ħ �^.�{jÂ/�%�?5���ݤϴ�?`B$��(�|�����[p[>��峰;���`��6��1?�CH��2��ȱ��#���FX]ωͥ�h�8�b�WmT6S��Rn�[U�1 {��xyA��cN+j�w�[�d���P��~TI%C끷s��Ż��D5:�y��Z�뷒%��"މ�, ���|���d��ZZ�U�!Đ��,�.b@�1dE�4h9���<�����	8��HЮOg��0���������P�,&Y�%����j�����f��1I��m����C.�ȷ��ԩ��ڸD��Mةd��s�:��4�y�T�E5�2�H����:��dZ94:�&�%M�x�c�ef;�uV��㲕�?@�S�V,q�H�0b�ޮ0@Lڄ(};����T;a��O�u���YNz~��H&��q�-�Y��1����Bs�/�>1,��?�4}�}���B�<� f�Q׸�h�Xd���u�o�7�G�9I�9 yxAJÍ�w�O_�,�������G���whL��T��٢v�u��Yj�ݚ�׮]�Xgӌ�O�`!F]���-��k�,�S�W�
|��ȁ�A�bA��]��'T"x�Ѯ�.N�ˡ����uBD!�+]n,��6���F���&;19��r).��ϧ��-�EN�h�4������\HF�;t��7�=L[\�)E]xY�:Y�/�
�����tyV���T�9GH����ҀP*#:��6�:W���k[??�]���xj��H8<�Sh�Ng�t����tF"P��Z5$Aj�r:ٲ�����*������
v�&{�wVx��� >��y�K/31R�o"��3���;{LmP�(��:�]埬G��K��w:�����!���f��Ԙ�"��?~[����)�n�
��0�R�:�P��-�<8��y�>�_�q<��R`�����5V0G��@�e�Xj�`y�2�>:P<#A��Rbբ�Q��|��,	R�cv ���BYC�)��az�#�o��t���8=q�5��`�*V,
����6X���Q���L�;��hz���������+}���(G�H�|���#����=t ���_X�F�`I%���U�w1�jd��bR����`���]ë���`'�7X�P	�jn�.E��n�)Ou�`W�>����7���iP&�N_F�Hw^����2;�"�C��c/	����c��3�kf%�+��̱v�>6�C��$	��S.��y#�t�y95,���d�����9�&�5/�����c�!{�� ��P&މ?�����a*t�$) �}I�p8�
��Q;����<sʮި�pA�5i��C[F�\�'��?��9�!����LbOC�<�6�u
�}�'��ȎPK���[Q
7�`a�a��T�������<D��������?�3�}��	�O�&wi��ѱ��*�5/�@>��� ��r�%qW���ܾ[�]�{d���I��t�g
"���3�}�7�h{u��)���?�����f�g��	/���׺x�|gȄ!��B3��?ڪ{'s��Ho\��JV}o�-}��߮�q�#�K�=�"A�x+�k�Vh��hi?I<��֣-�J��������a�v!!��cg��o���g�?���Ӻkl�:�̒��p՞���r�/g���	�si�*����i&���P��,~~HK�>G�y[�U��r(A�%�ǵr6W�ED�5�y>.�	D>m����!Q�"�S�)Z̓�.����tY��t#�gxͻ�3H(�@���E��f�G|��Z�jh"�q-uf_)����2S��=ӧ�s��T�X��آ���h5Yg��`�7��~��g�M�鋧��s�Й��>t��COw�A ��R����䭩Z�w��-��!��z�T`�4}�ݽ���9�l����~a����&TB���j!;nU�J�����g�D�hm�}o&��L٤���B�Du^�/a�@�y�Qӳ�qS�l2t=AOqS Ħ��.�Bmq��U�Y�p�Rp�
Z5f���-�F���N[8�G�D}��V���Gc$�ua�%�ɉ2���p+ҳ^�F0�[A�WR�;�k[�v��Ih-��1T�cC���4.�դ�jv�n��T�e�u���*rC ��q����QZ���\���ü��k`���/ ���2Yxܣ����;�&-0�-�-�|!�WZ���Gq�X0k��*4��?X�3}r5�ؔ�晟nW�]�)[\+�ʡKT9��j'�O���R#{8g*IVМJt�_��ibƼ���R��y�� V�Mm��S+��	KB�U-x��v+Df2M[{�͵82��"� ���ɣ���=KR0դ�9K�~#t�VW��L��˦x�Ol)#��i�Ӻ��S)�t(�R���R�j�F(��<��O�����=�9��zr�$��x-�i�-��x�k }�9�FǊO 	���6-H-��g�^��`�Vԕ/����'T�<��R�D{c�6�w�.�a�_/E��D�_$r>�/8�v��B��s�Pա Y1�aX�Ba��\�U�`U({:N��]C<Uk|ٳiݫ�1��*1�������gI�A��NҒ6�.��c�Z��VX�%g�К{�(���I�w�V6���a�5��+�����Oc�l�{��$�yf25$tIk5�'��SO����d���u�=�|�onVm�z[�9F�a�/����}��d]�'׭>�kp�t�3�>0n׽T���2��6���\ '���Bo�ӌ},8o�꺿lvV����8�w���~KHP�3�{0��~�
ҵ��p򓲆�w��EZ'*�X⯋)#,�l�v+�?ٞ���>�ǔ�n��!i܉���%��p����wf�)�&���P0q�?V�bƅ>���>	����o����i�Zc{�"RLrǽ�:7�u)7
�G�`?���V�KW#?�d�u����4�M<1��s��DgO9��띎0��q��#3�H_T�YWy��R�Ε6˲�H��v�� �!���G����~�?D�؎��� V�����0��9�;C�����'x�Q9s~>&��F�qrf�����b�L�GͿK$ ���5��=H���LC�~�s��Nu�ö[(���R�"�(Jǈ�\���(�-¯�(�/�hg��ziD-}���r������_���~��7=�T��A�0���ի��	��ф���N��Z=�1oӽ�ȡ�m,�I��(�Hl�>��J𲀞#�^�u
�M�S�|�Z�xf��G�[.+�v�0��u�Wgfd{y��2A��ȸ㐐��ӿ7����1��W^��8W64����}����#9	��������},0��^R��<�2��,@��O~;�T;�q��?�3��\�u���W��v�Z>r�d���a�JF�m��\ D�,G)ڪF�o���i�y?nB�-эV�����~��aE����T���w~đ��X�h~��g�W	�|��3���`�a�����{�"��Skc"��U�uH+|��W׮(]e��~�4�&��O2˶�z�"6��u="��`��Τ�����'��M�B>�WH��e��gh���čtD<+�w?�$���So~��桒 U�O��v�W�������Q����f��ƒ��X�0a%�bMkj����xo�e������	f�&�\>������}�p�۵���[�䷎��dy���W<!S"L��*|;�_8�^���n��X����rcp�{Y7�M�Q;%����F*=UV����x��~�F�Lm���d�Κ ��j޹�y�����\���A <�๿���5 �TZ�2�ᦷ�z'\oK�K�ؕ"ݷ��`�6
��;�,�'�r��O|�?K����?,���d���v��6�6We;E�G�K�2L���̦cN�.ٗ���4�-�'l����FK�)ȋ�[#�ċ�*v�z>쌣�&�DD7����0������vU:,��4Xt�#�������?��MY#!��=L�:�g3��F5�ro�v;z�ɔBl�TPvá�P�dX��X�kJ���Z2l����4U�B�r���.qy�����l3��T�XFɟ>� �mɏm�S0��$Ah1�����13�H��Z����rx2����^Nf�y��]�-��̈_���%��2mk1�/y���Yt�P���[}�����$ʠ�t~v�U��$V�_�4O��6�3ڟ��g�SH2��(r�"���M����G,�����"��;$��`�M�"^c�h<��9��I-!ze�b�>�Kap �;�p�����5��������`�ǥ+U�B�Tz�/T��ԥ�ɹ�"�o��:0JhC��z��/�"(�R�'�Q��?�u��$gi��v�v��
�������	�IaUz�B���Q*�I�������1���}�IW�#A�{_J���7�g�R6h���� C���j��'�1�T��
�."\�;��H@p�N_F�-=4���C�~s������Rb�Ǿ;�LD�0�U2��|��`��J "޵J���ɳ.��n�8hx��s^M2Հ��F�,U�+�MU����$_a�\���X_A�S�Ę��|��܆���/>��TȀO�� �� �������1&D�
�[1��Z�ú���u!��BO�x��}�ǂ�܎������{~�M���l��W	0� %��[c�u��۵e�!�� ��>�h5)b���x�eG�&z��E���Ŝ���V `(�d����h(XC�������(#�g�ۮ���U����n����FW�V�Ȟy-\�����[���4���o�蕲n��̺.:T��"?B�"�����^�IT]�n������vО�X���8�}�Bgr:�x�5�z2"(� H$��z���a�ʔrALE*%x�a�j�5�IMP�p)�首�m�D��-�~Vw%�~B#������}��k̴�͉x�@�B����W��"����,燼@�}�r?Kr���j�D���x8�����WY�����}"&�vs�����'KmR���!��ތ���x�@�n�3�����mǟѠ����l��p�� �=�MjO����F�N�r٠�N�W{@��R��gg��3B�����!��Y}B	�^�sJ6���H��W+9n���e��O�:ۑ;-�U�����}Y�+����ҥ�z�Pc�£�{Ġ��/��!M�|�T��\��z;_������{:�k���U�o$1vt��'�:�Ȉ�_�`3T{`y1�]Y��W��/.�Q�s���ewG4ƙ�B�y"ew��?Tc��t�?�1�#⤚��4ޖ�GDKY�Oq��A��ID7������Ák���;)�����_	��紌+��1��'�vA����$ڪQo���}�1qM���t�K��^��	s�� ,%�U�k��nG<��㓒�Ap�2[��/��)�.g%�@�?>3����	c���N��*����ad,����ސ����4�����w��!���fov��|��	�⊟��]��B��M�K1��r?b��6C4Vd�_rK�^���A�����\��7n4��^cvNh�8;�F�!G`��y6��j�qp�Y�c���?Uڅ9�f�(�	C(���!��%E�6�S��um��5.϶���"]�Q��Y�J��u~g�נq8d#3	�xPo���V[��}
������V�|3�<�^8��=�B-���zWmX7�\�^�G�c��Eu������j��*I�yȕ ����1J����I��}���2I	�H���-9�B�*,Y��!���^�A?�݀�B�S�V���)�#!�Ʊ�w�������$�U�	��J2,	��
U���l�1ڏ�9�n����m�' Z��
x�iP9�� a�ڦ�Z���|[�\̳\��˿?�J���{�^i�nm��%h(�h�|{�[��>p�����D ����9 mX�+{�����Ux��[Y#o����w�x�/>;�˲�K��5ή��B_�q=}�X�V��>�����T��a)�!���8Y� �B�u�P3�iƒ�`�'��{�{�G��'����''��_ۉ(~�G˦��W����]U
+�2O��|$TmL&%�קV�F �K�M��}��UI3�j(�$%��_�!�f�J���)�v\$js��,��<����|M�q��y���)'#+�0�h����d�6������;ð
c�kù�а�o�#��0:?W1e����1�t���[@N^q���2���v�����Wj����w�0��m+[�k�\�Ճ��w��,4Ļo�}c�u���rHnO(�lNw<]�#ڀ۔a5c����k�v�4����%ۜ�����BW�y�v��k=�1�O�sq`��%r�6Ε�p�_07C4Ҵ���b��<��	��9�������	S2�MU왙�����g�4�H���@����X�P�־�m�I�����V@�R��i�����L�3n�	ߝr����{��R��c�{�0�����=V�2�[|(4�s�B
��h5H�q�E�����5Bo~pb]b!�W0��j܄���e�7������e�h�Fϵs�<p�Y=� �0��yӲf�0鐍�"��U����
��c�Ϝ�JC����I|"]lք��fs�0L���Uj��F����V�9�S;��f#jȗ�t5�{HLrv2 8V����=L��p~>�XM���������I����{�'�ŷb���2̈S�ͥz�Ȝ����0-��bh�du�1w��R��}e�r�^�q�G�����A��1��s(�NO5˲������TM���ك} ~����E9���[��S�Y���&�˲~�ZNNֵ�)_N�&)f4�T��b��	�=�5�m��l��"8= /X �^��e-�Mէ��G
��nn�>��+�@��cƜ�v9��[<�*�J]�"����l���JJ�龄�U�_����G `9��-�	f{���p��+��Yɓ�K?b����S{2�B�>��3����ͱd9p~ABڿF6��!�+�P��AJ���,��^�21��TUF�~��VR�^>���?��*�uh����ߢS%` ����8Tqd8h��7y�2��D.p@R�9���_��4�*:�r�n VL
����Z��hS��'ѧ4���b�_�q+�|`SU�۔�n./{��K��vu��Z��jJ�.x��L4,Q�ж�1�$�D.~�+ ��>ѭe�U���_u��[s���N1y��'�<(�.��/6Z��TɌ(�~��+�x��nz�I�f�V�b�d,�Ć�Ɗ��R~�C�z������D� �s<FWN����V!�ߑ��F��w�6������}�R�[X2$�-�	������_m�Ι � g�پ>6�X;p��Wc)��c��ڤ��.���Z�0�շ�4��W��_�چ�֮�� %�G�Z;6���)&��N�k{O����]�H�_Z\�C|���:z�@5�)S�d�>(X���+�o��l����\��Ȳ�,vuIG�:�r�n:GR\��<?��\�V$��MX�fa�Akǅ{h��B��s=����B�Kt����uBj}.��شF�+�E��
mb�kw�B~������(��P5��~�1H����h���Y�I��75v�+�}��T����>=��n�,yհ�L��YI:Aa�s�2���=�	�����1�0��@�ۗ������E(�N�wx�ϚXt��h+�+��h�ࢆ[�d
~|?V�R�ߦH��V2�s#{���/��ᙽ���]Q���&���A���>@i��v	9[�+��bz�(C?��N�9۬1���!�+m�%NՊ��ݙB�W^=Kp8����>�v����$�]F�|;o��J�gl.*W�r�I?� 1t��|���'K �Z�C������S��������ܑ�>��<�J1�L~~1Z�l��*��������P��A�k��ؽ��p�">�T���\�K�J�p�O��)g��a_Oq	�m+L���j�q������=��*���?d���H!���l;'P�J���p�-��"Η�`��[^m�v�;�ޭE6l����E��f��nyH�y�=�9a�5�WK2��!A�����V�T��R�!#M��"w7GA�˱b��\�Ą�+�Y<��J�#�^�'Hy�����.a����ԗ�V�5c>�W9�s�{�F�Oh	~��35\�}�����j�kE��Z��M�X�88:�U����N����x�����n�&~��7ً-�+�����ҋ����]�;���
��"oͅ/ ��r�l��sNRi�6*��,Iǻ�yiL�h�&��ָpm�mk�YW��"H�Pa��� l5r���}p���˞.&e&wG
e��*�#��>5g,~v�p%��h�|�0�>�G���9�QQ�˵)�p�k+G�zMFp���6�/��A�0��4��H�̩�����o��嶪g���/��<��k�G��L��E9�*�U��'d
jC��L������a�Ro+�ǐ��@��lfd�����y��J;�[h�/�����-�`�i*�	��yUo慉��w;D��G�G��;��9YT�=\Xx�zӛ:��}�����EΈ�6����|�{]���'i}V�iA��_��@=�ïD��<�P�!�|r��5KC���6����)�\>S-ג
�r�>+cO3�4᜼4�g�%��e�:�]Oy��c�ϛy��H�B���X_�Ȝt�<B�j8~6z���d�g����];'���	.7�Y,�7t�l����ߋ}�U�c!����`�WZQ�~o�e7���нQ� ��'����Ą&G�_���D�:����~�qw�>��I�#$# ^���h �KB�!�3�Z��n�Y/A��w*F"x{��h���_�9�gL�|���M��<
{J����7����I���p���զ��Yq:$w��)���EL.@*��3,|��hQ�r�=V���c��C�j�����l/+����0k���eh$�5�+�}㪔�\K����[tE1cS�E���m�O�U��@w(.zj�/d� �N����0��\7��y�Z]x6������bm�܉�b3�.(��t�}	=B��w�ğ��HĺGH�r��Y`}{��A���'����ghr�i�����M���)�G��y¿^O=�*�MM|U�.��{�����1svX��aRc(X=�����o���(+�^w#e!��g�*��8�+7��'D������+�0	���j��п׿�l��IҘ��6�y�M�����k"0����~�%��#g�������2��9Or��2S��"l��`�wqh��M�p$�l�jQ�9�k�)yIV�Tx���y���@��Y.,!��?�������Б��J��f�.�"L9�"O��|���T�:[� ��O�����b�bz�_7ȋ��t[���:y�j|�GL�`L�|�@���?	.���{��9j����_d�j]�8��'0�ԗܽE�t�C��R˵rn�}�N~$�h"��p�0ڨ�����j2��c��'3ϯ=eCq��?�F���V2�܊�u���[v�Ow�*�/�^��Λ#0:�z|�騫�����p��@��$@�@
�����U���T�Ăt�\i��M�wD�9^w}U��N[�P���:��^�Le9y���;S=o���/K}�7�1ȁūj9��+
�Q50�ːe���Ȃ��p	Ok\���M���=��} ���i�	1�s��ԫ���l�f���S�iN'��q|�o�<@~n�c��Ppm6�(`MnY*�H�a�����O*ǒ�^�.3M����X<"��	 O	��dr~*ι>K����Y�#�xs��b3���V�c$��K���
�h:򝗙��4���QД�r�QD�_��:9�V����$�l�)@ӃiK����|⿭"�����fl�b|#�qa[��0%�_;�IL~�>V(�'�icκI����O*Q?��0_���Ҕ�����1=�G�-B����?N3���|���8�ץ�Z-���շ��֔�e�m��$C)��Y0@)5OY�sx��E�ВMV���gҷO���d�7Fi/��CU9W؀�_CG�t�2��k���7����k��p������C�}K�$L�LkVz����.�پڱN�d�+�6�_M2�ah�ߎT{�f]+�F�����cc<U_f�CV%��9hq��c02��?˩[�k)�?)k�Cp{]�����Ln�3AMVb�_���}{oIy5��A��8�3>׹ w�k1D&�!;�h������-*r�uN�3
��*�h6�_(�O2�a�.VK%�#��Et�H�F4px�"V���`�H@U���G#Nl{΅��k�7��Ub%U:i�rU�;�!_�ukG/9�CDc��f�Z���,��?��,�C�����&>~K0x��w��w|Y�3�Á�d= �T%�ފq�@������R�QC����Uw����g,���sj����� �59�#Ԇ�Vۡ����y>'$�a=�C�o�!W"�L���Ēm?�lY�ٍ&=��h�Z��Ȥ�V����.�� �.���ۡw�}M)�Bs`�y�F!��0P�X &+d���eBh���q~�/��ĸ�& `�jA{ʈk�&o�2��F[~z V���~5)�eر�"�^]���%��W
!��[|ǉS�����nx�q(x��#��J�W��p9��1V8�6u}��:�a���G{���sr��n�EAկ*�O&\J�B:/�������.��M�2�bװ�\{��{��8�"�IP-Ye;��@���� ��R?E1��ʑ�P�;eLS�<��ϳ�̔"���
8&>X��<�x���NЖ��=�����ۇL)��+��Q���1&�/t}]�E���n�x��F��K��w}}�8i�=_����W��:�@��o�1#�y/�I���Y+cӭN`�,k�+{���v�WU.����ԗ�	R��n�� 
��	��x��W. ���@4D�Fh�oa{�r�B����RM�!�a�Շ��x
�wEe��{�.+��N>R-��B�޿5F���0��L�ZE�K����>x�7Ȉ��-!)�_�I&r=�x���E0�]t��><���&�f�(�M�����ވ��H83�/N�y�mCw��.dsXm���AS�DmH����]Ո7�=��M�@B�]� �2%��dP�����OJ|ݜR��V}�3����ǜZP\�t���@gT�m.g{%��~�p$�wU�Z�0:��P鲉��b^fIf�>��w���t��+�Ӻ����r�ve
�p��)CR^[`d����M>�gF������U����#go��kA��pwUd/E��%�1�?��tu������g�l�c|$/	G�,��ƚ��hR�<.݅߀�Sn�~��k�T����R2#��w�� :�nU�q��A�Wp���2�r�`J�U��ǢUu�Co�Āj+d�F������Z�us�^_�5f4{$u�0[ޤ��2d����jSПY���P�E�d��$�V�Y3{���5�{��H��g,;H ?�栬��+�9r�&�sL1 �ԏ����+Ѭ�N\��J��u
ϟ{kf�9S)�}OX�A��/��t��`r������7��{�r���c?�9��Yp�b��U�~�:gzZ(�{��Կ���{Op�?Dt�����r�޿3��2"!�!����/xY���z�%��F����a�����3j���/���H����c���! +k��T��%	�؏�d�N�Wᕣ�W���0UJ����p���}pjJ$� fz.�b��,I-ݻ#(	����@pI���L�鵈��Ҩ�2�@�g�����˖�5Ҙ��j6��h���YH<�v�O��v�Z��;�b��{��>\�U�+,R����R�����̰��p-v �2��2e����k(�:{���va�V��*���g�h�t���#_M��Q`��H{�?�K��
��n�FB�i�؉���2��y)Q
��G���shqK@��wI3��ک}��!B��rk�cs`��y�zu(+fے>'0>�,o��p�V4�t6����>[�� Y�O�r`�a~|0�?���P�!K��R�ٹ9�a���h&�|c��.�mi ��>��1�Ymis�L������86����ZkBV`φ�8luń�#��jz��o��QQ���F���g'^��꡽�xRޫ H���l�^ԅ[�0,�����5�^����-�l!2/s{�؈�E)riP)!�<�Fh�w��3�~�p2�}��7�ƽ�O�_�f��}��z�����^�.��:eS6ɾ���V�u��)S��X���ӹ�`L���cd�m�����+߮V�V�VR�J����g�K��~�Ӫ��.�Lĕ���db��TjX�	,2G	=���S�Ǫ���b�F=A��tU?-[�o�3�{$b�pC�f���p�����~�#S�ӋA|
Ɗ$��y'g����ꐖl���<�m!�������@������"�Ю��-��z��-_�,�?��aS�����|�_�����8fK?��DMǷE�Y�6�K	y��խ���x�$�X/�������*<Y���*0����	�͏�7n�]��X�j���s��o~���jM<�S[0�Olj�o���Hф��mi����mT~q��&Q��	C���~Y�቞�]q�-^�[mo���-����)S�rϜ��X��pG����P�b+�l��Hٞ!��a��U��3���%��������(��1$}�*u���9����s�#�ژo�Q�c:M�+�Ɗ_;�b�Z�������F������|�b _���v�A��T%�9,��ng���0h�ެ��V�w�O�wJ���2�A5�p�K�s����p�cY���=�[��wJn�Q�H7���`��x�)/9��c�Y!�I'흙c��mz>R|��8#�<�����Ig'�P��i}t�ǝj�>?{��^��ֻ/�@�1�)�l����njq�f�Wj���x?�7��� �Y��|�6T�
lH�
XJ��4���?Ա�A'��P~Iv�/�D1�m���' f ��m�)or ҎD�%|�u&~�1Uv� 6�&f}���EoZ��_�a@<j�lɾM���ww��$��rp	�Go��o(es
�_�3p�@��XG8��l��<jn�V�FtO$�I�9���R��%J������_�aEXCb��]�LY���"Mn
�����)��x�M�ځ�7�@8�u�(��ט�W`1'*S9�/^�Xl�R��=%K6�wh�0#D�h&���N���U̯e���2�����
�[�����(!��"�8x]W}K��� vҩ��'w��a�6�<u���p@��?@���Ù���9�o�\_�[��i:��Ć]� �+�1��8]3d�f)^��c)fXX%��a&�������wj�0.<�0�r���1l��5�*y��ě�ڽ�lU�	<	�gp�-7k��k�4؁�O�w��&��h�}�5/]���_�}�^:������i��l"��,��rT՞ZH�?�;s���o���U��1�=x�yq_�V��e�<��F������a�o�3$�ȹĀ{���5�t�s�ӉN� 2ۅ���ے� �ڬ�B{�zퟲQV��^�E��^�1���R[*��m\�5I���a�N�6�v�c��+2MWv@P)O51��)T�܋�)�g��`8�S�#�i�RT�k]5��;�2!�����>��f��d�������Fe2�F���B���SE����+P=#'t���Z�1eO&,=���fj�HD���%�Y�xx/+X����#������PK-�o�m��#<Q�`�a�T(�g/'��D�Ү^?ݲ��pY���pO��������CY"l�;w��l��#k�"��?����c����+�HJXt�i׬�L���r�FC���d��������S�d!(e�FWF<R���g)�q��-������9�:m�:�[l��Q��%  4Y�6�*��F���)��"!��d��^�)  Sjf����W����n��J�z�BS�:D%��k&K"�B��w���ϋw��;?�5��w�X T��[,�ZnPT�bO��j���1硖H�MB��߉�ZY��L;� ΡE{l��	�ٔ�F�ҍ@�<�Q��*i���mzt������ӗ�|���mި�׬ۄe}9�\��q^��#@rs�$�c��3b6��C �%�,��̠y:�0)�Tͅ��Y�n���ƞeW"��E�sT<?���+�b�c0��S�zY�6"���S������dqo�hdd���TLE�B7:�yt��}�����3d/)s7�`�a}d͖:�'9=0zea(j�{/+�{i�wekn9��>��	�P��z!�G�������x��������$�{8����%5
��j�p�d���-��(����Wu�LޅU�Z;q�G��y��S��e��a��r�ި��(���v��SP8�a��r0��=Q<�4\�LS��,�n���_�L{�k��Gݦ(�B��H ΄[Ә����{tO#>U��1s=�4R�ߢڙA?���Qf�J�Jt}B��S���ԊY�=F5r��~-�h\�B2a�۔:�V|sOW��u=��9����N��{I�R-�cJ� 8CJK�����#��`��!��$̜��$�s�L����V����0GUo���F	L�C���e^ށ.g 
��,��{���t�*��QWg�H}E�l������Pw��p��"|>�g�@�+Y���	4�]��~�e̐ɍ �-йD00��=�������c�_����s\�4n���j�`K����U#F�"�R�Ao��j�M�	�q�G��uIQ�@�Hw���l�v:k;�PJ[�b�u���l������P��2�L
�9�B�4Jr�k��Pir�ز��)B��i�Z6_����-$I="�T�.�*�o����E��-���t<6he�+�~�{�Aȯ|E
�e5�]�I�8E��c�hݷ�V�����=.��W	 �vW��H��N�Tv�y>�}�v^38��2lT�Q���1x�z�n��u[���`^-�c^Hv<�oe5��%Ⱦ�?{�B�5����p��S��dբf��Ξ�$\��7B]�~�ݙ�"H`t�(ƚe2w<����n��?D�Fnt����H7�Rp!�~�>sgv0�^,Ѻ�����LF�Gē l����nΏ�v��� ?�)K�H����Ѱ,S�W�8�V�]8p@�)�;oi��Z���1��i_�-���z�@���� >��rB�sޡꊾ��{��i��Uz���וc�Ĺ�c�.�����g^%�6���$��N)���3�V����eV�m��{��WKM=8�w�s����boX�J�l�oZ$��b;�i1�(��з1�mN�� O*b,�3=�f�ŵ\��6�~mDvSxP��pv;UD����tL
��o�/(���ӸC�ep�!x���&�ړ��)��c-����;�����uW�G����oi�nQ��Ŕ����C�u�켲�3�F��A'�ΕUY�Z���'��4���e��~���Ra�������6�.��0�jث��jN\'+(�!܏L#���?�n9��C���>15d��˓�>��k����NN*>��Ｖ*���Bx��� �z}Q��C��Kf�f�zTC��u00�U˄�����r�������<-�F���d«=$k�j�"*��(;7�|f�IN��;,	�r�u2K����Y[�;��;�������.HVy��Y 	v)�A�����H9�f��F#�S%<>YG���
�hfsSg7�y(�hj7��u�;WBf@��}��UE���:��u&=�0�_[E׊��=��gE�s��	$␏�Q7�me5�^�q��~w+�����'ˆ���|5�԰�b��Q=Z�Ϣ'd��"`����?&��{{up1�ɾ���7��N}�a,�c���a
:�odFdO�2� e��D��9�k|Vj� p�WApoE���F\3�H*��+��)��k�C�AHM�<��!m��Y$yZ�9��I�Q+�<��-8mJ�|��m�������� ��b��4NSb��Q���r&K,�^��J�'�*L���5��*�\U?��8z���2Kq�h
͜��FkrY>B�D=��*@�5��H��S�Tb���� ��
*�1-�KO�2,}��~ ,5�R`_��U��\�K�-tha��j�sP���lH��P���v����Ж�V7qL y{!LQX�H�ʫU}����kè�y�~��۫ �DtCar���#��Pr�S�Uv!��W���v��D�-
��	aQ��ֱ��c�E��C�z`�8ڃĐ�}�ؾ˪<J�[*E��2j��%�/�CN[�1���LkcT�I�8��E/��������Ʃݯ�o,��V��_L}?�xV"�����S�3:����.�UӾ�A�O>�D��4WXÎmuD'���)�ь�[H�����E��&�n�̊�����`)4�!�Ϭ����[�h0�%��3tlu��<�����}"|��QV&��
T�n��dgD	8~�Ol]���o�X8�t���$yG�~�c,�,�
�����i�6��%��->�w�n=���$�\��ֱ%��e�$�����s?��;�3Ss�S�?W�;�\Y",�6�������hB�2vL�j��R~���`�>��	-/M�q,â)����SД��������A��B����vj��
���d���xMԡ;�E�9EM�*�X�f���{�-E�of���Y�}�.jkE�7o3�߆F֔�k�]<���鍾Sz�[��;}�U�/��AlF�L�HOԞS�pr�|����.u���{����t*_���C�\I�D ��qR�3tZ��C�Da��_gȓ�++|2n��IѰ���/24|�����s��9g�q��[��M����m�m��gGw���;���rfz����f�^@iz"Ɔ�%)�K�q��F9����2*�������,#����-��42rI��5u���evpm�X��Qu����� ��6N���N'�Bר��!4�ņ�A��,�ҟ,_�2NI�DCT��Ϛ�&���%Ef�̥��ip2Z:����L8�!˩���q���n6�̮ݭ��u�$���2x����Q/���e�/�41ɯ���OiF�[��	�w!�
h���%��K������f� ����(o>%g��6�|�Ti��(
G�a�`�|wF!s�
бs�����L���ľ�X��� hE��������Ǟ����]��q�U�y3dv
(���bJ�[:����~�]LJo�QI|�c!]ݿ�/Y���a�b�"�Y�?��:�~�}�x;��t�%n}� ؆��E�&Oc�gE��_T-
*�F��F�h����8�����c��X8H8#��T7��   m����ا���5��G>k�=�[+!o��ѭ�}����m�.x��DX��-̄K<������h����Ia���[�QT,(�[�l��#VK♭.���"P�>+~���UNd�ﰣ�������	���S�LX��]��kTCt8W�Iۖ'0��ڲ;��2L�c��0���]wm��Go���9�A��|�i�����-;;"��<�n��9 yEN|h��t��q�¾�ظ$f�yV�yKX����B���;�c�4tA1?�~ �m�!A�>ÖG�u�6��K�7��Y��%/�6o��!�q���Ǝo��q=�[���s��A>��x�[J�S�@]���"�k�����U����H>�O1�OU��,��>�>ݪl�/�H;�	C�>	����>e:����;�tą��t53��wb�VV	�MϷ���e*=6p���X�<)
,cB�������/z��$�r#��Γ�L�����჉נ����3`���r�`�iH��?�������
��O���s���m��Ł���'�DL�b&�:z	&y� d���X�y?�N!���ޒ
�`��½^��Np^��ҹ���ڻP&U�h�!�H��R��~�f����UҬ�1*ɼWTقy�E��ĸR��v�J�l�9P[��$��Z�����&Sh�k�[J���-tG��yg�݂�����?�]M��;P��Br�Ҭ�Qi��y`w�
y�];@�)aU_� J�б���2��(�'7�a�<����>�to\�Œ�C��S��wH�S(�&�:����C�!��+�z�J��ỵ�n�>�qڭ��gH�;�`�z���R���� sl�O��Gj���n����- �Y�T��{�+c���j�韫���������"�L����\~�^��'��Կ�q�1i=�>@�͞�λ�﷦����$&NN��c��dx���x�����>=�t�a0����{*P���4.]���e���)N߳s�'�Xn��y0?��˥>�U�x��z�p"�D�u� ^�~e]��!rD���%�b,��_ke�W�7�	%�s7�G�z�����<�A.�x��J3I�M�.m��x{s+]��6>~��61L,e�����ah9@KH�D�����Se˶�`=^��M�H3
�o��"WLi��q��� ��U��[	��5k��mx�A�U 9��k��;X�&�W>c/4d.�?�4�`��0Ԋ��-Վ�dؿ��/��W&\�b�J�z7���?�mF�!P��@�	pd����?�D43Jp��Q屠_��y%Gx�48C��SvZ߬�Y%l]���ŗ84�#��+e�k��/��������z�p˔��(j%z�y��0.J�J�m�����#`3�{{�bc�#�މ���<�Z-�Cά�
�t	(G�y܂������{�
�;�0��'3�d�rT��ޘ�@�~U��<�_di��8LMhz���N_�ޜ�ʁo"�rM����X����B�2=W\Z��y�z;�āy_�!��ȗ���f�� �s��!�5|C`�O���-�"��A
5
�|�A��n�����?;&�!0Sn�0h��2M��1*�p�`���R�z[c���"B��:�l( ,t���1ni�~�Ռ2�|��kO[F�ؔj��Y�=�Vt��d�Hc 4`G�Z�T�t�Rݠ�c>[|7;���T2����3��.F�	��%��q ��+������G��MT?UF0�~����C��RK
<��:�L�+����������i�0i6��g�k*;�EU�P���*��Ձ=��Y��hġ�+�Q��W%�:#��&q��*ܱJ_��_�N�ᇢ�n1U���	�-/�ꞩ3�\&�R�m{Ʌ{ͳa\lH��$:��/cel��~�W�XƆ���s4��Y_-̇Yw�ᡐw��G��&��b��������3�2�^�9���𞁚����a�`���P��8�0�����k�P���~⤱t��F ����o��; ����#�dD?Iٴ����u�f�B}��?,�բ)�ئ����P35ޡT\�`~���D֌wN�����c��ƴ��\�y�d���ܝ���?<4KHn��?�Ml�Y�����2cOmT��V%��l� �z��)�<ώ�%�D���#+��;��a�,�Qߒp	h�S���g�KYK����!&8��F\�2-f�=�B~^)Gu�p8����7�2�ݷ�d\k:D����0UN�D��-�)poE����j�/W�7b�Y�U'�X�l�İ�P��_~��ݖ��q5ȅk�t��_��9,�*ɗ�s�kN�3��B-�0�������W��j�[��g V�ˆV#�����g��3Uؑ��#GL��IH%�Ef��?s�����ch�k�Ÿ		`��͡u���ZN�-	/n����Q��1����\��E�.B	m�����9B�ː��OѺ�΢�^ߤ��������u�H��N&��O���"�X��t� j+i��CsOޢ�nW`l��{�uf�oJ. �Ѥ�:N���R��&��ڻ�X�7�hۙ�рn�6���g�0f�cHg�7X-��YH���ұ\�^/w7H6�-��+�0=�ﯦ�m�;
<X�_@M[<�z�r�"�;o0\l`)4��Q��]����&v*�(G���N�$D�U&`W<�Eu._R>��MQ{z�8��>ܝ�Cܐ}Y��Ef�P�s�9\���tbB�����f��ڒ��[U�Z�mt�VHm3��ǣ�:�N6�42�`k��&ž�H�*�?��H|��U<�:tV�d�4�$t�8�S`���_ĘB\����S ۋ~�_.u�;�λ}׭r��Hɳ�k��VP/�n��b���O�˕4q!J��q�za�Zx�;	ug�2v�h�����'(����d����4$��E�u�/��c(,��h�b�]��doͰ��aH�&[H0u��G%�8:��)���߭�A�L[�r[�j�xr�L�K�mB	��l}Ǝ��0,�����c��Y�������İ�l�QGyJ<�ґo�d\������7g��۸�	;)���/7j�9��MɌK��_�e���	��Ou�h�д�{5I��(�S�ͱ��l����
��oAJ���k�-�+>g�G��.���9�;=���y�4���,ݯ�	Bӯ\��X�.��q��O�w�V �9�mB�,�h��wrM(A��B��l�tW6Y�ޜ.Nu��ʁ��.�/������^ۭo���:��;��&$x?�HϠZ���Rf��k�4����7���q��@c��y�Vf>���r�D�+(8���>}��F��.��|�S�����'a��8�q�1D�i�������Q����`f�91t��O:�Wݙ�y�g!!����7K(�A1���/=@(����qE��co"�[a@�gz�t��k��}��Ԫf '�ۋ�F��E[`5�A�v�5q	~^���Q�*���k��	�Ψ�v��b�����ވ��0����֌�{����_�.%�DK�_�8���I�' ���#Q��)\(�f�>���X7.��I�,=��8�g�af��^����x5|F��)/��	f�^�^zw���<�0p��,Қ1qtڣBĀD�<����uv!���2�8���z�^(�[r�h,?.8s�o��xѓC����C�-��2�5Qξ�Q�Z`��F�:X�;k��Q�*	�{!;�,�n�l��X��\ �]��(�O�B]gc�?������<q�����>�C_�}���9L�ރ���ɧ�[����J?��ݸ���m�#Nz����
�cc{�ԕy�WYǕ���ʲ=�-���Y�*�V�����YQ���<�:�KLVHki.h��<�K�J��������S�yyj�%����y�c�����&��o�<�(��D��PX!.d�6��y�yb�]�Fr�}��X[��Q�B7:irVZ��F�Ƴ���Q��v4�>��5��/]�2mJL�9�g4{h�d�4�9Tt��^��H8��)u���M@�ہ=�4E�ޜ_^.�~m��$V ,A -�h �L�O�1��o�5����?ۆI�>�%ZAh�k�#��~p/3h�2_�$ԍ����v��PQ�r�q������f��B�(�\���.l��i��Î���0����H��7�|۬��e*�Ҟ�L4��;��`L���a�e�L���O�{��2�M���[Ǖ*@���V2�e��Dŀ���F�By�Ee4r*#��Ͻ�$4k���{�[��J;5��ٮ��]�_{Y�8hU�}Iz�J��z�]��x��s�P��&&fL5Yv,1a���<ld=\%V���� �;����m<Y%o�Z���9����y�;��3�5�'�H�/:���~�./�tm�Μ��� �z�/�ֲ^��?:��Ȓ�s��7�2֚��v"Ԃ���ݗާDN��u����gQ�����8SV�6��	a�6PχJ�3N����w�.e�=�0�=O'S�aw�.ѡ�I�\X���h@�D�F�Z���E�*��IpI�(��k8Ӏ������>�1L�rˋ\nX��?o3����`����@��H�J� �+J�
�7 �ǵI�q�Ĩ,,��9v��"Fej��%n���=��:'�j�ݬB#-������A͆��K~f��]�����&�/�!=1�8>b�7<�"�F�ު��F��at��d�'XSms������dm<���%� �ɿ�U:Z����x�p�z3|
�4�^#��X����'��$���@<�ܙ����b w�2�;���I08� S0�w]�V]AP��zؤos�'~�Ǌ�b%�O~9#v�{*�Ahɿ��dA�<�Iy�Q��1��\��u��0�	�����4���t�����
�p���;uB}�po#��3̓�}$RpO�iw�BU֥!�Q;~R )�',i]]Ϝ��7G��]�;���0�[$�mǎ���tH29jWr2F�tx��.�y��Վ�$��Z��]z3����m8�bn�ث�߃�����Jk�PJ	9� )�&���ȍ?cJ]e%�@q|6��!��������/�^+U6r��ʕ+(�����"Ocpd��L��Q����@ �(��i�BŮ(�l4e�����H�\ࡇ��-���6��h=����}�T�_�#�I�ʃǁC������!�a��#KF�L$L���u�M���Ny�S��2���.������E�'Qf~^��퉀�1��$��dWh����g���F�΄�Q���y� H�]�+��Ю=����#̹��)|��^5B�ۆg��e:}ݨ,9�d
\�"ww�!�32%��T��$,�+�U
������D$�)� ��y�qo(?�� d]&�N�T�`Е��=��D������W���L�(L�I�����Q�#`�q�J�:Ҽ��r��q��	�!�(T�E��j#e�� ���)1=L}\��d�A�'qa1cx؟��(��s��2:��+�]:߅�/�Km�ϸ%�3 �*\�7# 2%Xʫ�{�}�;��fϢ}<�_��*�b��m��z�:��/;����m���T��"l�6���LՉAw�� �jPV�6���~G%�+ȥ�2���H���L�����C��xC{�7��x�B�����xv$�U���ԱSf�3��oa0���h��X�u�rr§�6�i�amH���C�a���Zف�+�*��������,��1���f�1zk�3�$�>%i�����x�\dJ�h��dԞ8y�Y�{5��ˠ�'��k�I;�XBk,�L��g\P$��^fM��.qk�ΞuU�wW��:t�>CYQ��i�!i1�B���%8���%�j�"�Uتb�7v{���k�ق��A6�A+6b���X��@}�6r`1��ķ�r�˺0��� (+�@�"�<p��=�j��dBH曆��g���;18"u6uЙm�#��r���B��*�<݄��b����JA=���#�́zi0��i"i���L�~�)7��쇀�$�>�Ӫ?ߘM��/�v^!��<�4d FS?��M(W�/�^�78R���$X��O2��t@�-
j�}0놰�X!e#���Z)۲�0:5���
mӻ�=����^��:�H,���5O(�ݺ>� �3O,�jC=���1�HA�4� ?��� ir�J��QH�9��x�!���B>���&H�+C�kB1�fP;&sV�:ܶ�4���)���$aȍˑ6�6��f`|ԙZ�#���`�H`}�P|ZS��p�[�v+�A�������#���;��kjcfv�K�
��9��4̤��M9;���)Q��\�vT*K���a?2\s#�Ø6��F��R(���F��X1wT�zv��X��BM��^������S�̆�ò�r�����E��1u,,w+�I9E�*�UR�y,P��7'��hz%T\�UQC�T(�ٺU9D ��:��x�~#�n:Z�*�ak�4.�;����e)�<+��	�hnw��A�V�0E�n�O�8
�q�U���~��d���P�8��*m��z��|~[f�q��rP˖�	ѭ*%�4� 5C�<8iJ����&L���"��ƃ��l��1�j��d &L���s$=[F�T��#E@��5f��?�]$�)$��5	��O��\�X��|�;n��0y�^��S[������RUĴ*��z�9��S�M��fǆN�n�B�Ȉw8�v�[	���y������y��cW��Hu4��R��S�kg��k	���xh˦,O�!�?��A��e7ȓ� �8W�J*��`Zy����qc��3oc�I�~j��}_.82��V]�)���By��'O��B�>M��k͇��F��'���V�n�dCM�L�:�:3n���@4q2g�����W�i)\�+v�?�mDx�� 8�	\8OS�w�[�a5C��p=� �/��;��q�^~#8F_9ㅣ�Mt�s0�*PnH�d���T�m�!(]�O`�+�>p�����7�f<���S0�31U�H�U(�8�`��gr��,��'7Uz�/��#��8��c�t�!�����8)��~ty����xު��CN�.��g���Q�LfH����Kn1�'ó[OY����Z���>D��S{��d��,EQ���0�br�3.w�a�z�|Ea��5|	Pe��yz-;P�P��ih7��R�����g�uh>t�������W��;*��Ty.��e���n��O�e�^L<*�tWG������T�k�b�{�Fs��ŲI��=�o�X%�����]�}�S��=|����Ȁ�A��9��%t�_6�����#�5t��Ǘ�^za�}��B�7���=�8�>�e!��8c!\���#%�C��x���q�qDa�!�p>@��<�h��r/z�ee���3_\
�ST�v��g���Rz����Qi��������,Y�X&�����Q���]^��J�h������!$��%��T��=P6</�2,�Ɲ�~<yna�Mv@��g�.�7�ܠb�IΓ+x�%���|T�:�*6ԖѢ��
)�2M�D�?{�v�Z�&��>����d���7�m�guC����M��:+9a���'���(9��_xm���4�ܺ�,��U�7�Rو7�0x�o��3��XC�
���L�
��H$W�F���`�RX��r#�m<ҋdѩ����aq�+��o͕&�5�vG��T��D�C.QN좞D���4�������F⤜%0"��,OH}��[8�P���r�:5����v��w� �$"
�$oO������1/�X�^�("�Vr�rk���Y^&�퓻t�� ��{R��-�΍`�ϲc*ʟ�wߒ�.��::�ٛ�{}��	�fޑA�����������q�`#�T�iO�Tq�A{�-L�f*��@ǎC���޸���ʅ��߿��j���&']�e^�fr��5���ܖu�0�hvǩ�k�rw�I�s
¾�]7­�Q�H�FS���������m��+)�Qf��}�O�e�s��g;v���|[P& �v�ڔ�vŰ����y��wh3�V�Tv޺)kt����69�)�(=�Q��~�$�:��~r�]�.P����+R5�C�vRf^,J�#+����Xc�@u'=�nL|���Q��&v��`��-Qp���F��1����S��0���$�oU��6�N�9�_�`��nY�?e}�+����0�ǘH<�9�1P0��A×?�ui��\e��/U~RV6��I�����+(��ym!6�%�f%4���O��e��(��I��)�F���v6GEia�w����� Q5��^-18��L$�=M�K${��q�9SyhymܨD6�� &0o���]4���j�wl|��$si�G��R��D|�T�|R����s: h^­0;�љ�r�M�հ�Ė=��D��x�4�6��BfFh؎u�c�ʨ�k��@����_�p̾��"t|9�`"/���;��-йc�FNt��}M1>�@'�l�P��j���^�a¥�!��DފT6,�!�m��C��;����#�ٌ��5S��5�
a����9|R��Pscq� ��ݦ��2�6��|�����IY�,��d�ႆ�����a��9�B�֓i�����	j�+|~�*G{�S��i�D��r����*�5V	k���z����\�u.�t�F���xB�
����b
[ڣ�&H�`$���s��<h3��B��^@
�._A1�U�M'8�(y�95�969�N���v �3�����Sxl���j��-'�S�o�T�.����o�����;��ZE����trm��G�*�������JKpVu6�u����Q$wݱ �mG�8!D���ה�6��������x�l�+Zt8�0�/��}Bsw�F�f�b�;��q�5n�#%B�е��AD��D�X�7.�V�j��c�ヌ����}�e%�]�8����2[=�*h�cm�:cŋ�]�����հ�'����Ύ��%�OV�Kё�6v7�\�|��5z�ƚ��p���s��=9)�|���3�W�¯���2��B�z7�3�g���f����ܠD֢4��CŅ>2�����f���6�;�v��(9ZѰ����S���|a���+�N!�J���^A<bw&����p�~�Nb
:��p��>�~��;���(��r�c�;�-�T�9mI"}�l���`�b���>�C�}D�f�u�Ͻ#O6,�=O�M�
�ql�"��{���o�a��Ta'3W&p����2�ѥ���9Cn���i�bո15��̒G�b�`ˤ��g�Ǽ3�G�CW�A!Y[��S����
2j����YqIhİNt�~�"F5��X%^�a�O���A���i� ���-�ܕ.���g>�k��˗��oX�:��G5�Vc�T@g.����CI����?q���Ĭz,i�m�\n �s����"k��iG.���@�p�|�	�F>�f�iT�5�	���.��~�ϧA����s���Bx�]W�|X��&�x�p']��:�s, ���<Iߒ� ٯ�&�x��e�@��~��� 	wc�m����'L�尌�g�Q��7 9�A0����/K8�p��FÑ�b��4������s�9;�%(eyq�gȶ,.统4"��
e��~X[��l2~f�ixx�R�,>�G�"'l���!�窌����R;Ldq���.�rIg�s,�8�|'"b��Kf� ���J���r���LK��s����ݐuT9�E�V�ig	pm�g<�#�o&¬ijѳ��o%ި<];�}7�FK�����߽w�J�;:"�����W�ok䶚1�:�+��4��^A���W�gtF��튡�c������]�d.p'�G�ɡ^ۓ���U递Σ��Qhx�ӠY�6����	�i'0��WJ��	&����!%�V���tQ[�[�h#g��DsX��쀐^��n���}Q$f�L~ .�1�p�{S���<���ⵃB���yƉ���)�m�#�9 �9�mp��0Eǿ~ɒBB����6z�٥vY�Jy@��HCE-�ƫVA��CJF@���^`B뒶�Lrb�_ �޳N�P����)�X)O
珒��R�S��e���H�����&��&����&w^���j/\a��5�����|��S8� �u3�+ŝ�c[�/���������4���k�
D����lS,�H�Ƥ�ћ=�p�8���I2�g�g��۠4����f��'+�Jʍz��@�S���e��=)��ERJ~���QE"�q_p� �R5�X��$=�j�WOM�o�S�E�@��V�^f��iV��/���+Z0i�,�i]68�ɀj*��rK�t�Q�y?F�1{�s���2RDņ	e9��`��;^E��Q�,�P��
��}p,��,c��9���|�)�DǺ���ѡHπ��L:��ey�$�)�}����<\J9	9�U�ޚ`3�L͒=�����R��z��'�"*^��	~I���Qj5�:�����n�,=��sz�sG��S#8[>֏����	��CΙ�&���	��;L�]�����O���^��g;34�O|�b,s��/x�������`�\�&8_�,&ey��]VՒ�֊aލ��p1���VA֨���r�('J�o4�2���Re�g��[S)E�o���'Ud�eR�'���(����ٳJ��zga�j���gLՌ�V ��V���kmu��KO�^�bJY��eQN��.4�kޭ$���o��vX�.3��ԣ����db��S�|��""�_����A�X�
��.[��f�yH�B��F�O��A|�u4��i,Z�P08�L�n��9��=����46���`��U����9�8���Kʄ�f�ţ)��� i4��<��sMĺ�U��P���V/c'r��5�p�|Y;�Avo��bx4��I^H78-,��}�|P�X�r��%?3[�1����H#�G�)���i�&�����k���`���e���v��.��RR�(��$;�(�ψe��̲����K7�]�p��x��M�
a����X,P�)�Tn뼋�$��7M��U�a<X7mS��l����U�'e��TPT�"�YB�����IO��f����'W��`K{b0w7s>%5�����#�-�ٝ��Am�����-q��'`�������gW� &��j��E岮�����ٰ?UHA� tb�u
L�6|�q�yNi�lfb�O1"r̛�Qtp�Ց5��jN�)Ļ�iL�>*���F�;���n�Z��%���D��h%b倇�+�q�Lݒ䙸�~Bݔ�[$ 6(�K(�k�sb!�O�`�\��P�^_l[���w�m�ԣj��)�0q<�XҜD�cB��h�L�>��#k��2 �y�{�Z�yg��ٳ'���X?-��1fǒ��^����`�+]�,���+ W,�N���D�6->����F;�K�ϳ47��X
L�K8��{{h�CV7؝ȓ��YUͪ��Bs�ϝ#��7�Z`��FsPkI�?=�]�^�n�zn���4bp�BDW'�/��Q���C�M�R�N��5�L�PO�y���xe�<�Z����l ��.����e�H봯8��/뚆H��ɔؖo�����s���Uw�xc��	�n�ЙӰ+&�����o�kߪ	� ɣz�q���FdaSS��7�b�rW_ϓ�Y��	��_WÖ'ǅ𥵞!&����H�͂5��8�TVrKd{8.ږ�0����{x\hf0��B;=��C]]�2x�6��"s���N"��;hx�G����'廊�|������$I�re�;�DR5��,ΐ�X�$��[)�
9�	d��MSu&�q��>���ژ��&�<yXD�iS�Xba��nR�֬�5����Pn�7H��!*ϸ�hqE���"Sp&�`�D�{��_���	���;�&���gH�k�2�Ò�6	%|��Sb8�y����{�zĪ�Ҍ�7'�2�A,����s~Ɂ}�q��_$L��26#U�)J߄�O�aˋo7f$�u^��k.��):?^rx����0���:ϱ��?�ya9~F��F�,��!f�`l�çT��q���]Sԙ��#���q�mH�R�O�C�a� ��.��E9��qc�J��q%݉�n�=�#� ��t���$��a��7X�Q�37m(bmΟ����CJ��������f�Q�����;c�e�j�A��$�2�� �7����"%:��.�p�W15�/֋�y�8�	���b;�|��Ɓi�o��B�z�_���&M
y�'�b���JU6H)�%=RA��#W:F"泜�mTv��
X�A��@�_�}9���N:��p�'�\x�s��!5o����Բ�'Yާ���p���SNzת�7f���#�J��<{&���������l��j�($Q��R0�S-������Mzԧ��  '&N��C�t�B�m�-���.�s��RCup�/:�݉����c`_J�"ܠ6��b�[>�Af���a2.�$�\
��#b�4�Hs���+ ��H�"I躜Q�L5���~\�?�,�%`ā�R������9M�K����#��^J$�&D�L#!����g��d��(��vo꟎7`�K���d���g����Y�n7���s�i:�Ͻ`��Re� Ĥk����@��Z ʄ`K0Wu|��tO����t��G��p�����I�{y�j=�h]�m��+�*����*Z;=��0���Lw/��ps�t�4ꗾ(�~��u���~|q��8�N���^�y�6�-�\���9�ңT)�pR�߱�%ARP����#Gq-�E���[6D�D��8VrI�t�8��VJR�c�W���d�{�L�-Et��Htc��r\j��������<��T�>Z ?)r`��6��<�8[R�;\k
���N�/O}e@�m�PI�E~F�	���oBz�J��3Ij��0`���Ӑތ�s.�C~�%{ґ���3���_���4:LQ�0c
C(��^R�A�NL)C�]��-F��߻2-ױ�}��YA>X	ڡɕiܯN����i9Fc���d�Ԧ��ա��-���:�Řbzy��:�ι*�{1��C�qOQ5PD1IJ I���ڶ�8�?�Pb�J�c���z���D%��\t��������@��`;U�������iЫӿl���6�oxL�}���;J�_/]�)��B=��?"-���?�:9�OΑm�{oO	���oZւZ����}�H!
N>=���%Z���[s��8�����I?Bؙ6�v����\y���`X�B?�v�[{x๙���j�o��Ѳ�����PDr|���S[óq<�����S�&<�3�����%�r�B�=��RPCǃ)�T��~V�w/��1�/��G���Xa#��#��O�h��:J\�H�jǸ��Jh�����M~�"#��Ɵg��XW�ⳗMp�n��}�gq��㿖5�P�_���\TB(>�o	�y���4��Z�7�֋�6���"΅w�.$t�v��O#j��E&��"��dY#�����I2�`o��a
���iz)�q�ć�O���~��+���$��zʥ�ٱ#�QK��,�t�塾����`�c<�hD~H�I�M������A���^���(@�E77�_�.C�e�6ZXB{�K˲JW]Z'Red��É�@�<��j_��;�=�M}�nr��o,�=Hp��YR)D���v�AIj��q������v��>s~$���V�� H=��0�"��
CW_b����2��2az�&�����rn�����SlsM��,�����JU�U�6�?�H�BpL� ]b,�~���qߋW{�r���D|�QkjE�Qݝc�Λ���)�����DJ�M�V; �B�ǲ��61�Æ$*4�bj��R���\�K�k5,]��}���b���F�p���5�Bā+���(Y�av�C^�X'O?��"�Yt����i�w������L�?VM����daBǹߴ}�u�6�#K�	�sτB��G��Yx�84>͊G��&%���o"���y�/��"b���u;����G߹�m��5���&��YWW����m�γ�j[��^��ǈ iG�-:j��Ͻ�m�|I %���Z�����RW�d��#�H�DT���R2�M=[��Ļ��产�L�=�/���i���(Dz�_��o�;hő�� VM,���=",T:��6�:r��w��Q�sGS�Lm�Ko�%$�]�����}�3�Jds�_n�w�ƈZ��zw/Cѭ7K�����hP{�]q�y���J�z��XΑS�@��Lg�#>�f��6%�_��"x=:b9�k'I��磌�"����]��:f�ќi
�Rd�v?/ȡl�����͖o���NA{���4eN���)��,�w��)�0��ܮ��}��V�rz����.@j���|r?���k��ߵ%Ƨ/�ҚgE�+S_�~�eZ�O�@,Q��L����%[�5���H��j�
@W�*��u�1VR�&�+���F���I����s��uV<5w��_<�f�DɒO�'E*�����
��4]�\�̪����m��ܑ>�r*KD���ČQ"{�_�F���a�f+W.��Dq�p����>�T ��n՟3�6�I���ȀY ᡓ��%���RT�%�N=W�z,ǭ��=����=�o�j�bKq�Q-��s�8��=�K~4VJ_�۟����*e�� ���z6�$�MM�Mh	}�Ho3�Ky&9�<�OJ�/���]���4W��kp%�q������=WM?�$�fgUG�Dϝ�_�[����z�F��EW6�1��OV��N��-|�ٽ^F:E�Ր(BH�?�N
�/r����
3Lѓ0�����lMf�� ��0ARګ.�yt�8ѹ��0)�r�&���[�4׫l��L��E���-�i3��Àl$hPZ'���1
�+���#@uU�T�p�/k�����_�#Q������v�{�Y��I��D�� ����gI�Z�5�Gń����S���7�G�0�}����`%3�øy�X~.zF�Drf,�E	�>#s�}YN_���cH�QP����y�ĶA_�!��J�Z�LX�QU��ѻ�6jN)�@��`�����8�U�~�,��G�!hM����>¹�m���/�Mŗ�Hh����U�z7�Α�{gDZ��>q�&��h�b��5�5����L��'��W�OS�_����*�CAO��E�Y}�|��� 4�w�#W�;���WY*�b�9�)70K�sE�2�������	UKh��^�����e�DT��j�Q�g̟~!����΃��;3%�KQkh�p��(C�U�ЗO�j��5a�뜟�&����Q?5U�Q^a�<�o��E�E� �g�fR�$s�$�s��ïboT.[2�c�g���{��*�q>�a;��߀��v�M�z��ܸf�2���pml�Do�X���{�x/ 1�R�ˢ�=/u5���	&}���}��;�9=���[�NVE�J�2�(#�<��)�[S���`Q\Z
�|L�A��u���!�1d�X�7�~ͷ1��d��E�P���S Y<V�sS'�6������V�M4�5�j;A^����?Q�,��;n���0���	�s�񸁕���'���g�.|�7s�3����N�"3�8��
�8�g�^���O�u5?Nz4��G$7'p �ӀI���x ^4h��ÀY��yX'r�3�'u���su�]�����;�g]W:���Mع֧�?���!&}ý�<r�C �m�&��l�Sp�����Rf�}���q�l<�$�D��AN{k�Z�{d�h�,:|�nEā.�w�4�:����X��\@3�4۽�8�0�����+�	���+�0��v���<�1�Q�W����z��T5f����q�v��|��e���@9"<o��� <��*��:���!.x�Rh5�ܻMNt#�����N�~�l�r�vg{�/'���'��7��=c���^��q��>\���	���2G�����b���vkJ�O�	�����{Ԯ��F��|#���<�A��MK*�ܞ�;�ɿ�q��9pQ�X������4�_&�b%x_������yR��ѱ�����y.X��s�)=�$dw ,n[��ѰGw��y�H^z�g9�KJ�B(���.{O�D�p=�Bj� \�!],}	�E/�M�q��@�f��Cl6��˨�p�� 4�q�_AAM�	��Eʑ0\����k�/��7��)���M��XWS�ɭ��M���A3 ���&Q&(��H/��	����[d���;��ٴ�&l�%�`�ӑ����SU��aЫ�.� ܻ��S&�7�{Ĵ�K�'�}
^�H)W�S:�K���e��%�6+�y>e@�Hи�#H{t1���FD��X��&�3����
���Z`�h+��Ǚ|[6'�ڡ���_H`����8� ��x)��Y��o�D�����E[n�nv�x���V�BI�����_?�>�U�V�F�č1bk�����{(����8��e	�}�g�*�_��ip��'��\,�L���E ��i�@
2J4]!��hS��� \��KC���S�`���Q�m?�܌�6J���%��g�~��6��\<b����K��[����G%��2B~e/@d�QBO�/i��05d��X4�G��~^�v���t4��;[p��G���0g��@x��V�
Xп�!�eN���А��z���U'�����g�������\ �*U�h6��g���.P�U�x
fD��x<?�������%H�w�&�J},q�5f���V�B���O�ֳAHP/�/���ZFy�Gv�������,�?Q+$���re c {O�@D�R����/�$�������C����<��^i�+��k��lm�[�oͦ��E��'q�5��>�nI �lכ
q�M�fhGx57q�����q�\�$�ͮ�\ ��|Dg��h���t�3g��I^�'I2�6�����6���
{�~����*���Z�	����0y�6+�c�Ȃ~O�tM��GAaSO*�D��m��s�D�����jY��zmy4׋Z�fA�`�z7�� ��ތm�l����6"�ɷ�0q}XZ���?�	���uy-%�3��F�����O٭�5�8�+BŬ�X8�'�sX�9ئ���E�+i5�������M���������__�g�S�g�l��;7b����h��T��i�Jz�W���=����/���X؎o
���_�7���>!~�7b�^j/�k�z�` �\<���5�KFw��)�BW�>�}�0p
�H	��=� �џ~ٚ�{~�5$���T#C$��G*�ݙ��k�J�q��WP��5����6�b�P����=�~�9�I�;3�����+��$t^�[^ը`Nh�>����^��rs4a��W7CkQ����q��OW*����.�F�x�N�p�_^�g?&��窴iт	h�N�|$8|����AT���6��W�^��&q�5�pK^Mn3��o?s� ~$?����5Ν�Ƶ_Ĩ��;�k���4��7��1OY9ނ�+�rܜ�+Z�Ȣ�CٵS�D[$sш0��<I�J�m�^I���b
��a�/�y Oe��uk��ƣq�"X,����\ �.$���Y��3f�Yv���W��� G6D�a%R���Nw����Gg�!���'�9�U���#�����G�$Ɣ��P�UFH
--��e�1��ߥ�m}%��!8��-����P�eC�_2%���c������ʝ�:<�nӜ�;�"*�#:xr9���6W�
b����а�̛�� a��P���NJ�s�]�?��p#} �F��1_ԇ���:k�����%X�S�o����߾!=�y�r,��~W!�vz\�.� ���� ���@6<8����TIw��Q<�Fp�n_��`�V�%�{U�䬪��˴�9���6��������t��9x��](� ��R�n�,���|⊦�/2FGT�L#���u�X`<Q_-�;ͭX�"^=�fq��Q�Xg��L'��O-e4�χ���h1l��X]�E�nP@I\�R�1)�b�EYW�*��n Dȸ1)��D� "(A���*����"��O��#_*��+�ߍ�'�`ي�����AK�V��7!��C������Ae��|�5�W������ A �K6Ե�ѹ�[��)�&[�@�;�$���4�������h�o6�0�ç=ڦ�/#�h3�R[Q;}	�>�f����p�޽ ��E���=�o|���;(M��O��vġ{�so?*3R�J��-b�T���#
��hĳx�M�s��e����i�6#�T��^f}*�=蹒�}�B-�
��]��l��֎�c��ʮ���?����F�j����Dp"�r [�B�w�Z�׬��D!="�&���r��	OWĉ�Q�m�FP\�ɀ��_��A_�|O���8l�"���%=2�S0V쭓�2%=0'h2�y3�8���f���3��|�7�D?S�P�B	�~�	�X���{�ws[�p�n��gYD�6>��.�WG�I=�X��t�4ݟD��/���_ �d����3p5j�B�=[0]�L���; m37�b��������|h02	]��JT�t��`sps���,�=����vO�v�i0EB#rg	5漒h�w'�_:��+\9�'L!�L{�>ɓE��䈈���O2c�O'E��u�rF�[���(Cwh�Ŭ~͒��BJyGqz�����3��̀���T�{8�Q����hQJG,�?P0����u��J�����1��l�J���"�)%�Zc�������e�"!�"�
*�w�(r�ʺ��V�2��My� �w�BqQEˊPl����]�eF�C?7���{��>8�gs˭+�h���<{�k��&|�&bП-�>"�~<���l��`�P���&R��dԇ�r� d��9.o2����AB��McF�>�rC)����^���>�&��ZR@	��b|�o��N�?�nV�n!�T�/�v&�7�X�Hu��C"l�:+}�&�'��xD\MM��x�`>��<NT�!\�.6%��#�����cy������0-~�>���W�@�r,�cf�\Ї<�YI5��/�ڇ���+K&����k�\ؙ�$�-pFRi˔>˄>l�^�`�Q�3���A�+��t��H7a��!s��Q��c��u6����%n��i=�PΞ�֍��_X��Ώw�FHԤ������m�'3�(
�B�&S�7�ޢ���^{� 괭��%y�2���[78��Y��ާV�q'v�mQ�x�Z��	�<�nG�`ؒx7�� ��#��(?�E�vj#�嶺j2�\�8=9��ϗ��bV�Kp��2��k̏�J�	"O�P m�G�-� ͫ�+AqL}�^Ƿl(������<h���=���6�TN��`W�N j��b^~�tB���I|:��j���BH6(��	�1&u�m7�������LJ��t��
�q�M�&�#����G)�Ќ�%�*y{t,zD�f�Z �����ͫ�F�`�a�A&���������׹:�Z�ly8�0,�b�h�SV9]"��{&�h�q3�����I���Zw�ҝ�F��`>���X����P?�E )X@�
�B���D�/j�=k�Q���Aw�I�AF�q�I�FI�	/����)�o��Ĳ�/T��%)��4���đ�����u��π�'�.�*�[cUO��u�A�t,�O���6�ȰH���w='��L�'��L���N��瓟�3l��׌�����`>��g�ZĈZxZ �%<w�54�e �pYp2X�|�%�(vT���KU��M��R��#��WgN�����f��U��z H
��ղ�j���7p�ȯPoAշ^�1B�9��� ���ό
�N�E'�;X��������FG���&	N�]�C�M��\��˼�Mu�v�4�7��c|l���c�^��i.о��@z��#��+_(�|�9�m�#R����~b�_����b
7��~;츍2j�P�����X�1��>�	�)]��+��(�f.z8�_}�l	I��iyO��ƝQy&t;l�	օ�n_������-~�@+�*���c:����H�;׺.X1�~��t/p�&m;�>���෷����)P�z�"�B����hbh�/>�y��B1q/�}/U~#iM���I�cD3��`��	L����z��5�ed
��7����Psڐ�:WE����4��O����c���4���ʂ��N�c����:��8�Az���F�e�M[x06:[L���gk/�s���s����Xv�HMN����f�.s���9�k� ��.7�&$]�MK�#�]�}�׃��Μk2&2�뷎7j:5�>ܦÖ�����9������	7Ec�F��#��{��5{�,��q�:c�B�w����A��OnQ����Eua��W�z���YT�vL�E����\e�=�i�0.�i��Yg��ڤ��f��o,@q��%���}^���Q�v����| �%�b7f׽�<.�2�uUp<�4%g;��~]�u;��(�s��cz[�#��NoΖ�q�e3�����E|�JX?]��lG�K�fX}[���Ȭ
�l�P�%�J��ߔZ�S];�b��Y�'���&� ?���KhV=tl�-m��[�e�Аӣ��7
���4ԟ4����K*έ�ڝ�%�ez᝜�P�*A�\X���o���E_}��f���ギ�U�2>���QLW�oguc�fU�i�;�G
�#�kLvN�Zt9���!��7U���>����(
W!&U.f K�j�܁M�?]_WS��UםlG�#s+�_�|��hX�y�hj���%����&L��%�ݘ�	�|��N��"	觷����yot��1�dtV'�ƫr��{��-���,	}�x�K�w�b�Ai�sqU�o�>�閙#�5?�9S�oPC�1��xS�z�������k����2Gf�!��b� �Ў���)��B�zfg��i�ˏ��&`�:9i�k�Dtgo�]ܢ7%]��A��vH����h�����mprb�/��(M��@b��ğ�����+�!=Ͼۂ"���lf��\��3�@|W'�,%��Ww�����'3f��;D��{1���:��/��H1c3�,����_�C`���dr�Ҁ����f|mc����H\S33Qq������+PKpp&牨ĮD��j�.B~�R����%`�-")�����6�`$�<����F���k
�j�rGAy9��&xGzͧ��9P'&���ӻ�k�g g�A�����u�zI��t�!,s�_[Zմy�mڣ)Λ�8Js�������0��@�O,��F}<X"m��؝��0�/�'��Ԁ��OC?>E�
�΋�>��!6#�Jf@�qй�!��Q��ћ.�#��O�����i�k�e�?�-�v������c����o��{9�����{@���AH����� ��#����Y�g6���ſ>�V����6 5-��X�*j|��9?�6[��wco���&�e�-�q����ݚ��L�����$ �߮�%��ױ2c1���"�W8���-��40�5�#IwxاI���쁮�0<� =(6Y��ٯ0�9nD���!k��^��E9a;	JbJ���p��P=��|�Q�b�B1�N��W�%Mw@�?��G�O�O�W��n]�H6��1�s�w=�4
�;b�[���7�"���Τ�D?V��sjW��'��b�QY��ω��]*j��$rI�� 	�����I�)v}��x�����H`ܺ�[�������F�����xN�-��=�sJB�����$�>��ON�!����u���x����[���y]��hF�%�,QŎ�v�vʳ?L��f=RfD;W�Ypz d��Z9��������T��;;������9
Pغs��d�~V����ZJ%�\��؁��R���*��{�(�9L�`�qu�1:&�1/��pI�S��2'��:C��W/\{�e�p�fE�Q�$�,yP�O�|�1W
���$k�_ѫ�F_}p�Y���)7�W�O��c��Q}�����q.m��֪��@�FH���"5s��+�>�Xi9]5x��朞���`A:�k�k��}4ip�����������[u���f��`���g�eFK��|�*8�x�*w�+ fc����;��)�z���0�!�RU�\>p�������{/Z��o+4�>>�sغk���j�U_�<s���j��IZ���M���!5F�U�S�O�3^�I�h������V�ד�Pc7���I��wbuu�x�0G��j�m���-$:޲м������~l5p�u�_��	���aؽH�*u ����+�d�c�?"��t���	�A�/pn����.�bU�ԫ.�T��t��P���hR��VZ�%�M��%�����m�!��sq~KtV�w;-��[�A-ǹ�|؋���O��T�	��ܞW/���B��[e7���[��:|�릶h"/�H�Aw=�R�\&h��7�H#���@����ܖC&����<�rh+�_Q�KT�Ql�K���,�הC�{�d2��,l ����>�쵺RP�+! ��U'~q?�����[8k(�p4�5�.�D��'��-�D9�~�����ԭ��sя	UC���%/0��B�,��&��c[�c&N�t�Y�)9���b*���ӥ�����2��i��q��%���
��a|��Si�y̋������6�Y�_pӦ�¤��x0m*�,Drѣ�\)'e8�P8k�����(�k&��F�u�ώA+��orm�s�s=�9����MD&G�*�P8kxnm��ɋ�e����^�m���l���9�69N�0�s-ydN��àqOZ�I�&U" �c����]�����iL��$@�]k�+>����@%K�n�uE���:a���kT���7�.���*;_�\���I��_�MW���@č��eOB�_���F"�W��kB��z�.~�t���Ƙ���˾�����ᣀ���Wk�D�{}g4|\��Ӭoq�-������8��e��I��_K,���텧N�܈I�L�.����<#�ɮ�/�8��(`S��H��괶 �_��%0��;��1��b�ߝ6����qkZЛ�Ѣ���6�=�0T��qF'!2��G��ynƸDcs|ګ��B�V��]�2��v׶ ��{�%/m�$%c�mu�^��X:�_���h����cc4K�J�2KZ��D0I��,�ݛ62'c�Rasq1B�=S�9��$��V�j��J[��5��]$F�C
��O�dу�k7��{ߘ����4՛9<�^�����+c�GO�l{�ql�F�������,}�cha���9��7�޳n�0E�&�UKE�"��Ε�R���������nh?xv>�=�	�����.-`��:@{s��eV��3����n��<�¡D�����-�I�ZHm\][�6�q4�$������6��Xط4g�z?��=��u�^ȃm���X�t*(M���&L[�f
�ݥʘA�V������441 ��H��� Ǘ���jsV�C��;b�I�ߔ�k�-��@��a
~��f��M})iw��T4�b��b�_P�f��&����\P�����`���/���k����WGCA �c����?^~(K"�͕�1�w���M�=��S�i��}]6N�?��hS��؟y���U�;����֜g�t�:�IQ�|-6ݙըY>���t9 �b@V�87W���Z�f�f�`�\Nĝ'%�X��f�b5�M޲䦟�>q�A�9��g=p�*�����&���;��+���}�AC�������.�y>]bE�8;gf��u�^&._:+�>��Q�0��:��}�o#/٦y�����Y�V�1��%$������Z��j\�XgS�r�+��X+P��/������j�:t�� �: bxB�'
�cՖXP�Qkh�~6����%2�1��4��ж�Ò!;@�f|T� �����F��͑6+Y荳^��8�X�����p-�5�Υ6=�l�M<��q����\���6
с����	|%?��N�tlUuZ�/�n�j�W���Y[��4��
�'|W��Z�����L��g�8aX�1�E�	^�b�:}�^���Q��om}�m���-�������_�(�v�(�U�
�Fͳ�5�C�d|H��g}9q�0%Y�������a�R�K
��C�Zu�(��nAnD/����r���T��iT����k�wpղ�+�Q��1YU%�o��m�����y�oPߒ�Z^�d����%{���0�]���u
-s���I�����=���`���ye�Լ�77+�k��뿘'~��ښ�vTr�'���K�O5��d�(��id*.d���6�-(���~����}�RgR��f͇�W��[ ~��O���2}���J�`����ʭ�j�*C!_?��kK����YV�
�eR�����z����7@�L����h���G+�R��	�2\
A4QϚ��۫�7Z��R���Uр4���5WV�;��2?\@kY	����~LW>f-I��lF2d����1�A	���M;P萮�C2�M��������1�6�ޛ4,O��{��♁�B�S�X:;���)ڒ�JF�{ߋ��������~��o?��L���%�������}>���cE��S��{��A �Me"k���]3��F窱�����ԡ{fQi���me�K,Lr��3���A�nEg-����]ςǈ^�������F���k1���kT��x�I����2}������H�d"�Ҍ����)?S��r�м{\�3L�uH���;F�\�;(�F%����JY�_-�J; ������(��J�O�;�V��+2���lL	n�~�A�.z����)��n��~�=�>W(!4���4.8�7�������=E�/��i�u���{Ӡ�TY���
�<�$�B*��|�@p��y�Vnb���}G��;�>�An [O�^�� ��X���]�m��܎�N�#y_������V#G�3�o&�՗��~���-)GH}�����9$裚 �r��@�ť�w���2�F^�]6d����ԩh������~8��x,6�Qy �V* �,8�
8�e��G�zӲ��N�����l���g�����[@B��u66��N2Ϛ����YRh�n�ޜ��#gyƚ�7�2�	�d^�y�z�	��.rhᏄY�/�Q˲y��D*oC�|$k�y%���������l��䲭�`���k۹͚�1��_&Pc~��m�<D��pʮ��x�a����X�$�(Qձ^���ju��Z��ғ�[��0�����B��}��z�&��`��'��6Iա��\�?���ާ`R��pr�(U�myz��ױ�ǿ�5��Gk��1����Y�u/?��R�A{`q����c�/[�y2� �K�`u����69����u٠���Q��Hw�6���A��)�ˋƻ��u��/
6ǁIwgb�sH���/hS��бHF�哼l���H �)��I����/>�	X+L�m�d��<G�"i��DPǪ9�CK�uy�vJ,���Q�!�gܿ�H�sG.���R:ܼ��r:a�䈨�!C/�l耱�潎�^�=�<n��l���
���kȱ�妦6��^��#V�V��}�J��zP�+�t��P�N�9S��k>������f����6�����<�t�q�����q��r2J|��"*���s�@�?���|og�����5�.�N-zi3H�lnH����N�	P�oa@#fV򧶩>b7Nܐ�c~'U>�^m��\�WM�I��e�а6?^���܃`�bL(�
��D�±�����h��;�Ǯ��W"d{�pZv�[�e,}��x�._�]�v4���h�,a��ᆚ��.�*��޼8��{���k�7[H�~j� u�ן�b��D!�9l#��G)\&��Ld�`��$5,�s�6���$�w!�!�^@L��܏AE�iƄ9iІ��W�2.nA�j@�Gְ&�l�}[yw-�d,`���y	6!n��Y\(f������-����K;�|��~�HM����S߷��ݣ�a�~���$+�a|}p��������һV��T��NH`_��%)T]����Zq�D��E��O�_$q��2���a�e��"��:m)l&v\,X�����g���8GU�Ua8?��1�YQ�
���yf"O����p��?�sl`~Y��y E�gȼ3(�]�q(t<�r�+-iW���Lg�@	`u�{�0��*K6@T���=��0 �x�[rǄMD���Y�H��������(��ؕR�q"��Q:T�̷v���ڷ�Z����o{�g4Mv_�@M����0d�k�d`���{I�5&�Gk�)������X9aA3�deɚ������ G�uA��b�ުY]�'�$�xǸ	R�.0B�9��9�S���XOt�Y=�$���V;C7}S~{-k���}�'�InN� ��y�i[i *F�En��)��c݋��+?W���Y� ����Ǖy���mE��U�ɰ� �����C �G:�bB!�q?S���D��� le
A:��}��G��[B!�*�n���D��b�D��d��q�1lңk��2�W>��(�A�"6׍�l�G��LnW�p��.�-���������ډ	�s�� �#dZ�x�|�μwm�+��E2��]@����]��_��7�v��c@u���xBrW5�������RㄘF����GYb�RЦ3�gk�M��)�?�W�YG�qd2�b�/�s��۶_�9���&��/�����'3�K aă�M�i`���cL���c��o�:S t�	�@��Ҟ��r�!@*NC����/cX��N�֧�Y �iM�� (:ӕ��n�4a�>��<~�^�W]�T��	��7&O���	Ȟ��
.��KdꌲTNz��¢D�ܝ��.����"h1�F�6�4r�ў�X{#�;��z��S�SM���5�`�_�2k���TZ���o.���=�~:n�����}mS�Qʹg���9@�~�a��X�T�:K���g�+��O-eT��L��yE=�\�����8�>9�fju�U��|���,<������]�����E:H#5-�_���3��<2R�x�����$&��1��}�k�K!�S��nr��A�]�:�l���f�Z�)X�N�#�+w����tVQށ�J�6�/��OK�xP&M���a^3��.�~;/�����ly�:�q�Y%i���vI�}tW��{b��%�m�`|�3`���	�ίo]�����]Σ{eT=3T�����pH�����ߤjCͨդ�E[� U�4b���1~[�=�L�jWߔNt�+إ��}�>9���Wh�MKr�
�d�@�R��&��3���>����yn�C�����J��Eˆ*�� A�����"������m`��o��-%�n�Jy��flW��y�vUYXs�U;���v�6ج×������u;��d�B9�y{rK�}��ov
Mz�����5�9��5@���8�$����{Z�c�;��xV�{?b��NcsL{�-~���3�y�{�����лG��F��70mb�ѐ�.aCr�4��+5�p_��ó�5�9�cbm=-d?��zz����J��0�"�'�t=�����M8�C�U��0� �Ο��,�AJ���t����3E�����]�;��k_�q�Ľ�����!�?i�����:�]C�^M��AN����瀞�R�� ۖ���Ui�{#�k���b]��ɮ8_9�>Qo@���+d��`��<q�؏;�&�ۯIQ��tW�^�/6[Ӿ� �����щ�V���^����o�ku��}N�6��q��i�5��},0�?Pݞ��p��Va��3���Ѩ虄��_��͐�6�����p̸���$r��L����TԘ]/>�+QL������
�x,c)p���C�WBg���1����%�}G�~�CK����2���Tz��m���������!�q���o�UP�yj���נP� x��!k�9:��v0=խ&e�Z�3zy��B3fi��̿���>mrl�F��S@��SL�nI�]�s�ꄬ+SB��fL� �wT�:�6|��/�P~�mWuʛ�k�Pˢ�J�x�K�����v�s���?6��#��iF���E�c��"��ZRhNDү˅φ	�y!ː��GE��ղDe�?[��	�����t�nHn#���`'<xxq@�9	�e`r�y�P%�?B3��ѻ���t��S}�/~b��#:���I��WXV��!�݋cˍ�����|��y�}�D��`R�+Y�3����4�������ȅ��	�����n�^��eD��<�2
�ۗgt�L�BP@�|�dRb]�F�C-$���p�DH��,WŭaR[��RI�:��Xr1�eоi虚�%˺r�D�n�?���픆���!��:�~�Eyk�cHuom�J��W4r��E�s�L����)Χ^�$�Z��\���c.tSe�횴ll�;-~u�\��>��>3%x�����O�I=s�c�R�����R�b:����S��gC�D�c�irS6ekF�)"A�1�̍,J��Q�޽g�"��]�pip^��R߹��v����p����K7*~XB��.r�_k�A�&��i�Ӵ�Mo�s��(
g�oǄDSH��œw�!�X����t��H�iL~ Á����K��E���ET4O1I�S��9E6�^iU��m�@�3�GJ���,�MU09�tp�ݯ9��;�.�U�z6Vt�;���5���	����!w'�?hƲ��1|�0b5�c�[�,��ba�w:�4��uc۴D�3S���jQ^��;��A�u��^�y8{�{�"	������Hn�]Sl�'}�/ߘ>���A�?��>X�>؃b�FWFL^�@z�/��X���*��r^_�{�����$���.��i�0!�#�
�o�Ԝ��Bj0nl�H�*�:�n���)mK�4�B�X�|�Na!��h�ʾ\�\��g��jJ!��M�0c�ҕ��m���G�i[5��ȳ����/<��H����^L^�hH,B[f덣 �2�͔�m<���cT��P�?`ٿuiGH�y.JQ_dJ��7F��
w��90'�&L�C7�˞|��0t��S���?�jL����ŕ7�ԗ���F�/ɦ'�7K�{��s�͔�UNHI{j��Q1{���ۨ��t�Vg����V�@���W�^��:(	m���5��#��1A��Of�BX֩�;��}8�[R�wo2�#��0�m���Q�vl�v���3�S�w��?q"�Y:�N�tN%{m<ߣl۠H��Р��P|U	f�HҸJWr�'LŸډxVS� �[+���ﴏ|�I�[��5w9j��y×��
	�9,4ڸU����0�/�#&|�P��jEmN��=J�����RbuΟ��w��B�8���x�0�rl���e	 �����$ �������R�����Ӟ�T�q��w��8��y��y���+�N?ڐd�8�k��A5�]p�bSO�!�7�x�d��J��	<��4']0��HiC�!U�K�:Rۀ���^v`�bo �
(���?�F� 5Z�aK�go��P����Cj��j�x?�iH {�� AvAՕ砃�F<v%3b�@�����Š�'��1��!�Ǖ6�E~m.������°�'�F��~�է��6\�X�"�*�Y(��lL|���/N����`��@�V���K��Ӗ�P��ZbU�T�,��%��b`@�?.�Ѕ��� �>����$2���d�%8J��A��;��gZ����/�:!`�.r�˄��
X��A� ѯ�ꅮ�WJb���?�bo�F�O�=�f��w	� �n��h�t�I���`�M��j�Vݦ�����^�������j�&��נ({�5�٢J�Jn1JZ��q�r�,�ZNPhv�_��b�T���s"<a��Y�7�C�~4���?��Y��4QP������n�E����s�J�����9�C��D50�scH6O.��n<_�/����T�Cz�����q|I��Z��"O=�! mcy"6��,�A�4�#���lˡ֠&�ra��W_���Mh�}�^xS}3<I,�C�@�"m�@ŷ�F0	�B�\1��O�J���54d;2I��Ỏ�*Y�?��|s��'�+�	�5����@X��+.`j�@.*� �EcAQ2�]g��m�����UAB�y�?�;���d�����H� _e'�SPeH�5n��b��%�̓?M��4�����6[~f_m	j�W3��<�*:Ȼ#�;[3e<Y��бO���������r �Yl4�i����ݡ�2�$�"cI���ݣ�������y&��/��Zn�dF������Ͳ=3��keB�pz8ݰ���kZ5���*FIvP�������?�����Vo����Y�\9��l$`��ub�<�+�������k�Q�6:���E�y�O"3��N���Y�3WD�`w�u�����A�ڵËm�'\��*�<�T���|�l7$>}N�b���=���[<����ݎ�u��b~���qV � ��	V�]B��Ċ���ҏ'W��I���"�+ג�QP�Dl��1������M���Y!T�K'�DG5W��8�CZ�\0�w��ՃVc���:kzH1�{��ᾁ~�4���.lt õC�M-���9�(a�dȤF�bkKc�%�c����D��j(��	�r�d�O��rl1�e�t���A�WsV)8�RM������8�r`hc���$���z��^�ǳ�@D����!��BP�F���Am,WAs	���X����%��mdQȹW'��-a#���M���OD(Xx�\����8��!�ڌ�昜��U�v�/i��CS������rۅ���`�~���I?ս�u�)����d�@�͋`B.��͐�[�e�pp@݌&>Ȝ���v��'�����r��Q��'�#Z|�}���%)ݍ���ˤ	�'�6���R�}.�ʣn����~1 �6'ivӍMnKEO�2r�`��mF>T�4w{�{l5���h5y���j����4컩�|<������k���tܯ�B�y�Ɵ}J��$j��l?uy�͙e.��s�a����$�$Z���,O�g��n:�x��\�`�ަ4��z�=�e���Aڒ���ޠ��y�~q�!������	q?�8��<Ȍ�/�t1Ըiç,!��l���'��q�����^7純����������,)Næ��������i���Kz1�� �:ծn�('Ș��E���-����n�׋/�Ygn�ǩP'/p��*5��lN\�_�X�6�ç��%���>��o��x4�;��Z:�:@���y�[�T4���� �d������1�5��5&�7����
���ӥ�[�3�p�^������b�y2�xo�k�,-x�W������;<IN���9�ꀦ�w�Lw�&d��;h�<�~��.=����-O�*K+�~͆˃@E]ƴ�'A��~�^<?m<���/�[Q�?��_�u�#X���0R�ڝ|~����8���o�����	5�)��xE�����1WO���jb����_�Y@2���F�����M�p��_��ثITZyVC�C](S���t(�+:L�
���Mh�z�!^�)e�C4����X���|�.�Ig�4�Hi�";PΣ+ v��pف�-�եYPᄲU4��Nr�8Pb+_�7��cL�X�	[Mę��t*���DL3�}�hxg�z�U.�3d�8V���;��tC�sC��>�E��A�mײ���G�ߞ�� W+ě:�K4<���f�7�J;�H�������-�'��p�I�j�n_�K�m�!����~`"b��	�<:���l�-��5�Gr����P�L6�@����е�1*��t��_9|#�����{4��(�޶�|.����e=1>E��oK���=�҆�YZ{��X��-�!�(�,ƣ�?3H})^U6���5����st1)L�1{��Z�/��ᢿ����<wKa�����VΌX������h���F(������<�K�gm�V��w��"n	
z��mW퍂���ƺ�$���M3��[�B|��<�=`O�G^<��ZI�66 L���q��bSZ^�F�*{رA�Ç���.�ď��G�z׏�|�+�ۗ���#c��-��cE��n��'7�1�31�JUZ]��N��}��\���ƃ����V�Պa��]�H�Ŗ��\���h�H�����©6i4���48=H�ӺY��L>��t�0�5�X�p �K·��/ԫ^�c|M��gѠ�g��*+��ON�ru�d�/D!�G�����o�cA �i"���\�m�N0o)X���7�罭M���NSp,�����+7��D�E�ګ������SM�҈�rN	SgcU_ݍ#$8Vho��,�I��f�>���P���ʗ��x� �z��F:!�[]�t�G=^�K��pLo�U������n��"`��OF�/�/��X��Յ&�]\��q���!���̓vO	d"�z�|��D��Udt���T'l>7.��Ϝ� 0%��<���^�~���G��<�����~�H"0I�Y�����C���wrEB,�y���ι�A9Tv�l��cm���d�¸��7�)҂�ctZ}?2Sh�����>�7)X�b�*��q��vA2(@ӞdK;�ˬQn� �0cA�	���-�6T�g�F�.�1���������xr�ͻ|y2��p_�O'8�����6@V����G. ����������=���VX��DqP>��S�ލ��T��mr،]e��ԏy�ۇ�u����5^��� ���؉�7��bf����u�*j�W�g�������5FFy@�$ S��0��,¹�����	g8�V��i /�ׇ	�=�(#�ՠ�}i����a�6'tA���̩�I���j��"��� �̅�ѧNF�sl>�n����'e�H�ڷ�1˝{;��5B�N�|���}��b|pns����w� �i�����hk��vrn����Z��V�3i���N�M�;Dq�h4�^����mOaTz7�3�$�܁*=����#�p*��'��s̉ޖ
��j�IEў��PN>y}p��`D��.N�)J���-�����nRU|/��ۑ#�#.4^+�(p��y!����������|��x!�2�t΢�V�>N���^3��[�n�ay��ݫά�p�VĚ�w����!���yd�
i�!R�,��1 �'���v�X�!�)`��e�j��F)���e�����J�v�������Z����N[�����)�T~�e/�@ʾ�nb�����D�P�؉0X���scZ���R3��9u ;�RN�d�'ٖ�E���1qs>L��IĆ����%�����j�M)���"� ��	�8vh�.z��ǀh��l�yg�q˭�.	�us�uR���V�JxD�����.�ݰG;��Jz�X�/�
hm�����(�S�0�8B0+��i�VsSJ��` �S�lBD�fБ�P4��V0|C���B)�n �I!�x�IUN��S�/�%�9\{��z�W�Y�uz���D��~ҹ_R�B�lÁ���������+�3p�|��F�[hb����*N E��uC��ŜB��	r
�!�1% �j7�a��N��w}u��81�gO&�\1VJV�`��*�_!tqQ��{�������D�/�{C�������4	6�iG �=�����VQﬅ���=(ji%<���6�+�ߎ}�o*G���G�8N��3Nz�n^J�M���O%$A��d3e�9�f�ђ�*�nA;L��<��?�7���x���ܙTĈ۳ÿ����`�BȔ��G�y�ߍ�YЋ!����Dk��Q�j*�)~�9�xJ�M�����M�!�q�I��	;�!\\�@��v�O��m\0!c!B�f�e
�+����iA�(̻e�s9Λ�}%�k8O����/P�Q;������"\�4�I�>v�`p@�p�d�����IP;�FR�ICJ������2��Zk���R�>k?*noQ�>��UϾMZ��%Boe�Q�k���V��p/:0�m4똽C���~�`_j䬟G�L� �՟)	���i���y����T�H��<�Qe-ct�� �o5�2dx@>(i�< q�"
�ژ��Yl��X����ռ]�ٺ��{�7�6�X��[Eb��5����{����l���R�TV�ô@o����í9�_΢bBw��~t�;�@���%�5Y���@)Z� ��V#(2�K�kԻa����R��|���&&�9XJR�ss���v�Ev�LT��(y�L��|�Pl6{�G�>-��B���L%�����?�dӆP���BR�'H>�K@�\���x��@���ǟj���O���^T�����d�L�\�'2� 3p��mvs�;�^��#'��Q��^D �
��>�������*���9q�`����E�+��� ���s;�9���Gv�Շ����j4���e7�����& Ȣ��n�Y9-�zJ�p�%��(č  ��tyF�\��d��3�%u�̨������u�/B�PH���{�sH6?��{FZ�UL�;d��Uu|�!��}�n�1�L��<�'��9��H#�9� �y�2�Q��6�^���Uz�6�xV��N�~Lt_^�5�nL����zYB72�7w�T��&x��1���"ґ-@͡��_���{������aT^i+�~�dԣ��*�6Vn�����-㵏����?ߤ*s���K��L-ú�޵�(-�����b9��~2�^�f,���}7M���
S��$�KXCxaO�2�����z|\`��P�!����
<�wutؾ���������?f(r�\�ߠ�Tu��Cl��9���F�i�@\i#� �U&y��Os���j�\$��o0�6�;t-|i�D�@Rm�zݣ,a(6%�op��C�\~���#��������: ���G#��x���T\_��&0�f2���c���SЅ��[��>�Ł(�4r�IB�N �������RF�y9m��q~�S��E�~�i-����B�~=X/��z�m��GW�6���Ӌ�zIimr8�nܧ輳N~h�����L����P/��;�L�9�>sc%���	Ȟ�T5WE�Twj�,�t�	Q���C\~\�����X�s��z�l����D�?|�֨�Uy ^}6j��mxg�;��J�U���xr���6�����l���jhN�"�>��C�fǿ������-r��N��4#Z�R���c�Q�MWN6e_j���x�!�����M��gy��77������0N��^C��>�Ȝ��a�_-0�'�Dh�j{�}����e��Y\}a���Y��x��ov���x�tx�䱻��^��P�uC@���B3��� ����R�B�dg����E�a��D�}�Ǎ����n��Gی͢�m��J�������ubq��ٚ%^j���q����e���;�=�'�R�of��2[e�9��k8�X�Ymv	��o�}gn��$��Yzȍ~�A��A2X��=�'���k��p����!d�U��el<y��Ҥ-���}�k�:���QE�^�i�Cwa�=��3��e+U�I"�]d��?~V�9�<�[��`�?e����j�})�/���Ͽ�n��<��Eϵ�'�2��"���ۭ�렿����������?g��S�2V�E>��B�{ԩAA0��3��!��wx��8�)�l����-~��o��=O��|pE<Sti�B(\J�nc�uD~ ����<�x��ӵM|/�����ON`��l�xː���6���"�i�l-
|��A.�� �������1c
j ����%k�Y�N�U[�a�-Lr��c�p)�P�h����8�nV�x�n�@��=�9��ܤũ���z��Yn��c���<�)�Bi���r��)�F���^'� �R�v�h���&=
�sV��?{ =��?��d	Яj[Wi��
T�o�%��@0��Ξ�_���Ե�~�D�JD����o �P�2q-��/7`�;�\W�y���?I2��6���Ub'���`�u ���0M�)<�M��U�;9��
#�WZ��>����U��i��9b?����H$"~{V�y���$^<QB<|�߃�<�V���Ø�����T7u3�SSz�s�W�9�Kd�86S���]���e�{يn	�XO1����}��'2j�2�܁�7������k���  �r�Ϲ�I�BK߃*�L��4a� .0,ZÍ���s,`�ڷ�s!��`�a����v�m���׬���ҍvz*,���{���5�6��a�{o޴���|�g��c+�c۰g�IH��c1�暈O�F�����x֧�3�b�6���B�p6���Չe{����)�Bُ2} )�LDh�]��f�s�`���T�j>7��e�S	kh#�#@�l�1�	��X�Ԏ2�"��p��z����$�"q�����7i#��"������Թ'hD�#}��փ�*��9���ߨ��x�Ѻ�O��w�~�X��\��I"��{�d#w������Dy?�ދ�e��T U@.m�bٳ��q�ly�����R3�`�ʫO �΢Q��v�-���n �i�3�UU��~�j��Q�hb ���[w��1^�&��k�r�x��]��D�T�jtoИ�,\(@
����������G�F�}b=�!=�9�2���js�%��;1\��|aaf�K裿M�S���ؗ�RfJ�سϚ�!a�j)��ҥisҔ9?��4Z�{	�ɿ}����nhM��)������j�n�U%���U�.�vlӦ_APu�{ie�$(�;m��+(1ɢ"����|a���l����ĸ�*�u��*�0�׽){.(P=�
���o�L��i�.qT�b� m�!n�?qvuw���!|�	`��kj�H8Z����]ێ��gk��h0�-���a렭�UH�;��9�<����/!��'��9z��t0Wl����}���U_�ϯ���Kr��$�ަ(�5U�A*�>�`~f��`��DLh�K�n7f,��XnV�W���@�Y�c"�}>dC���iO+Uō��*���%��e]���}<��<�!�"OGYD��V�.���[�$���9��}�%'�T��{�T�S��}�R)��l�R��<��
#k	@����I���`*��]y������Ӕ��^c���b���u~��u���-,Ef�ͪ��rQ]D�P����؝��OH�F�������)���)zi�[��t e�s����?��$i�a�f��0p�$v̕H�a�y��c��/[A\%���zK�6�Kl�7���=V(�!RA9E���\#�Nʄ����>ȼ�rPKwWe���C�q��4��ͤ۵��<�qB��=����:�=�`�:2I��H��a�p��^�m� 53�+跷����}��j���������YW�.����V��v?�β�#�f�u��e�q<?��F�U$p���\y�6%�b�Vr@�d�p�m�N��f=Z>��ãK�ܐc�琤όd���	{�=��
�7l	�e$g7�#�"& �O����Z�fK|�D��(($_54�"��Z��*�6A�4���hZG��n�@�DLA��~�}��m�Ej�3�Y6\2��^�4ݟ�1>����(��o��i����1T�!���Æ�a-��(��&?2LLo������c����6���w���+�9�e<S!������[�@'��Rf���Ps�u.�����C��vЛ4��Į��d`��&��g:�=�pmm�+gf���$T�"�09s~V��{�!��G�[�;�;�5쇿E}z�~�֢�[���Y�?������2P ���L
Of�C���o �`��~\���OJ$
�7���Z�֘0�"��7�U�cA7������$�w��>��c:n�0"V�>݁��y��^m�q��E;mA����5�n�/O��vP���-��,.�l0%v��:�]��Σ�ù��?��i�5�Bs'K�M���#�-�z@,"�!Uf��G"]"¶�G�D���~L2٦	�g�T����q�kP���O�͔˽�G(S�hr+ʿP��L��'}��館��r`����]i����E����S�ɓ���I��5��y�ju퓖Ys�,j7�w+ߊj�/PVBձ���7�4��KY	[� F�g�Nt�E�Su��ʓ�~�"r__�,�.Jw�������+��o�����ʭT��EM�n��������[D����[���� ��IͻZ�2�r ��ѝ��|�J���O�7GڣW�pɢ)^uk�j������Z9�V���Q_0����\#����	���x��[l}ޙ̭��H:[W*0�&ya�7�����2F\q9r$<Z|'�D��d���s�L�@ͱ������3L�;'�	h��l��[�������i�����P\�d���Iΰ&{8'(T��GW5��w�_o&�T�����[����H�k��k�uؖ1��*�+8�����_�@&X��qP�cM�<h��
oCL��sJ���q.HX�8����Z5b�$Au�a+3�aY��wyr�"�c�ň�IF�T%���#�~�g�K3c�P}N�#E�(�l���&_o��v��=�A�*� ����ld[�����얜*��~�G��C�&q�ߎ�|��X��i`%n���-_Kt�&��9��\�{�u��١�z1Y�|�*�� ��׿4�U�sV)���a!��R�u�ý��GY�]Mk6E�����m���;�I�����R�4ߛ���G&�Z��9�p1
}�Ɲ��{�P����j����w�g3c����E�7a�&�`~�Ԋ��79�9���~��0�I�>�\)��0=H0:����k.���\�k�ʁ���u$I^��B
^o��,�~=`vO8�7�b�ː�x����lwV���5��:c�����P�;GOm�w5�z��R6��f@[��������X���޹��?���
�b����)���\���K�ve�$GZ纴�mu�a��3���j�{���F���HWW�WI �*@�ݙ{;HA
[�b�N�ӿǒT2������sC��]\u�$H�~�̃��n����ݿmu��=�K�?�|�����6_�qCXdK��gI�N�F]�mJp"�(���ܥ�& 
"�i<W��5+ܬ!
��t��kX���s��*џ�C{?D,��~'����B�W�$�4�j
h�w��Fq�t����n���ǕO�"��r�e���T��{N�|��g��8��<П�$��q�ւY����5��w���UK�f���bÁ����Z���7�偊���0|���Jn/��~�B��m ��!Z�7#.Tu�w��
�LE�0���%��e��� �@++��Db�5����@��V&Ni'w���[���]�B ����S��¨8؛�0@�GV|A��V��e�z8j��`D�~,w�>�_u��is,��?��exAo�e�w��i>���,-ͽ����)*���U�P��4F�0�>9k��A���	�	��c����u�aB��3Y�ݻ�	bx��#�j�(���RrbC�޷Ju�����ǨO�A#���K���2尃������j|�w�]�YUX	�Ε�1L�+Eڧ��䤯�?c�������lh���L�|��X��g�P�$�x�1�<��V�>�S���`O}��K�Z�Ů�p���UV5咭�7��F4xσ�E�q�f\��_dQk���Y����H��	Yݞ�F(��:�Z7;��i���i��"�E�y�`��w�j�����뫀C��:#$��`a_��p���w�>��=�'v�-LN��,\u��QY�I[1�kJ�a�g�-~`����1(Z�%N0��!E��l?i'm4����[`�Da���?#1Ee�>�LP�u��Y�PWU���)��Z�;"�3K�,@g���fz,l6�f�K�����A����A���e�H�����:#��P��r�v3W-^n�:�p�����0S���9tӌ�x5� ���/�?�� ��DI,E ��i���vni���	Nxr��)��4�`;k�.9?z�$F)�Ӂ�<�X�m��[7�T�c�/U�o!Z�ON%`K��}���@�K�T��O4��=�p��I����S���Yk�Cz��k{��u���gA|�!�B�	%p����z���8� &��c��u�a���(�偔��ģ�Y���Z�D#�|��Q��D���;�,�r�_P�bd\oͷ�e>L�bC�_����-��5c%#�]�J�FZ�P���#�8N	)|��=z��Y�.���g;����"6���!��3�
��&n�C	x��`} ��t������V��Ve�%Ѓ�A��t+�!B�f=yV�mg鐂�
~2�n8��{g�5�A ����X�m+�.*}�/�������6��vEّ��ް����ӫ.5yP�y�۵e�[��TՇ�Y9���^�/�8vG��i�`�'�'�(��\��l�R�+1��E�a7B6�2ѭ�*xJ9�T��SX%�
����yeC-p���#�si�ת&�ג�M�a��`F�IwFS�QɅJ��8e��Ͻ~܏��E�,�Mhq^��@�sߩ{z��.��ו�P�Tٗ�96G�m>P��u�U�a���'R��Ʈe�H4��5���@�G�G\K&RO���k�U�5'����}۸��lvr�m/Ր� �Խ�sz�s�N�j�yk--��I4@��q�M<�g{�A�d�[�����jҁ�eU&�M������3e~�rt甐��#Z���z�Je
����}��	��G'��h3�'���IQ��`���.^�(~�/����0{����
kf���p�gb�i�O�y���*�ľ�W�Æ��f$�g����Ub�x��=��M7)�|dU��_��M���{N�!G^�?ǵ��t�t2�]X��x�B����&ő6��/Tr򳎯���v�0~ݭǞ��y�^�B�	��6��ԥ�A��F��z�}r�=�-�����]���8#6�k6|$g�It6qyz�ڟ����3�2nkI��;1O#��+&b�6���/������)g����Q�*QC���9�Dgr7�`d%�i�g�+Ib��Zo��&W����<*�ew�`{�>����th���q���P�����e��� )4Ӟ�J������-V�Q�����	,��f���a����t�!9��#;�n���hf*��ˮ���t�A"ъ��$�5{=})�vO��:�A��S:DY�o��K*X���ijEp6����M�e8����a���?�+8Cv�Q��1"���U���5�}�x]��T �On���6�$���-��uMe�5�_f��W��봡4^�9_B�"9\_a�S�%A%�
�q5]���f�Bsߩa��F�� �����jc����\�2�c/6*��c��S!������,?[Q�0�7�*a�<�6��w�B�\��kr" �{�����)�|O9���؊eP�r��J2��耻�3F�������
����_2�D��P�7���(#���?���3r��P�sɝ����q�!��=�Z���
<�Q��ݢr�׏~�@Y��M�[p�/_��NR�IԖ��ʬL�Ԙ�Yܽ�w]��7���4�DٚLdO��VB��f3�8���V��m�<���JRa�;<�H�;W�&�h�%괙[4��T&-^I=�sr_�pN<V�s5siG,��=��Kj���vC#�a�d_f�>����:��5��b���j�f^%v���U# KS�c�c�m#�41u�<����Q�Z��8���U�����#�� r3!�B�ʚ:"�����J���[
��}eN�\M
i�Jۉ$�� �`j`O��A��/��H���z��33"���; ��u�7"���C�B_s,q��w�i���&ċ�
ms˟�0�dڳ7:ʌ�SdG�� �G,�	Q� ���?<�Z�"�<��Te��v�$~�i	�^	�v�%�UQ���iN�X��݋�0��Q�������
�{���/�Vh�떧�^��İybr
c彟a�t'$�{HE}d�r����h:�x�)���<B5���Cr�Q܀�9��Kq��e(��r?߷"����sϿ,����"s �<���Dh�Gj��c
���4OC�^����5_h��o$?_zR˿������q&V�B�8%�d���1�F��ն�� �3LL>�%��!j�0C��»�VcHh�1��뉝f����<���z��D�~-��U��BD��s�1��h��*�������Y�������RM��N��N����Y�Û�����@�E�*��2�
�T���HC$^�0A]yGڮʨHڬ�ݙd��|�[d<��f�g��jlR�Vs�C���u&Ι�!�˯�d^����я�̾�7���d�� �� �c�a��1.�X�,�QG~I�o���\���-r�1�PU�Ϳ�y��t�����C+�`x1��n7��+�`z`��"���X���Nϱ���yV�e ����h 9�������rܞ�E-�t� %4���oTe�L�;��� ȏ7Z�t�q#4?-Wl1>2b� ���m�',5t��`�v�7�H���<��۫Lb���S���5k�����,�����k"%��������Q���ml�Es�������:S���]~��/$j ����T��"���)�����6�}����'⹹�z5c|�Z�O�eF��(�M��� �f��bƏɧpݽ]?&��9y����G�ɦ;������Տ�A�N��l����+ay��s�G�ܚ�ˆ_Gr��f`�̎B�Ne����A�-�S�`6#�0(�����Oӡ�-ߝ\F�:��+`]��#[G�p�}#A����lX���l�h$�QU�8�@Oi�Kv�U�˛�����7��bͯ6���0ݻSiV�mӏY�"FXl�ˬ]��*��o�g=�W����Ͼ�Vy�0��A�음��|�d��P-��H��C�	?�#��^2�:M�C�Ϙ�h�]I���Ⱦ,C�T�ӿ(Oe�`H�.�h�f>/.M��ǩZ��w�M�¸��i�M�c�C��H=�1����^n����NW�� ag@U\�4�|����~��{}Y�_�����"͙�q��V�<��/��q�	�+�|,�W���W�Mu�_p�N-��;�l�I�m�)[x|2Kل���.��U�������J&@��$�]�{�'fY�X�I���$�f�� 5l֘��d����:����/�)	��;v���Z��j��ߤF����K�y�h�A����}��Ӫv~$֜�l���U���F�ؑz;ѳ�%�I�3-�|o g��'��X��~��ŌD�=�1�@P@'@�73�a�l#��ф�k�便����@)5�P�9n��+�j0���&]�P��s�����R�v$P���j Ӱ����-� VZI�l��gDn4��>�E7{���B.Mx���C�x�$�a`�9�{%'G�~�:n -��E욜�B����բ���8�TW`���dK��h  Ѽv����;����fI�p�g�3әw�g~�S���h��t�1��N�mK-��f�,�/f��4���\�� Py�E��;s���ڎ
�0���Gc�{�k���'��f8�\
��`wei/�|�\4OFjw(2(����܏�"A.�OQU1 @��21lFz�_�8����h0�eFa*�_��kRZ"��J֔M��9�sɔ<Z8z��0SXH]e����GB<��@��b�5@�2?/)K9�[��n�ڪ��_V�s�8��{K��2�٬�Ҟja����@�mL��W��/lp�%�L
ܵ�y1���Dݯ�F�W��%�P�qK�v�u?��g���:��W{��b�<��c+��T�IBm��E��V��p���Z�"������J���h�8e?֋,�����F�LK��"��ĝ����ݔTW��4����.ܜ�EiX��Sh�b����RiI>����8�T�faވ��c`*���:p[y[+Fg�A���=aPE�n�d�_���y���ן_��(q�LoT�;� �%��^����ؽ�	yA󣋮0��)�����x5��@<�c�G�7a�Jb>$�~�~����i��I�9=��0�GDә��k\5�Qq����I $�>�����YU�&����?�?�T@�jC_���R��c>�UXM�L��$�W��P]��t�%��m����_�k��c�����e_�7�A9U�7�C���s���Z�=�T�J�~����³�����:�Qs��кISe@$���3\�4��L�ӧ#Yg�*��|��1W����Q��m%�Y���q>��b�̿Ķ�]|�� k����Pc���U��񵥯�M�L=#�����U��#�ԥ���UbI��o䎃�a-?y�<?Q���z�n���@�VN-���]��Z�V`C?#��J���Q7^"��\�2 ^����+.���2�՞�~UwT䳱/�xHq���S	uE]ҌJ�HX�i���ݧ!h�	:5@�-�&_H��@�p��mў���h�R���s�HE��?�*�a?���zG���1����i�����R�,Rn��@���bn��	�E�
O��=�7�8���'�.���6[�L�c�z$��;R�/ �>℻�;���)��������3�Ռ2`��0e���uf&c&���G_I���<A6T�9V��<H$��
�k�� �Ne�/}���A1��1h�|I~�u)p?��nx�U:&�o��i�jb�@��?������8׵�z���5��%�I@�p!Du���T������7� �x.���� \n�s��ǉ�v�T�8�a��p"�N�g'��#e^�u�-i�.�9��wL�9��˓J#spE�:�{��T8�';KzA��p�ع/�F��0:SI��̿j�/
C��r�a]���&Ri�ۍbڠ��9�������YD���e�"��%?��j9�E�!��i��ga�յJ?��c������W���{�<���t�=��}*�]yЍ�� �H͂O<p�,���F){���_Jȏ�|�+�V����;
n�ƝAxs�p�=h�%gB��y^I]4-������Xd�O4O�c9^��a}��F�ە���M�*[o;����m�FlnS��
�&Գ�GB,��UcI�|0����~b�)#|�s��)��y�":�wYZOc�I�B�<�̘��Zf���z�\1>.1�g�(7e_s����JfNT6w���������;o3�)ߋ ʀm��(럒b�<��O��[%��{5D@��Ǭ���S��˱�
����!�]��b�=^w�Ϳ�Y���O�"��j�U��#���st�e~4���$�g
p�^/�MR^i٥�$�ML~��'I�[)zs�f<��w��m��\m�zd��I�.�����DΓ� �jK���'���ΟBoE���� 3��x��dV�]�A��b$�Z�/�ф-Rs�Tw�W:���@XQ�5�u��ן�և��{���v%>�>�Nq�y��N���8�]����?:Ih� j�%�&�b}M����AP�|w���S�=R�v�Š^$=����;��0�q�2ӦB9�i��Z}e1S{Z�zF;k��{�F�i����õ��磳��������AxĉF��k�mq;�/
@�n[���N2���Z�Q��V����q �~;k5��[���ό=����\1�I��e�b�kМŰ��)��-K�e{��12X{����	�w�ڝ�[#�?iTvǡ`!ѕВ4o]ג����=�m=�.�9��~B唻����,�"A�h�a����JP�I�Y�B��/":��F�)�f>��8Zݩn����S�&��8��z�CjL,��o�K�fM��@�ykbZx|>�jw����l�я\��Մ0o#qN^���:���{�C��M�Ȕ��AZ�I���)u�j��ؾw�
�w��䡙��H'�����e��TS�n~���N&�J��K�?E:�����+�$��p�&I���jݿ�с�,�u0�~�.�
�n�(�9!�	0��-�f��I�<S0H| ;;ǲ6 ��y����AS]z���"�`}P���Ȏ:��L(	��4:��d	�||��":{D�~���Edxʊ�zْ�=�y��'5�	p�*=f��ʴ%�<�:*�(�=����D��ջ�������Z��U*�ݻ���f�]3���_?�/in+W%���%����k-�Z��&ύ~�S�5C�ejv�(L4����$�Qk��p�G(��Dn�����Fמ�%���EJl�M`
J�|is��|e	7�`�SMf�%^���kY�(k�@m�{�uC׎6uN���Q�@ �5Pb��Ջ�2�1U����Qq�e����E�m��y���v�G.�0ܹ�<��5��B�MP�+�4%�S2��G���<	��1χ$Eh��e#�e	�E��Y��e�k'1�w��c����[�$�ڪ�I������z��T��j�s�x��)s�����T\����?�<�O+U42��|��6��`D�;��v��6Fs�o����YN㞱�7�4BV�b�		d;�n]?�3�=�z�Ti�u�&5$S1�ߝ8Ji�x�r\���B|��1�5(�x5���_�:ۋ��T7��/N�w5R[j���H	�O~\��ײ��p�جu�t�r��Zʛ��p��dU�p�\`Ϥ�Kf����O� h9iֽ��")�F����R�.38������LV�9�!W���<З���o53G��*�=I(o�I8��Μ����~L�`�}0�^X�LF�L 0��|��N�j�ya�"��C��sc�|i�P:Q���o���-i���p�'��z*���f徹c5¦]�f>���İ�ނ�6@�V��bM���t���`�J<���<�Zw	�д68��������g��?>�����P�ŕ��0ϕ����4j����@O7^�!ѫu6W �`���D��5��f�viź�]�IU�{5K���\i�:�0:�uSz�>�����9����l&�m��v5,����ayij{���ސ��n�^h�[wU�aY)���`��y*�]��!�8�e�1)j;���g9\���Q�%�CO�i���b�cB��&�n���.��}؞"��%ρ,r��5�Ɍ��K_�D��!�.4���!��J_��a;��es���W�kIw��~���jw	�l��7'P�H�������.K��h����$*b	�����.�S�:|#�`�������h5��"E'�R2&*<�:N7ק��w���̀���jgC����.o(=�%~�j:��/�h��ުĴw�iT:�9�C� fcB��JҎ�=� �]�b�T�d`$Z�y��[�Z
�T�'oF=���\Ø�,X.�*���k+:��M��;Y���nt��t�d��A���)�}b_�1F%�7�es�v���B=�,;A��2T�`�pAu�'u	c���zr�;z�-�ׂ�Ϡۉ�$�9S�6G���V���ƀh�J%�5�2�N��i��${l� ��;HDT'��U)H��� �Rl(�G�pF�v\�z��q��E_�S���ϟ}�"�����Ĭv�0a�bkz�bS�7Aُg��	�թ��$�L��>\�G~m2��/���CY��T���l�郻3�Ӆ)�N㓴	cR5?J�)��q��v�62hRG`o���h���T��]^����dU���$��=�����yt*��W��/����B5�;W=�·,��BX�2]R$���M瘧@�_�Æ�,�6G��\��R0�}�lR��rڽ����r8�|$�'�������W9����n�U�X�]%�5���C,[�y����g�?q�`@nl}��~��˕�ЃNsՁ�N6
7�N����>s��E�SY~Ic�	V���	
�jO�6�Y�"Tu���\�½�i�8�'`$��%'��\�Ħ3@�k�-��6j�V0 � F2h�j�yCUԷ��@��{s���A�?~6�##5(�g.U�s�OR�;�9��V�̸�Jq����q��B.r�+�'S�Ѯ1mK\�"@�믇�oj��3�?a�G|<�I'�Vd���V�!
�� =���W�}��$�Lf{�<�����lE�M��(%:#��Ks��4�릗Q�{˶��g����,]��D�#�{�L`�#)/����d7�C&�j�D��Z�n-�#|�5���ۗC#V��_���v�W/��W�}"��a�+/~'�~e�[�IE�p�h;�#fY\Z��-Zx�򰍏��;�ϙ�)��������ou!
!���o�F�1��UK��|Rxt��	!z������vHk(_/��S�ȕ�S❇,;��%���.7��!��BV�U��uQ�3�}#��)@��b�k����@�B�?��Cn���~����˟֩P�2Խ'F��(�Q+�|���(DF[����u+q6�6j/ �W��
��b���(�T����lT�9B�^���ʛ��Dj����ܻ|nO�GZ�m�G>�F��X�^�[
>NnF�X��5t>����ţ�.�?v�s��`���&�l�ĩ�j��xM�GW�ָ�I�6-�W�]��u&�ZP��-�5?� 3���Z�X	��'.����0�dթ��ѩ�Rͮ����9��w�X�0�"��[O��L���d^�t�E0�q� ��G[pU�h���3[ ��	*���p�rT���蝃l�z�AeLs�0���{��ϳ����W[Z�Ew3N�'�H:��͜��
v"�Y=��+$���4O@��:��($��c]tQ�A����zM�vK��U$x	K�:�X]� d��v�֪&��K>}�x_]��zj��ү[������;Y�|�)� �nѨ��Nt8&	m) ��BT�z�Ŵb1��R���yi0~`Ħl���7f���.���k��ngj��GS��W\v���z�������@��a�ÚT�<�X5�lC�"wLӷ�r��d�zZ�&22���ZL*a�����e���m;c���v-hzJG�����ఴ�n��L;���b3 ͜Nf��7a�&!��@�[Z�U��f3��p��-� \vv_[r��B�j_���2��P
0�������A�𿁘_��m�I�ԅW�Jp��8Go@Rqۚm j
�zȒG�؃j"�B�+�B��\�b��e���ھ�ׂ`ɑ&ѿ�+5��vV1�Մ[$w���l��Z/!�S�Հ:D�xMQ��#7�������@J�������%�����"�8�*��9�ʔJe<,���ػ �f���~/.Gê{?�H�.L��Jv�sb7�!�J��A�}C����e�KJ!8,t��o k��I�i�;-m���8'���c���tz���[��P�b<������q<KK�(ԧJ��kq����Os�nb��HU>�7��q�Q?ثP��E0�?�oI\ó�]�;��[��'�Y|EZ?��7SI��ʊ�?no 7�t~�73%LC��� �v5�i��u�TM �G E}��Z�����tRB�̌P�g��_1�Q|Mb�����%*�^-�Cu�Z��`��hi��D<����|P!%�~��$��w�,�����O c~�ч����.D/���&�z3�,1�:eTM<�Z�;�爼�K��w_�l�8
sgb��K��ǜ�m�� �&��j��+�-�6��2JT�w��s~��V�D~�bre�W�ң���?�$O\�c觽�I�%�l��u� ��Y~l�#�e'y�ol"v��{��c�PwX�VnP�g�5,~_�����E/��l:Y)%�yjT��?=��k�f�e$�f��lL6nY�}±�{�rM�[�砷�u,&�#����w�H����]�^���ƙ^�pyq�.s6nbpo�N<��,����x*�}�!�p�lD�����u�q|�2MZ�fҿ��~�WQ��6���n�4�$�_o�B�G���@���IK��_�̿T�ܸ�pzu<�0+�~�+�ނ�~.�,�3�$�$x�h+���&q�n�.� 7sªџ���pskHI�1H�ɟ��{�f
���7$�jù^�TD�Y;+��fb��Ӷ=G��7�Z)���l!Z
8Aősa�JEP�KK�
����N�"SU�N����Z�r�բB��H�:��坮g6�˫&����n�i���1��L����|*�5�����R��gWI�P��٠� :��;eic���u���<���眸M��.6lE�?B��@!{?t�����H��FU�R�&�8h|��W�c���9e[��f�O��1�[����r���`j8�Fs���ӯ�ʽ�l3�\�'iw�r��<3�hI>%��6,ny�9�	�~�?��x�7&�n��퐂���¶See �����.��g]�"'��P���2�Y�j�~�@��qM"K�D��4�ɛ�#�a_;B h���q)���YFi!���.�{������^�txjp���s`51/H�U)V��u��w���8M=0ŭhw���H�&�7�T�A�P����ߡ(N/rBW���MA֙��gu{@O��h*��F�W��!T+_�!�>�K��;M��+��� �w�����C��_IO�#�������o*?$Sw9�$7E����VH��6��ѯ�!�����~��jya�h����!�3�gE��(b��oy��}9dB* ���oS��y��uruʋ}��ko�/�d�������^XY �(Ue�hC�t[��$���S��Y{�ԡ�.g ��Ԩl�ui�fB���r8�E��U�W�PO4��!�+!mS,Qo.$��p7�C_��'���^�ȕ�@�(|N!�����#�!����j	�J+Q�?�7g�Ū?��������]���1^��uG[�8"f�H�=j�.˭�<�h^�K��Je�Imo�+/�n�����Q��yO�ͪh�HDv�w<�'A7���+�m �k�v-;�(�2ԛ.Y�)s�*y�96�6�:5�?@�R�"O�L����Q�=g�Rt�����_<ٮ���h'.��S��������I�POD愠��@h/t��j�t*I��VrZ&���� =��H���>��G��Z�>�=}HnT��kO�y��'�<�z׭��R+�F����<#evh�����͵R�|����hB4�0���gጉ�:�]�������܎{��[��(�����W�˲Ŝx��pPXP�ҺB��C@��"Ei~�x��r(�>}/������������H�����@yG��5��)G��������q����;�nb�b���&�~za�N{�*lw��!��k|Xb�bo)@-���r�H!40Cĉ��d[�S3�cl���Q��R��*���2+����\),ܪ�$F'��ҵ_!��}�(w��鷣U�d��a0���׽��w���K��sFd�o��\S���K��\k|�&�I=-Vg}�H��rl�<Ĥ��kCc�َu}}��1�!ArQ�ZAR��??E����r2�`&�~�P*C��ў���׬�ms�@sץfq�~�������}�BQ�t���xŮ��`%��Z�-Oɧ`��K�s�("�U{��qhS��
-��0���.UU-��`���b�[x
2s�~yW6]:�k�ǞO6~ro��쫪�P��`~�	�"ɝ0y�ˑO|i����r��B�2H�� &�`���c���	�-�8�^�˗��J�e� �oI��+���JwR��Kh��}^�9�^glU�/��_!�X�K�Ґ�5]{���e`W��Nߍ���+S�dV�ZC.��/+n����yvُ�a�&ff$�7�|�_g/^(�-���P|C��=�˫�!/�l"�Ăscu��lU��	��3�A�l�H�&��H�\.����]�t �Z������\�B� A9~#,�㵾S�+D��䔗9�X�Q�/�WR-0ƪ�Ĝ�ҝ��Eɂ\N�ᾔ����ki�G�[����&bmc�hK�?����:�o�>�/��\��;=䀴8�#jQ3ڌO�$��2�3�#��@'�Z%xv\�����0��_���`��{���_���7�{ސ����2��Cq;�#6޶8=g�-�����M�F�'�X��-�a�h�86p2��%b��J�V��-�ý�X�a���J��RB(� �K��eD��䜽8"<���8n��4~�*�L̂5{�{6G��d-�Z2VnE6/Թ8���DՄs;��l9��±�x�8N��9
�}�Ϲ��I�M�v<<�$���q�Q���P�0��(�Ā3?�b�<������~�˚��uV۳|n��1�k�n���l���G`]��rn��J����OӘ6@xc'!F�^5��FF�;����@��'�i[�}[\dh����G�K1�Q�2����,��#:�l�ln�EL�0�"�� �'�\��w]�K�L����f�N�Wg���_�7g��3;(��~��{�+�f�2�Y��Ah�|�v
$�Bx�x�vn,pi�S+�ݢIka��[������-q��6�D�d�t�-�b���*�s8/��Q���O�ߜ[���?~��^gT%��}�x�<	�5�B��N"�{|3����%@�`��b:�tX'^2����Z�o����N�{���/�򃰤�sƑ�{�7y*Ck�,�ɢ�N�,�1&Vb��"W�R}��$�@
ȁ�����-�L�����th1�f��jC�z1TU�	��U�c��$��OQ���Wإ��D���ny��ፕ�r���P�\��%���ub��x	��/��⿡�>�e�k��a�>�������2n8Y��m�y�N �J{�4�@�9�և_N{��Ŗ/cn%��+X��a8���j����Zheq��!�@B�k�(D����M���5��s�pVp�&��7�T%&������ʧ�����!?$t�"��2�Q@c�����s���D��AŐPQJɖJ�kPf�9�8�aEm%:t��z��OŐ�W#�P����I�i3z�D/^��-OP�쁊[!O-۵���@h��k��y��������{tTځK��I{��#�3}-?�k#�e2=e�Q�a�_��z�s�OV	#|���/�֝C#�̻~�ƚW �;��0�W�xf*^Y� >9���ؕ��/��J�_������(�?��K�^z�5ԛ3z1�x�;r�L8d�+*7���x؏�"r>C��;/eIw�Fx��	���ڹs$Tme�c�{i-G˴�s�)���չ�2����D ش��|b�Xɢ���{t �|x�3G.�1�_K�����KeZ�M;O�1K=B����c)�K��)�ύ�X����i!����u)f�60���2�7����Zkp�H�_�vGVcsS��ۛL���4�t(�v�����4�$�[#�<O�Ӕ�M>�G���bk����]��L�?��p�g5X��~��<�!�+�+~�+Q	
�PCM�Z6|{�fU��J�+%w.'Ս�9P��A�y�-9��! x��g�����U�Jld�bC�`xuw��3�#����eI9�ɏ���"Ѵ*]C���	${��̠�\�3O���|������*�r���e0<Z��,�9y��2wO`��DlDT_�z��k|��Ϳ0a�K�f
zpY������w�b��X�V畨/�}�v��&Lb0���'��;�B������Z�#���Or�͘
@�*_�R�P�SЯt�QW��o͓f�f���Ů�I.I.�]A%n��H1��1�D��̧��J*:.�����;��IxP��Ù5�,o��������j,�*%O�^���p15s��70u�X�~��� K�<k����x��
b�L"�:ZhrH���F�����F����:��&3��` i�?f���wO��M�<G�OO	&�n�W�KR��}O���Ԫ��0���1:L��ݤ!�A����"k�f<k�����ug9��Iw�[��n�4.go߀ȷ�"��	�XU�o�'�tu���%fw9)O�?�����m��j�T	�X���X�N�T��
2,E�wrj��v�έ�	�6��O��S��B9z3��e�<?�.�jr�������`*�f4��Tߙ; `���<xj�5�ׇHBp�+t"1�2~�a��I��,�j,�Ɩ�E�QC.�'0�*���X���넌��4�K�=Qn%P6���b^2�<��� +cu2߮S�-1��"���Kgp'�d��+�"O���k	��4�[R�0!���Tr�gy���3�N��Z�!�6�&��"������Σ��#-ƪ㓮W:�����8� 1�����S��y#So�f�_��Ӝ��BbJ&���c��mkd^D3��ƿ;�\���~�e��rT�Lت�*P[�I�Gd��q/�����/����zA��>�)���	1�.��\jW$�PI�g��m�I�sx�$�<���J�^q������D������ �ډ��K��{9gfQefְ\Gh��M����~<�Zs��l_x�R�
"V��"gҙ�q1-{���Z\K��
CY���n�Fn*��%|��i4t���ھq(�o���_�)�[StD5g��� �r�U����cqҧ��Q��&vz��D�-|%R��,��o�,���11�ؠ��`*��y1֮��b���̿B��@��o���/'�r��1Y��N|e��|��F:�盎����mjʇ�|X9N�?V&��{`$?��T䋕P�ڙ��%�@�Ni��.آ*�'����g��1�[�a,�2�8x>溔����G|��qD��/X<?��>;PY��bW����+��J��]FX�~�`��d�y:"�f����<-�M��C�`Ȟ��,u�G������7EI폠=��-�
D�1+0Uܫ��n��2����2���ʙkD_�!E�6n����3�oJ)��˶�Q<����Ku�R�e�vE��;�@bWJo��Wn� ��!�m�Y�d���B�z�`���ج�b���?�x�O���U���7���8#}�v1�w��q�wQ�{��v�,��^9g�U� W����~���W	5K>F$���=[��b(�p.���ʙ�d��c��VN��!P�f�Y�p�0�P�_�`��j���K���*�y�33�R�-��*� �9����z2m4���[_:��hN�4�Yŷ��*�s���6�0�y�H�k���׳b�Oؼ��D�&�x�+�43���������`UޓZ����t�ߗ��>�Mϵ�B'�TL	^.b�'��|U!�'w���g����I��)����������p��B�,�Wa�1fhF�KtL�?8Z?XE�R���Q�:�K�W�A��T5vX��y	��d�(ocl�Ǭ�q��i��2�,�{�J6�A��f�#��z�B0��L��x�hlg�����E�$�Ͷ��~���~��5˺�vO�v;{K#���+����qmb�]��h(�O��(�������_~�}��:&�F���	��20cӍ���r�'Fo�y�?6��`d��	��Z1t�����a��\Q��J�u�JD"OG��Y�M�?�׍0M��6��z�m����-�0�]+Y��%�p�\o)�_S�yP�	 C��� M���m@H����� �H~�J40�ށ�W��q��v�-���lU^����]�dh7`81��CÖ�e���e��V�|�yu���;�4���/�yEn�.m��~"��5ٙ1��:5�B�������:�:�Uɜ���M%q-pM`���u^�`8���SA^����ѕ��F�lA���R6�����̀�+����R�=���;�"�;���9�#����q��˪
1><q�H�\~P����'m]�"'���6ř���Y"�����R�
T<����z:? �1}h�����B&tB�Ē���@��Q�>nZ�O�)a�f-�Ӷ��_G�B���Ec����RKO���֗�����쀌��fgos(7�~��b³��� io߸Y��P�F��Ob���g��P�Z��}�M9U�� ����:p��q�6?�VVG�A��d��^��������MX��tv�G��(%ޞ�����G����ר0�w�,��f	(���R�i��ϰ���B?;�ųj�ʲ�*/��>;у��ɱ#dD�:2_�&�N�yo�/�"[D��D��DO����Y�wLт�/��g�IL��װ~�c���EW�,e�b�	$O�/�K�?��9�xn���!�,��I��% �:U�k�O9#��'ǌA7oNI$���vi<N������ā-��S�xG�^ք��,�������+V��s5�� <i��e� �z��]�ȡDk�ƌfa���1S�6T���My����3��|r�/,���I!Ү~��f���=���	�T��l�d�
*Eb���&ڵr��`�IN�MN}v�!]/�8nb���89{��R�����@p�`L
��%���	�����&\�Z��gF.�����~I~�p���ʜ�_��"^���#��p'��C�����Cw���qA���kC},STT�1�rL㘣8!Rp=6�lf�4�;l�c׊:�J�Q��
�2�#��.����P��������ODO���N��w�;�+<~\��:�0�)Ef����O�O�_	U�¯n��c�}�"���w��:����;]����=�e5/���W_�ܰ���+<2�� �ۘ��:�W�y�^g)�{��=u�A1��NQt�Й5��ۗ�I���Gr��}�$�Vm���O�����1`�)�L����ƫ��IN{Ef[M���7Am�2���v,��\㊴�<v�(b3Y���s�%f<��a�zq�&E�t���*��:aP��•�i W4I�Ff$>hc����w�+���Y���RW�M��{��F�w�e�Urмu���EU*�zr䭳�I�Zt�"�E�I$��ߔ)�F0X�( ���{����F���5-4���*�q��ٻEN�x�V���� ��aqn:q�T��<p�M;��Wx�Ԯ��^^��7|�ք��(�I�?,�������$���26�c���H-��'��l�o�����Wr��"�������^*S�*�B�L�@h�{�c��%�@�>�[���K��i�r��ޡ�w�v�J7���;��(�l�̔�2�1�vu6e��(j`��q��x��XܲAq{(j����C[P�� �������d:�_Q�t��Y[C�3v�xY`aK?<�R�saH��tt~�!�2 -�����g��a[��w_�D��h�n�a��ն�f͚	�����N��ޗ6,!J�"X��C�)i���|�� ��ءb�$�l$@�M���#�RKx���Z�#�Z&F�������[~���pS�C�!���?mQ������;�O�P���O�l��6٠�+�r���k-z媣r6�Bh҅E:۞����+�?)�է�.�"b�+]E�KZ ���w��0��w�v���Ɲ����v�A��q�Ѹ��ٮ6ɢ�pZ~F�Y@M���c^{:�r�M�r���nL��7�ӭ3�Я)��m-�?2�{k��Lj�ه1�� �<��gpMA�wM[��J���M!S5^��0dZM���̀���"�X7��&omu3�׹ ٶ�0:M�R9�r*���~�}�l�˻������z�(�=����31b)�@Y��5rmR��5/��;����t�6��*�������͆KX'�,�>E1�������y7h�����4
qhі�V�����:��c�
��L�n(��G�Z�1A��mm�r��U����?D�^�4����]#P��i��S�C+��[a�W�UwY�w��U$�f���D^��",h��@�\���$��G'�-Dy$.u;^�Ī��u�55D�2A�'<�k�ǃ�Q�(�]e�Mo����] O��.]�+����3C�b����
�Rj�lGs���逖 ����5w}��ٷ��h��)H����5����͑���ʹ�AM�aU�9:�Az����/�s_-��}�M^�S	�o�M���*��e_Q��]FM��
��TN�J�\��%���>됼�����_b�[80�b�)���ͩG��Fx�uKS�!���5����}�������u��i۰D%��{%���]���<�����mAL���D$��� �������[�A⍌)M�b�$!D&���b#�Y��^����|<�MH C_��k6��h`-�7lǀ�J�8ό'�u3:�U)�\u䬾�"��ѧnO�%	�l�2�@E����MI�}�
џ�@h��U7����u�^g3�Ns/�Mڈ���Ͻ^��b�G�3�P������+̃fV��z�L�a�k)��9�t82J�Se��� �z�]���0fo�մ�cS�I �H��&ق�n����&��zϠ�4���k��$��e��i��+�\�bˇ$ӏ���.WlB�^��_�y"����˩��C*����zV��`�&p��X�䰝-mlۏ�-3�ډ��S�|n���,6��X9�D�=!C����[~���˛����j��Y��X����a@
W������ٱF..�_�K�����wO�4"#��wي�X�ݫ2���%S�:@2���A����3]�P����{�����A�ox�oI�Ɯ��"��މP�9Gy�V��2��s1
Q~�"�3����]��[����+�k	�s�XH@�6�������C��"J�:��|Fm�F���X:tuv%�/�Y;c�7�]�A��bp*%<N-��P~�������M}�Y��[uj��WB)�a��r;t�J���Y�v��o^�̠���J�'�|+ʖ� ,��"�Ҿ[���==6��@���ٸ&8z]Pb�:X���!3��Cf�u�`�ԽӋ�q�0W�O��F�o��s�ţ�s�)���$�G-���B�z2��z&	8q�l��;��de>���z�n��0dd���-��}	���\D���E�H��^\���eHy����0Fg�xL�`(.u#<#i�Â�N�����=ep��
�^S�����
�ҥ�b�'f}�tI��������|78�7���zD���@=�A��՗r����9�s&�~���rzl;�!��?�MR�:W���
ׂ�Z��۾�>c9?K������n���$;6�1� �,V�W6
T��>����X�x*�Z��v�g�wګ�z%� @D�܈�D���YE���(��y]��+���{<��ep,�}nr��M{1�(�����?�7�}R�ʬ�b�%kÌ�jhg�;�%�w�G�:�Q�Q��ҿ�������X�����Զ&[��^X���ϤמP)L����S	x�+�����L�`8X��x��	a����.�1ǋ��0��W{���Q`:��/j#-�OF3
R�@���e�:6u�� ��Ŋ)h�Hh�G��H*X=$#��߅ñ "l9<Z��F8��P~�
ѩ�q`�&x8�	/�2��*���J;��t���G�����;a�>=���}P)y,a���d��qY�[�ُk}�Ғ(����
p:��X��`T����
��%�ߦ�z���8�<�F�j_���Z0�E�(��[��.j��w
������a1˵+�	K��H=��xk�n��я��d-��E)� ��7������!r[z�^�$;�e����I86��h�t�EggB]��S�{"��\�j����?*Uq���Cwǜ@�y��ـ�q��g���=.6e�����MZ.K]
:n��%�P�^1`�ǟ�$�b+��8�̛�0��~ߪ����Wױ�P�20�q��Cv�- +���1P��dYW���\k�Z���0�ywt�p<)�YE�,h�i�ƢF���ߒZ�c��������ꆿ�(!3�5��ܜE��I�(F�3�X��s���*��n����AHΓ��	�Լ�#���\���iH���i�^l/�[���d%���FG��[PYN������`'��U�Z�%ˢU������R�2��1�~2�p1|�g`.��N9Q5���_b	��=g/��"�.-%_��*`�T}�82ʾ��=L�ts�fiDe��[3�	��s*p�Xi��o�^���)���7��ֱ����2?�eQI����\&Qշ���~?���W�����|#��
O'����n��
`��$�@�]��c_�Da8�ns�[��w�����Lb���:��� \'��T�Z��BM���0f�A8uZٝ�\�J�7��G~F�8	���W�uQ%@�~��m����7��ۉ����[��TE)�X� :��ͼ����;�d?��$-�,���B\T�Lo��b�V��M��u�p��tE�\%�� z�Y����7�YI�(�����h�G��t��%UB��ȗo!:}��^ _P������',	�0]�E4�ԖLX�����>O��OT��{�"=���_�&&�q
�x�� n�+;ֆ�����rʽ�ϖ �jս���}A��e�]�ç�����i,,C�qiO��}�eS͋�y��U�V|c�2؛��Jf��	(�Y'�lpj��]d6��< �V����=p��T��eڱ�8�E�k�Q��xg#��%�e7�l�u�;�'R���e��L�C>�����.ѲVBٿ�wHS��R�+[g����`_��&9�8���h떳\X��N��9���=��ʣ�+/��t��&�[�{lPA��g��?Ý�j��{��#���L�#+��(�2��q�,l��,U���z��݋2�_J��Ǽ����`Y�Ü��e�&�ǙᲵ�P������<�ׁEɈ�ēҊ�K�0�8�0�<�2���H�F͹��Pt�Ne�y:� K]��t��f<�i*B��p' !eL���G��aI�A ia���ܥ�P% �w�S*o^N�
���rv,��J���-����������_�n�^-���A�j	����!f3l��.��`���� �s�0dܥ��@%�B���9��6�g����= ��"Q�[��T�T�b�m���艄��F:}�(vY��C��{���e�B������2����H���}X{�C��( �o�Z�F5XkQT��͒o��Mx� A�T��q�Z(DU�:p�r/�ӣ��Y#d�'6a�u����3 lb��ׯq��i���BL`��˹���V��}�����D�X/��?|o_t޽��A�R-��S��a3����DYjm���(-p�L�Ẫ��k��B[��0��r�B"tL[���$]�H��0$U6�&5Z\�~Ӣ�K�6a�!_���i3�L�P�=s2�Ȼ����M]��]�H�$y;�=ǉ�}���1��|� TN��O�lA��7� ��e8]LNE�̏�.�i�T���$�9Gu�|���X�P�.vaO["���k�a����|I��!`b[i��>��|:/�Ac���AݸRi�N��Έ6�G~����\r�c�ؓ�z����د3�&���-c!���4�H[�B����"t��~B�����O�BK��԰ovm4"��o�U�-80z��[�U�yRA	�@t�I��Do!�Jl�K�]�<��n/8(z�W��u5��ܰ��+��*��I�(�Dx����������ْ�����ނf�w�U�{,[WF�|B4�I Y���T����{|_�RzE*���������yc���a�Kt������R5�C9a�p:�����*�M�8���^�����@6�Ea��.�.�V[N\���f5x-����֯P����u���I:7V�{����Er�(O�{�=�O=y9Ñ��[	zuif�4�g��n�)t3��1{��z�ϒ���C��E����X�~C���%3��K�:�1��呮�:W�o��ŦF�d�� 2�%Ҋ%ϲ�Χ�!��J�x��o�ҾcC0C$G����`j< ӳhq��ּ�jt����c�IT��/�;������D�&|l$E&�YZ`za��@��*�57���x.�8�ؘ�Y(��3���옡?h���@����u�\�G�[��y��d�,�r�L�j�ZT���h�ƛ�D���lJ�ۈ�9�\!r���t4Q��
�7)����-���)9i�	b��o�?W�t��=f)LDw�2�ls8��Et8S)]�Tq۠F��$�C��x������5T%�g$n�H�LD�d\1u�ꀊ����6����5fZ�[�)k.�Hme�0��O (�	g b�"��t�8۴yt ���2���ʵ��A�����Y5��)�`<�Kf����t@��$��~zW��f���ήh/�l�_Ѣn)�0z�S�T����)��-�F}fڱg�׫��cK��e� ��̄���|=,r7���w�nN [H���,��W�0Q.��G�&�ǂ�	����m��[��D*���P�N��Y��|��g|S
[�R��x��~֔�w8�ȿwՓ�����E����@�.�F�ر&:ڬrغ����.Tg*1��sWʊ�2s�h_@�X]!�^4ãr?1�K�<�0f*QAx����H��;�j���C,����30��җӗ�h�_���P�T�� �Jw��=}G8�p�nP��&�j�@��~�<w�۶�b&���������s�OTA�Z�f6������f|���47a������=8R�{�ђT(���*i�������N��[�-b�q�t�s��j��>��JZo|ˑK0_��Z�TP���a�0ތ2�����~�)j:=����rB�2����p�����*3��P �B��Yq_�t���C����Q��E,ĳ`���߃���@��D�HG;��TE]�17�{�h�S:>�_3��0#3��v{	�Zm��G3B�A����L�� !�A�)�YtZ��3JO�>
��r܏�@��XS�^��M'L�c�?�u잍���RFW�ɠ�9�I?��L�����gzЛ��RGF����F���\�K�4a� �ƫ��Ji�?ן��V���Qb�;!��`y(>^ݟ�/ݧ��8%Y��ʱb5a��" xڡ�Qc�"��~��P4��0v���y�3�ӄ�a��6���)F�qi<[4�fQ��x/�\8�]�Z��m\�,�䋯�u�d�欽�=�AtG/�z�S*u��:YΖڃ��Bp��NBVZ��vH��L)��[�5�_�-(��ߦ�x�A����;��a�������� U ���L�5��>��s8oD��6|��s���۩�iŸ0ɩ� ���!��/��rrD��a%%`�r���=wD�	��B N���7�Le�{%%���A���Lh�����B7Hk#;T�
a�TCTޙn��\c�K}���am
;@i>m��jY�<���*.K�5Z};I6��kʨ���s	�L�:��
@t���[����� %$�}A���D�i������W�x�Ә��{I,?6��睢	V���	�@F]� rgM���)α1�>�h���I�>v(ˣ�>r��u� ����4��!�!�A|@�)�0���� ��/ny�y�����K�r�t���#��I�8����Q��`��#��{�������n���^ ����VȒ��Աo�:-��xH1��h�e�]9_��Q@���0!�	'8 ��?hU�\�-�ӘJNׅ��N���o��9!�+풮0��%�4C�h��WTn1��.zl�d}7/�;�K�o�I;����[-!3�ڲ~���LA?���3�k�Ƚ��T蚵�j�s���X�/ �Ȱ�'���նY��� 8Od]�H���6�o�P�w��� �R��x`�./�8h�/�~{g�[�A #�jف-���HϨK@���F�J�$IF�c�]������u)�JQ����g�w�M�� 1l�>���������^�����3^���-��)5%G.����"W��M�/�~��/?V/�)��{�
�T��\~��P���u	;ۣ�W������ ��Hp'�^P$sӽ���Y.`�&��3���xx/�:צ�^���
G~���	Y$�t)�A��dq�$����)�
S8�=��;��Ou�)���N��:�g*)˶�Z����U6� ��1���Q0�Bl�zzdrzX�F�7�}g�<>��H�����џ�P0�G�km�it�����_?�U�x�C5z�u	&@�U:Ͳ�$��}��~��ED�m�`g��,@�H�\W���l`�SNL0a�l�J�C0��h��Jv������khG��yD��M\r�	�$�x�8�6RJ�2^!�� ��bm9���B��I��vB@s����]����y'�����D��R���&�>�ax���~�t��ЩR��@=8~]OvJM�jM�$�ﻍBu�`���aA��AC�Z�(� +��E���>{K����A41N���<|�!��ټ :��U�<�|���K��.r��ܼ�-g�b�}�����׊ne�{s� bS�6��v��'����t��u�ӧR|X�84OA?��od�y�S	�,�5b+�Ѫ{�u�)�v��"�├E��K#9�#s�	�ٱ眚�Q���� �Y�qLϘ����q���l�"}Θ�-rC�-����I�F�<~��ܞ�U�<�Z��85�j��I�T�R�wE��$�c�Հz��i�S)��.�1��!<��03Fvh�3B! 
z��gk<ʰ�"k~U)c�.1'��~�.�+[�RC��Z�M�GUƢ�\���,Ҍѳ�7�:0��~��12A�dh�f��S�G��2�Ct'l��s�/�j���wJ3�H1�2�M[b>���;���]*�j�V��ն��v��@�e��*��9F��\ =���m��`��8������b���6JiL�Ɛ����:�I�)\��Z�pθ[�s��ؘR��	��?������,��6���p�u|��Ib>M��2m�ʬ�]����9����K�iGj�Xk����³�z��2�:XXLɪ�j��/�4�#�J�7zB�0���jOsd��êys���#�������nq��AF ��w�٢2�I�����~����[aƯ��#�{��Iok�5(�,7�T�9��\o�ދ�Q��M���pJ�ss �d
�pH/�ju����m�@{>
Ϛ��,������Qm�<ů���*pH������O	�Ef�^��n"X���+��
�ҔՅ��[�	��6+�Z4&�]��8�0�NaC{$�`��w�� r�1�Է�XC�ǤÀ���C]��RO�	)\Z-v��ԈT~��EEߢ7�p�6��Jf�>{����,�jdݻ���h�����n>�'���T
�:L���P��)�+�Gm���&l��O�b���^��{<�߭4i�ͼْ�y8���n�0��h���,}&��;�z=B� ��B���ڧ��Y��e�������r!>���������7��,���ܶ}��DS��nۭP�9���l;��_�J���x!���)��od%YOMQgݨ�|yB�`#L�؉��y�,{#�Zg)������M����.�@J����"De�g�T��C�D��4eS���!��ӑ�h:��D�ÁJ0�`�Y�>�Z�2獘15��,^އ��Vi�	v!�r�{���[�-+`B&.%��t0	�P�:X�p=?�{}�z��$I���A��=!��(M���{�;h`��Qs���ɇD��W��vf>ܴP�7�ɷ7Q�'��<������~���ص��h<�,(_�����8U_���RV���)Y���8X��Ϣ"�.����)�����+�T��!Ȩ: M^���;Є���cr̤t�a���e�����]	{.�L�e�FZ��&R�s*�����a_i�H߻�#X"���鰱�j	� ��P��aN��X�7�J���V�O~��Q����y|�=.^�
�0M�Ҡ�S2/Z��`�y΍v-xжx{<����V��ͼb��m��P���3�b/���\�� �Q���kŘ��bu�s���P�)a�EY���o����Wj�W����Q�j�UvP�Z�y'�]q��,^cS�v��Њ}c0�}CS0�'s�ͅ/�c`�����Kj�@õ�I(��/�f�A�Z���_͌d�P/����,��Xj�~��A�ܧ��%�Y�����J�3���ѻ�9QИ���R���^s#wm`���-����V9BX)�䞿Z�E��"EǏݽ8�N����{�A�2�1�?���	1l��J��Q����1S�6�
�?� �Ɏs�)֤Yc���/+[���*� /���j����"��ufx!���GD8�@IB ��d�k�ޓEy^.vܹ�{����r����-�]U�����=�<��%��U<S���݅T��fƔ`�G�9@m�KS���"�I�KD1�Y4HH]����S��M8;F�^P+I)XMO˟S�)�����;������	f�*���~M1�6Z�����qo��ș�����oB��)�K���j	�#[q�]6s�l�Z�\�a����ۡ�H^ў'���k)�G��0<��oS�ʘ����y�J^�k�������U�	v��k�/$���b!r��~�<u'�K�㨱��1��8O��p����%aˡ>��fm+�&8{g#����f@Tςf1b	�Ƨ�u�uǯ�[�.����yN�0Q=zj�HJp�t᝽'߯��Z�M��� ��if�Q���Fe���.j�o=��Б��&h�im�
)��ҒG�|���i&y�ߺ��h���0L?۬Q�{h��2�0o4��e���Q�'=M ~�2ښحo����N�/����d���$��G��vIxmwF㭂��#F"�}��JI�R�q[M�%R���Id=���!��A��$��b���Ijl2[RS8wEĎH�%�����,�k�O-�mϥ {M4� ��Υb����ˢ���@Ï�\��>Z�2��c��4���q���9�h�
��a?��Q�ѓ����<�D�de����������6|�h����O[i����h�Yq���୒���,d�o�`T�n����,U�X�M��"���z#~�9�n��{��bN��U��T��HI���:F�_��b88���)���[u�i��)"<��Ʉ��.+��dV����Ⱥ�3�G�� r�2�/���$�]��u��P��2ž9��@�����v�>H�yύ���D|��e�l{	��}B؅��&h��k|��¹r�76�i�)5�̵f9j�Ƒ���X5Fj�����;&G�`/�[�2X^Ķ�� �Gտ�0���SA�(s��8�8"v�W�{}ح���l8(��a\|zҞ��;���Յ��)l�(��gU�G�x���ۺ��֘X�����Q?���i�}1���32���Gw�U�z@���1AA� l?�?=o�%�=���r��gs�;-Y���cW�7�1#�J��&#�c�`���n��d�S����1����R���@��̍"Hf��M��n�h��,(��v��΁{�w,��^����[��/�'R�V�F�<��z5�k-�{�++b 8�ќSh.�S	c���"D���|FH��\��4�T��"�	F�d<*�٠<��A̽�ϯ�~&�笴!�Ŵck ʔz�l�a�8eIք��#+�+���\�r������V��As��6� >�so�~2%;d�h��[� f�iB2D�rⱒ�u���q�nƒ}B��/�Bӧ/m8����,����򕧹��F�/M��b"����#8i4�O��FqT��1��݇n�JWn"Y��>�*�S�P���b�2���<���⛰.��8Gg'��al �s�Q��u��n��34��?O�4�G�=��I�}#viw�`4�N� `�Y(���u=\�^��Fi{^��%6���74����a����?9�{�р��+��*w�|�>w��1S9��y��x�V���B#�
6��&9�3��l���>���/�X"G8z$h��҆��:��q��.[�qu���>�u8� ���fg�v���wԪH}}�p�'��E�WFP�
Rp`��Q`�G�[!���?鎫��	�ڌ�Xj��@�������S�����>h�sTJ�n�y��q4�}�M���([XN��Ν���b	Z��4Z�&O#�Fua�eY}���@��XCS��T�T(	�B-��`�<8\F�.k�0�c���8���a���{��#L���ƥ.O��3��*)�?� �(9���&���@��p:��2�h;U�P5�1����r����ͼnn��N"���΍?�R|�p��������CW|�fr0�¡M[Gm�!����;T�|����{�YXp��p��_"��*�0&Z'�	���tZ���������5oED��zѠ�R�pc �j6������F5ʝ��s�zG��<6J�-��V�}�0ږ�Mx��S��|��i�==nڍ����q�o����Ơe�'W��];�����9��'�����;�ͼ���̮��+�"R�pا����g��&��&�����Չ�i�.)��vvbP{1J�A�z���t@l���&m�}�ByH2�醌�+g�ǐ��S\[�M�Qr��gv���&���ɊB��k�������͑�T5[�f����s�}�w�2������ne@~{�o���54F}E_���E��bX���v|v��%X�������:QS��hN�S+kzGI�@x�]��FP[��^�����NQ�)�%�p���D��C)Of(.k�ۣ$�\��[�DZ<�$�#4 �U�V,�����r��b���|ŭa�Rj,����O�A`R	�R��HS:c�2��Jz��a�����߼���ޏ�>���'��c�պ%����� \؄z��>o�)�n�����11�_����7r�-	�	��������:�֤�p�o�̨�I��b�)�>Ǻ�D�K��A��#(G�SfjU!�� �,#�s�d(�G�R_f%�V��ꯘ/��wT����0F��˿��] z@
&r�L"�X}8� �uQ~������)��O ��Ԩ�I�]w���Z���X	����$��؝�'j��
��툦��H0ȕ۸�p J	A�ڂ��!M��:n(��·�Ai7.FѾ�luq��)��*;64�%�������}��u	�'+���ʨ�_��v\�L>����F��@���\%܄�rQ1���m��;�j�Y3�;�8�,��A�ь�82����Og>��:�����
v�4�}y�\,BU��r)'x�3`j���͸anxUӂǌv�*�
r�РC4����}��x�(�R�=>޷���{u�Ϲ	W��ϕ��7�L��!���,;�SدR�n��Hݕ��H�%�Xz�{���u���?уͪ��A�#��o��(1Qf=q�M�F�K+	#�cˍ�\aJ��#��p���iP/k3��X���"9�<DuyD�%Eq�?�}�P�h��M>�͟#(%���� �Xmg2PRۥ�����fe�J�,��ό����e����"��N��>���"_h<g=�PɁHd���	����Kb+f���JV��D�Z����-�F�vp��m^�Y��ؙ�>~����f�B2SOL��n�vh-
W����\�����*���<����Yd�����1cp�ݘ]�sv{������'��غ�kK�8��������ܫ���%'����]T�!2|S�6V����Ռ���Y�]c�����XyF���BIoݥ�#���7�ۙ�~e�gat-<��7�֐q��rixz=M+�d��(�W�\����Z��ԥ�4d�5o��s&��Ǝ^�g���N$�i-#8��T�z�WVǧ?�(�MD>��~8��.4�%��qU�������p�A�X>l����7?��������">�Zx q�I)Ŀ"�CA�U�Z�z����ӫf��Z�	��T�^ј�5Y��7(ӄsg�m���^�'�O�s�ˊ5w.,ű+�
$�߰��5�p��d_j��Z�䮪V_?��^$�IBJ�û��\��s��`��R�R�*���i�`�N-��u�g׺u���Y��wrTR)Yd��tj�W6BP�	L�n/����R���;;rm��Y3Y����7�f8lyQ�z��؅���`y`�?R���;��V{AW;�^]÷='HWo��ḪVi��-
�@'?���L��
v�w �J��~�:�L��a�߻�F�ۙ�FW��������y���*�#�A�7e�P??�ޘ�zX��gnߑ��U#������/�d����Cn�pA�L����^5}�����j���n籣��C/6���4ݣ+�_����؉�������s��0'
��	l� \
ʆ������]�]�.��f	x)��O�~p pߧOؒ�t�?����1ݤ5��q��f|ra  #���0B0�C��l��� ��DF�W��5�"]��>׺�S��}п���c͖��92H'���[�8۹�z����o�'oL� ����k������7��@j��Lt'f'��e��#{������>������/��>E�6K�M{�̞�D����V��ږ��˟�
�������[���F�X@�-l��K�yW�=B�9]XO_+XpVA]P�6S�*Xo���p����%J�>{�[����LU��X�� 5Yk����+��twT��f��p�Pd#ӫPZ��P�'���9�̚!�Oݺ�6��t7��!Md�o�Hw �w��Y�:�W��>�md�O�JT�њ�1��0x�h�@�s(���B��W��Ԛ����D�}O ��5�k�w�m��H!ө�r9#n�7!�/���T_��hedK8��&C��jn��'d�N�ѻ�W�����ʤ6��N�ȶEs�<�����k��M�w�S�ĝ@9�%tkl��^-�vW�� Dsݗ\5ݹ�U@�pu�a7�06GL�w��k ��n��JnRt��3B�"��q��n�,����E',��x��U�˨������%X'y*E�E�t��!��}���k֒�_(ƕ��\��y��N=��V��?_d����D>���}`��L�Tܙ�2?�_%�=?��b���!�k����1�ȷ�:�,��k�_��I�L;�y2u��q��"�yΦG�;��]��Dw<�� HZ�f<k�v�eč��I[Ku�����om,�ѹ0�R���4g����g��K�-�HC��ć75��о4�!H�F���X�}?O�E�ed����C?s���c�d�U�`�.A�4l�c �n�@�d�طu�;36W سĶ�Ne%"��X��h�P�Q�
sV uں���.�s��TQ7��clkn$1ͯ<>��1�D���8�$I�����@x�؂J���x�=���ʽr_H�m[9�l�W����I� ��p���tX|��Ùx��	�u� ��|v����T�pG	�EgX;;��Ql�܈ӻAX'�bU\��_�&�|'����i���vvo]f����oag���w��j(�����S�o�Fdu��Tuko�7�M�di���uX��~H��� t��oR�U���%�$P��=�lYh�����emPe-0{�Fhv=>��Z�z����ʐoWg��Q�5R�6�]��E9��2N�����T��U���v��F�q�_��[܉1����=F����� D�r+Q���[�8��A���S���6�V���&����责J�vZ*4��-���$N�P_�V�*��[!n��2Չ��>�9DA�cM�.��V�P�/sߴ��W,ؠ[W�ڨ���p�Ct@�|���3�0P�B{C@��o	�&>M�)��T��ڪi6}L���"�9y��
�h�.S�gÈkYtu�����Ӯ�ic��y'�y�~�f(�ؔxMBV օ�ҳ?�s��߉����k���u �ώ,B!5�ݙ�m#���(=�G����Fo���|0=���&������Pśh�҅�n��0��t���M�N��N`�p�#*J�o?��kTz�3��+�,����@e���2G�í��2�ͧ�&�+�W.��=��0��+��*;���%�_��	�;{��<؁�
���=̍�1�n�`�������6Ԣij=��aZ3J"��[��I�����I)H�B��c�UM�b�^�$b�]�37��K_|���&;(>�k���G����n�}
�Q����)��U@aA���E��;c����9����
��tPdƪȎ�7�C��X��qq8a��4� �)�m�7_!��T���)�<��b��3�XV>�\�����-[h�A��3�%�����S�R�'<��d�ta~��uuOC���NS������ʸ�Dg~�>)M_��S\T2�q�-��_[�A^e�},F39��bF �K���w��ã�á�>����V�����͵YZ<K�1/�3� 8ɼ\��r�I��mLO�W�<O]D_� 
�JJ����#2[�$�`�}��k�ooU��? cՠè��3�Ô=�&[0H����i��?����HƱ�:T�A�8>�l������X	O.@��5�9�2�4x9 �R�GeH���ctg8��J�p�%I\
��?��*�MY`~\�T�Ur>M6���w�9r���P:�{l2u�>2+�Z�9�s�Veޮ� �3�!e���V�<���E�d�.�43Q+�� +��p�?��;:
-	�og$u�nH��H-�Ʉ+)�(ɼ�Yn�W���Oʒ�J�D��g�� ��j���SE�Qa�(��#��,�(~�s�����(c#]��-��s��8 �?ٟ�����n_,>r�#�۟��f+D�y0#
�q-w8ݪF�����L��O���cw���6�b��p�k�h�P4�KF��gi�V���Ib=���߸��(���gQyi�LhK�z�6I���F���{�;ǵ9P�
�����T�;8�����.n�,�>|���qO��h�(1��"��^
�O�+�D��EؼA��� ��c���K)��ڲ�M���jJ[�eK�(� �>=�Ω$�:�f�Eyҡ�����HFG�'V���
�dKPyUN���I������d�˂Y��L�X����F�-�)U�̍uM� ����ΐ�MZ�ϴ{�|��a	�X�I�A�l{� ��LM���/����t����P�����b�.���VSp<�'E7%^����k9ia0�����s�����C���/�4��%�:s�XW0J]�$���o]�|���RAax���]�3�ƹ-���e˗x�J�ޠ�L��C{l�H�6�s�i�m�����-+�� %�j['�^X�j��x�`/��/CNxi�;b�F�Y��I�q���H{wmAV)�+���ztV�WL�+�U�gJ*S�(Cl�tnaAU���M�-�Ѹ|5�=��E��#7�P�S�W� u�)�O�c돜� �����h�����'�v�!ruu�z�d|�~�N$)F��=�Y�G����W�����Y��E�oJEa�n9��7y�q���ń�g\})������X _ ���]� *��;_j�Mf`��@KWӉ�s޹>����z��yN�I���.�[�ή"�Tvzp��P����~Gձu*��=}�R;��' Z��Z�@�����rK�F��|��xF�p��5*BEV��Lw�FS�!�ze>�>cc��XҴwΏ��눁�qe�M��a�7�;���[�A<������,��1چ�A~�fθ]RA�n���z�p) �>W��=`��"�v��Z��o{e[WN&��9�l�j|F	ʄ��|���V����J-�^<B���l6~��H?���5����?�u.:\}-�����$K�̕h��P�	Ω�X���2"��KjL���$A�$�����p��lz�+s�R6�>zn�/
����h�����M�FD%�tK����|���邷�e���#0��&|r�ҥ���H���8K��<Y�AY�ıY*��������'�ـ��0����Q $�X�O��]~�@�N�~�����,���3������_��Rg%3�:5ݍ�lx>���~i��0���~Y
gͮ��s<M��������g�2���m�P*��q!9U��A��'@��Yh�	�<���
�J��촢����/���fͅON�CP��8��2��L-�]�X6|��tqZ_P���7�z����e�#C(�"�FXY��t6���������&=| g-��V<w���MӸW#/1*�k��#�P',n�9�)Xu�v���C���k���i��VZѢ)�z{5$l���/-�=��8�	'�m����r!�;UTu�x���o0�<�e��r)�nY�W;������I��*�#wCP��'˽�T0�a(YF�|���������X%���mה�o��᥄8�wZ���_;\�y|8,`��y���&��&Ӑ��l�rZ�R�ilL�^D���>& ��e��<Z7���a3�+�|�vPkh��u�ܴ�.�zlp<�<"����q��2Y̧��.�������&Z2��'�����\�0�˩"�H�(���\��덺�p�n�N4i���#�-�-�Q��%l/	(�Ù�*�L���l"|��[Nn�+��[�v�^���-��Ǡ����H^@��*��� �{�-;��ngEZ�����竔ԅ��Z-w3�qǣ�#x[�bꄞמ1��<67z����>�x�O��K��&FUmW+k�n���%��v�-u�_XK:������������Zy����@�z�w�7�t�Uh)xS�G�f=u�G`S4M�B�����MQ6a���1ᤰ�0�?[L��uCD���M6H)H��o�`�Xc�x
-c�!x �3��h̏�E�:x���ep �sS
f��e<�G:���l�}^�cct�q�U�w0>~�.&<0޴.ȡ9�BZgOMu��y�e���!�i�;����c2�� ���bњW���i�B���/�C�[F��1��϶V#%|��M��u����uI@âP�u7��$�+a�&� ��I=>�*����j�4!αq}ay�pN�yx���K��v�?��G;f$��
��������}���,�\�UD���!�9@$:ӣ�`
��cm2%����h<+�>�ޢ��So�
oI{��1��r�y=	��T苽������k~U���Ds����\Y�}�Lop��ۀ����C���H�� �-3��?+�O'FZ�ŰDQ"{�)�T�xd��a0b2����B��U{�rG��}vׄ�~��2�;ׁ�IY�%��If�sϤ���|�da"��3o2}<$�D��2����S-	�eu��Ѡ�0SD�k\�����t��KpXk�3A�E�g�+�H�(\���u]k��F:�p\�������I��c&��Ba����c��qB�OB\�#��%a�a]T���*�_;>��J�|ʮ��C?�J���n��Ōb&�]�q��y%ftd��-#���U0�����o}Hjf�E�~��J7�4Q���DfPk>��:�tVW`g��G��c�;�SY���*9�����+� �)Dˊ��(��&\�>�Ԯ���C���LV�K��l��z��A+����D&�����τ�����h�R�A�S-n������%��Ń^ë�ڮ�ezõ���fÏ4H��]���g�5l$ӎ�-w5��o��/7�O�	͌Խb$/TKkDa���� ���v�BB�0j�VCE������8�;+dK�F���RV�1�驎�% N�����c��_���Бw��`�xRD����{��Y6�E�VY��V�ę�w�g� t�e�K_�Ԗ�^Z�? g�nd�;�ȥ����*�$��PrQ�v
�)��ԝ���8\�H��cظ.?�p�{MA|BC"'�Ȱst�q�}|�4��O��	�O 7؀f��}�Tk��_�W��$6��Asٙ�ʟ�	������fά�et�R?���f�,
W�5�E��'
���p�&����Ƴ<bZ�Qёu<z�*j1�y�#e�-~��Y��t||Y�������]���vW�':��V��D��T]])�������wC[�`���y���k�I00�#��?5/]7<��i4�i�e�'W��iV��z+�%�u8�����������T���A�|l��qՃ�C�P��p�y4U���3��5���w=��2���@��*i�.���|�&>�`��].EO�אg���� ���(���4�FQ���9�X���>�R1.w�˙d�ben��+�)��&�60��3n�x^ �9�fBœ�,E�������(��+)ȇ@���rSĵk�\{Z���+�Ҳi=����%�o\�|�*,~��	��[{r���_���͘p��|W��0{��˛��H<���J&۪�R��M�-�[�"�#;�M'���7ՍL7j�_�1�;�1����р+�b�Cd>���V]��:��?)�?x��h1�d�6%��x܄���~���]i HO����7��./�ZL�w�=��nS�"�z�Wuz�t�u���_ 8����ҽapV��a[���2���Q�X���B����'�"�b0�xG.���s<� �u3h�[���'��Rk�
ǩ����Z~�=ԟ��6	��p������Q���Yz��K ���UQqνx�>C`�|�t�:�hUn�X��K6o�1����ʅ�y0e9ŕ���͂S6����j��X�}��v�2�_4�x�v�	]���C�U��ܚ�Z��0��
t�����	Ll�����U?5��Q�9̠�i���A���7��y���-5�j[�u����fZ*�ҽ��#Q�C)�S���Y+B�����'	r0��l�	�}�']{�y�������%�ʳcD�8ԡb�:�(a�"���s2Sj[��"r_��d�;L�"c����H�U���*�]��i�!��D	̙�M)pǂ$��JkX7�|3�r���I.�3ī�jĊ>/�/���0�ؽ�XD4�!N���.QhFs�,]���SH�ĉDH��˅Pq=��8���4O�Q���u�~�V`�͍��|0֗ûa���ݸ�U:�栠��D޸��9��G|�H��R�+��(E�O�ah''rsf�<8�	f����c��������1.�����y�\���:ɴ���G�Pڵ�w-a��D���Uָ���3�f�҆�K�����if�h�+�M��D'T&0� V�����9���� �WX��NgzV�un�[j��g�b�a������S���Sz�r������f�R����*`�L;���`TNH*M���v���S�vz��]���5�۞P��u0F�q/��q7	���鑲C�������M�m�� �]��d˛9�I'���f��0{K-�T�[�x�}��~���*�~o���[�Ͳ���'���.d��#�3����Ú�Z��!���
kC�'SU7�J���r�@�i�O,xv)N���,��5��k}p�zܼ��^(�[�nt��tԡ���r�U�꩑	���ŉ��>�I��	�;HR��[h��UΞj �!��O��%
�ߛ,���0�K�t$pr�U��/c)ֲv�rn/S���伜�؉rY�0��>b��s�� 	4�$�QO.��=IzWf�����J)~Bշ"�x�qP��e�@�)�Q�B��{��qi�\���i�;Lc��^Z�lU�9� �Ǒ�j��4�Y1O�s��!�4[�L4u?b��M�q��� ��DɷҪ?m�U�+��{/�Y��.$B��	Y��+6ܟ��Ն&��;4����}�F��i5Ae�Y{ȊZw"}|8;	��Bp����!RӢN�cLZ<hbOdI7�Δ��]X�,��q�{�̇�[�q����WD�E8MU�]A�:�T}s����Y�C�ed��S3�C�N�N����w^��bw.^ѓ�/����Иo�i}/�#mD#u!������CGڶ$aǫ�h9��0��Q����t�5�e�T{�5aM�FI(���E6x���Q�'��Jb���D$v�eYĽ^1�w�w�?�<������}ݟW<2����y��1�*�]����a��?rۘ�T���wMK���q��<I��q��5P�1R�b;��ӱ��b���B8H$�K��d`�֍�\,w��݉TLx�0w]ϱ�TF�,�Z��ew��;�l��ۃ��5�B�S�ɖ�j����V�����Hna�.�z�|���=��1�=A\=x��F��\��G����46 6ͮj�혎��R�s-ض����:�<(�?���*���5لZU?�u��^��iC��`;O<ů�6�@���.7�}�o�<Z�
�j �Wيfr Ji:�����>��uQL='�񚬃��l9FW���d����;��5�����"l	a���B�Ba�nE�5��V%��U,R�s ��LR�����}Y��2x�Y֋M��O�F�t���J��@�����<6#�rw.+:��h�CWNA������Qу�C��c\� �o�AX�w�i{`�+$i�=:�7E��ʅ\cf�[�Q���j'�Z�u��~NpZ����T8L�_k�|7����1]k���œE��@�%��	s��y�C�!'����'tM�=�
���>��Ф�x�C�%�!�F xY���٬�c!皈�͊�F�ƆdX�0�����~��������Nl�zv�� m�[���m�Y�jzX��4�F�o�d^0_�����ld�wX6L@�A�ֲ�T2��3B0�2���'>5���@T�Z�����#iQ�)�;��4`{��sR\M�2J��q�S |x|��,��^ۂ 䇩:̞s���d��d�g��9�+�|-���ʑ������P��P��\W�p]�c8b��zhA��W���u5�.=�(���D�n��7o���)'��Ĉu�h'C���|c7��f!=�~���ez��}G#��t=h��h�a�p����H�=葭"o��8����\��F��[�[�������?))��I��"H.�c	���e�,�I�a$�."jOuY=��)�����n�^����L4Ϳ	=qn��Zy�������	xa���Ui�d�v�d-�1nOY���]��9�-�j��0��S��V�L'�d,����P���bn�n��a���(�B����|L���憺�b�T�7Q�j���ܬ��\WRH��C��\�F6&��i>G����a����a��v�3}��a��-��թ/.VOa�'�o���iY��>�\��ռ���1�>���g�0���Z��9�ɯi��.?��s�d���Qީj��Qs���#�Ϡ� j���h��k+*ܛI�5�����MJ!c[��7���x�̲��@�`�ju��:p�?�k�L��w�uC���ӬZs��;��6=�[5]{�L�e�l�JM��<[�t���HAu�
G;j+6�M�U��R��r�˪���nu˰e�ע���� xR�ko�I_�.c�R2�x���.�6'��s��8��{�؁�8Z���D�۸Ȗ7[B�����v���Kˀe�|ǚ�X>,t��+V.H�+�Z����V��Kq�YxL��O������y�S)o[a��7� uF��Q����9ZU��j�)�9�{�H��|T�l���zV+�? ^��F��f
k&.���,z�zት��;�2O�F��+/�eH۸�Z�[v�F�L��ߞ*����!�7r�ά�|������T�BS�k��w:��sa��`�gd�v�!�EI��ot{c��'e�Mh��s�s��r7F��M��iIM�ʌ�����hbN薲�Z�(�*��L��Q'Ws�����S��f�,?��yR�GZq�1����W�6��^�=��?/^ڠ�������^��àA����l�~u�=���H�P�$��TӒn��H�Ċ�̟�v#�&�ENp��&�)�ݚ���Mf�t�m}rj�g�SIܿ��u������ С,�cϫŖ�Oo�.ui�O{3N�H������١��j93;(�k���`�C��k%Z?sz:w�`=�e�5�r�((TT�F�I�D��MbɣӤ���^<�.~�{*�f���
y���l7��0:���������?�Zz�W5P��L�S��>���pط:ǽ�nXŰ=��e�z ��"Gf& ��~/=��;@�R��)�u�(c1�'N��=ç�Fe)�^�&E}����'n�s�����h�_m��`�ltS�A�q���ԯ<@����恈��sHtwFuT�#*yF�^�N��e����CCC�z�Zƛ���ژ�̏fr��m��M(���1r�H��r6�O5���տ�y���6O�ыT��|�X��b��w�y��"5�����;q��Ѳ*����@��z���mh`]r\$;�=;��,�j���8]���
W�O��wHc������B���(O/?�l's�_����Z\����V�K�C�w�� E�[m�h�K�[RI��r�wa5���Ը����r�}n6��_�u,w�,�Gծ����QB�|a�O�C"��G"Vc��˿�*-���#�{X��U�A��T6�%��5��� �آ�e��F:�����Sъ�����C_��ែ:夻ծ�pͿ=#�"�0�>=�aؤ
�^e{��D���|D?�s�B�@6�O��1Ɯ'R4�')v��0 6׾�G��Km��e�Z(�z.Ϊm
1 �P�@�Z膳o����:���#����)w���d2Jz��l�O$�� �9���N_��0
L"��2͈I�Z�8�:l=�~���:w��RI#�����ASj�����URb��7"N�W�Zj�H�"/�n"�{*�X_�I��-��6Y9B���Z�E"~U�
"l�n.oP��,J�'9b)cʇ��s'
mK� ����s�i|���IDM"�i������~f8*R�_�����)���y��a�Nz�?�6b��Y�A'���Ȉ�S���[�~'�(�-�I���D6:s$��^�$S51����&���Y*�hՍ&���Ӹ˳���/6�R�Äa�w��5�������~��=:R��*�Lb��"g4Sp��)��� ������Yz�F<�VE���h��a�nCd�H�f'�*ipPwQs�9L��*�T@��z(�=*Is�@���6����bV��[��Tm�$��X��ӂ�_�p��Fj�^���$�}�#�A��Mj�X�lAj�'��cR�V(���5=��*J�jx�yn&�O
v	 �cj���?�)4�q#p��Q}f+�,^�ؗ��Xs������|���Ը�&|��>�{�f]*{��2ɢ�f0H5y�D/��R&�k�~f���Ę<�<<�<Tް��p�6�q�-b��0+�X�$v�o<G�/p$=.lͧ�7�iB�V,�=K��������ͣ�D�B}_[�~�M�rj�p���M���3�Є�z�޹�("Fk$�?��j�2�@;���&.�����@�oZ��
���E�p�m��� T�Ief
@eNo�܄�T�?�e5D��N�.��8ڧh��.��-)�e^���4��M!ߋ��:
Ȁ�	WZe�:�A�-R��dlܞ&n^^v�&���޽��?�Y�LgZA�Ͻ^8%Z[R���)�ʻ�v�Bj��Z� v�{�fk�m|���$��,w�?����T�Z.�3W[z+{15;G��#�zO�u�S���f�X��ӧ���l7H/v���^������~3��y���O��QC��͡r�p�Q��B��S�S֚���E��h���v���a�;=�Q	�t�,Qi9���n�����A(�f$�������@,�16�_��f���&x�x�Cƞ��	��{��7�X��XhT&a�_EU��N0�
�(��/PL�C���F�!��dTvK�Jy̽$����
�)����zG�����c*I1s�U<S)��l�{�Z��o�(�\�ذ�,!��h~FDz�@R��!�7�{�����b}َ'��o��v�v�ݺ3��&^ҧ�K�)�R&5=UfY�0j1`�Ӿ4zɾ�+"���T���[;4M���;�m���p[�<A�5kff{��fą�SN���ƣ�w�$=.)�� )T�X���%���}�I�[
�~��]o��T�nY5�ߋ�֍f=�'h�)�����u�
i-�>�3R.�y�^��$N/�40�uK!+h�t%���t߃�d��D� *k����c
#$�H�y$������SA���!Kb�^88��'�M/k�!�����u�W�\�����k� �k����aآ�U�f��o�q��٘��|U�P���RZ C���tCd�Œ��[��WG;����h�)+��1;���\@��ꔘ�åe��L?��6���2��Ӝ�ҫe�e�fφL���5�]M"�tM��O�������v�Z,�P+p�V� g����4?�rl�����O�����Ĺ��)���|�V�˰�����|F��B�QXm�l��%k����"����W��,9���EG���eѓA���b�����L���%=5��R�%^�V�v�H����?9E�A�c4M eȲ���'N0q�O����Ð^_�`�E2%S�orn��C��.���!�����_��W��/��O�q.��~zp=�>��cDC*o���OL�%J4�}��tn�X��е�Ğv+�D���*�ڝb|��t��kj��6�EQ�j֩�����/&��a85B����uF�H�<�� ��.4�).��Ym06-��e^���0���j���1����o(��b�.�n:ݑ{u�#�� �^(�%-;�}������9t�[�r;*	��35i���J�"�1Iup�y~б�T��4T����ڤ0�afM�IH�2��s������g�H=L�k� ��2,F���Ӗ�|m}jߚC�Ð��
P�DR,�oW�Ϳ�_�Qx�� ��z=l�?y�o��ϴ~�"�iakw1����j�3^y��A���y��	^oV�}Do��+����RX���{J'�Na��cv�
�� �s!����tb�A��[Wy��jNg��ZZ�f����c�,��8U���S�;�	y!tU��HQ�Ŷ|j���Nz�Y�>t�ܛ�Z��eub�e��l�nb���Yػ�q$�3D����(��B���Jl_��� ��P�Z�*�E"^���l��	�oעG?'/��
�1�m>�xŅm�����w��ᩞ��d�������Se\D�)�3)x�%N�
n@K�b&\��g��Yҩ��(�|���C�3�l>4dg� ���P�����J%����5��8���6��n������(2��IU�k0�zMa�p򮣦��&�+�}�8���/|M�N�ko��cH�
�T,����{vvħ�@iuJq$�s���lG4�^�[�2�<�D��k�]Ͼ!�n&�g��"��^�oP�^/V�Ԫ�ǬH����J�_����sZ�N�w��ٓۮ�$���ڭ&^2�[l.o2wMr�jƺ�
쪺F��F�|B�˙/�`WP����ۣ���
�@�zb�ؠ6���v�y��V�<�5�wr��%��ğI��0z�H����O D��i3:$k�
W�3{��u"���-�J�����#-�cPΪ�:媠��x�#�N<"6x/��/@�JA:�£]qC��j�H�2�I��i�М�S��_z���8�a��=���9;=:",���9���bd�\M��=����hw�X��w����p�3��d�p��o�ŭw���ϓ���-�� aV��x>�^�Q�j��͎��}Dr�x}�'s��7P�FZ�V�dc��đ���+�Σ �#���iU�1�Bc;���P<Z�9��z"ҡD1$M�z^���J�ֳZ�����F\X�ܕ;��۳�o���Er�`'Ǎ+c�=�k��{#3���f=�����8o��Sf��X��t�qS]mq�ӏ"�@0)>BO%$+��m�x�������q��A[��~���UWm��E���"�l+�p+[6X!�d<Z��[����gͫ3���
��~/�a����d�z�z+T�i6jKg�p�%�n���(Q�k=��ܼ�h>�,�v�q��Y���
���ow[�Dŝ} X
�sx���?�; ȳ��X�0-��
��ۻy4%ѯ[�*�ۦj>�0�Ѐ��"�s���yWʮ�b{ͣ��*�}N��������|�T��&(;c�D�<P�'�~�(�jALa\ò�eL�c��3b����h?*�v @	eZ�E��$T����2d�YF�Z,�x����G�F��}հv{m�/ioziЩ�����,�%��; �Z�N�#yWdk�;+ݖfea�|7 �ۘ����M�Fl�Q�[��@��;��uJY{��TnYp-?���c���c�௔U���{}x��#���j�R%�B�j����'��xsl~�.NP�g��Z�H�Wg+��q)���S�}lsHҦ�����UآbJ��E	3�l��@6��9��#����n�fT��BP���H(�$�<B����/��Kub�?ah���؊�2ac-$�����|]ؤҮ����vfu@z`0YZ?�B=�LY���v��c�Y�=�	ΞK���3���W�yh|`�m5hi��CIco�ey�W����	a���	���ڹ=�d���Gg�;��^9^�xd��
�clZ��*��$����!v���_K�d���N�q��g��j�<z�zM[�-=������X��VߥrV�P[_�,P�>��xK\�ڟ�D�Ƥ���ґ7��T߈��K���4���܎{N�~��_/�ݕ\V�n��(P�~����\�!�O[�9�I��b5��S�:� j���㪟;�,�+��b� C!1�����q�45���y�b�lw��+����MI���d�\�]�ė7�˺;�C��{4�>?^`�b�uN~v�|��P��>�0jk㐎ϙϞ4�	�3�~Y�����$r�΂�t�1s��"6-�`�/�����-O���I���J�]?B2�E2i ����ŤR�����L�4(p�:����R��'��k���B[�����3�0s=%oX76(�6]��wI"�������Kc�eVk7�\�	+\<���V��KАG��H<,��*0��ҥ(讣�`�1L�;��/t��7t����Ш�S=`c�����5z�~M�5�p�i��[uK�ls�zY���>�"Q��8*y�ތ�QlCx�$��}b�G�����_ñ|���۶�z}��r�GoE`55�'R�qg`f�D�bj�۲���!"�=5�)���_k6�^!g1{��o�>�)�]�������o����*�_H1{�g<��L��#�3��@K��ǝ�����9Ϙ�ܦ��%�:��A֟�k��9��&mHzR�����7��|�]� ��K��͈E��颏и��]���O�5I�fA��y�;���u����[��u���Z4�#[��B2y����V`p`;��R�ʍ�n������v�*�Qx�9�������]XzzUI 1���Mյ��d��c`g���_F���V� �[\A�@kJ!��f��,�<A�.e��B�8���ނ�%�5�auB���ʳ���",;ٶ�X��7HU��W�H�L�Ie\����&Vk!`���lyKmG�N�אa�Q�VMq���hq嫏�q0<�m����PȻ�`'��Y�� F� �Q� ��p?'��< Dhm\�5���x>��gV�5	>J1��;sL�l�`sŸ1\cMB���^�%9K�b��^\Η�׺����`nU�߷68	���q!17ɔhK}�4�c�rFU���]�Z3���ok8h��`��^u�!����z���XC��{���GSVx� �F���!�<��"A����ي��
;/E�@l9�+}i��߸l����股����L� �`:�ɾ�QA�3b�M�vzߕ�s"Y�A$l@�*��>�:��V�^���x�2���_��(
x�Y}^�u;�_A"+�ْ���7>����f���m&*�q����P��3g&��G��	�=4I�B�yLc��Q���@
�ŀX��))�肮=@�S�q���<U��U#
_]���Y��3��+42�a�I��8�rC����8�I�LZ��^��e��7��_~:�Ӭ�c��%}: ����6�����@��=�h�hM��7����vB�G\ŝC���px�I�ȱ��Ka�@�����^A4D'�Im�-���˅�$?�D��j�pЫ��2&�W*�2ǕyVo0v��;T�O�~����E����:�!� ��;�IJ�;�Q��=K��T(�g7�/H��`)�H؆=f�< ��;!�܊�(���r7���w�D�T��V��4�4��p oQwo�n*�)ŏ�����2|��+���d��/g1L�ԕ%F�|�+�s8*PH��s�<F�̍��!MTn�$ʅ���cx ��Q�	9#uT� [_jj�$_Ն��~8GM�y�
��8�,�����'g*71V&}�/���֚��(<>�\���u:�z0�g� �h����D�'�/+^Ҟ��lH5^�#θ�Eռ[Δx�oe����
�]�T��}�ݿZ鷕��zs�[8c����Cx�5�ʒ��n1���
��$���prE��S� ��[(q���#�S�G���&��x\���q��l%�S�<�6
xD%-���"N�C�+"�/���Ђ:y ��8�k*h�ɮ��fP��c���f3�e��5b?�4C��I{%F�<��؜)��r�?j7�T�*��^Fo�Y�EH��ިT�Cy�Y酢x��l8��eeJjĤ4���M�Q+�-\5�2�����f�����__]��+׶���sԒn";׶ ^�5R�mZ9���y���!:�>��i�(�׵���CL{DM��+�+����M\�A��:cT�T��S+B��[{��0�p�9q�L�vA�l�D�'� g+�\n��{4�#ó?m��!Ǒ���&��d�L@h7��X�Q`�>�t{��p�.�Gf4J� �dv�J}�F.�S8m=��1Av���b����s5+K�!tk�6�b��̤�,֫�x�
���7�y~k���o�i�Z��#a �| jm��[�{J�$��(α�<C~�5�`�.�cM���^��kSnlΣ��k ��VP�>��2�m6�4���Р��	ʡ�!*"�@=E�H�P���č"wlH�R}#
H�K�;����;�<]�����i>f616��%��8���l� �ѡ� �Nk�V'�C0�JVݜP(��m��YT������0���G`L��
��M1guk���e��/�(z��?�%ܲ���[m�^��Z�k�����ِD���ߎ�P-e
m7͆��A0�80����҃]��+^�U3q
E���ʩ MŽp��>��Ӟz���{�"N��~U�ܷ����b��6��.nC�e�d�
�[��u��k]=ș%��o�6Q���.};��7��P��O�ZF_z�S���J5������2��"�e���g�A42kH ��wֵj��'�|nq���*W��ɲ���q黾���W���L�7�mJ�V�)_7����"?���M߸�~��S+Zj�w*���ؤv�݌�o�o����א?��/��2^��a���#c��^���*�SG��C����id�/y�$0��=�["^���հ��?ת�4�*���]8�|V������]C"yZv�*���fde{���@;�n�v�Ԋ|Y�b��"�҂o��I��ޣw�<�& �Ƃ�&s�4���ًBzW��TD聦-♼ˉ}����{4�=	/8W0��ᤁ!$v���:x���xQ1��p�0�D*�\�����v�Il\8asn?$2�8����P�K�k��L (n^/I=L�*�/��#�4F'ը
V�����ʬ�j>.�aj�M�x��C�����"�)k�FO}C ̈T �6���s�׷�V2@����x��ɤ+Ԫ߽;�1��A��0"������Fc����3�0�<�����	�ZD����h��~������۞cS�c�7�֒n6�(�#�L������O�sB_�c��+<����p$����z��\�-YQS��w�KO�En�=)O��a�Д�F��V���(���P�l�VK��lO�n�I&���\�^���]�QdBl.dLa*	)N֪������79([1�x��M	�;� T�N�*D���d$)sq�k� 6���:a��sĽ�D��ֆ,ά=��Պ_o¸�~�h]��2b���W=2	��g�qx?�."�wc�����F��ײ��+�F��'�%ZD5o2�0�� %��Pw�g��tzj�?�瑀�c>s��JD꣊8��s�7VJ�<�c!z��8võN�:�T��<��#�"M{D=�@LpD	Qp$�iJj� x��5 )�wD�E�J��ż»��l�� �*������+���%g�~�`B?�N�]��Z-e�q��e�����׹t�9L�P�k�X����pj��;3=}�����G_����`���Ų��C��X����ۯ��&�6n������a>�v����̾��W��N�6Z��?,�4]�Qg�UQGd�-k�����&��qP���-1����M�S�/d����3۩#�ie8,��p�f���
6#a�4M�e����n'����;���9��^��GyO�/�=�(���h��^WhM�N�S N��[/%���yI�Q�L�l�l3��8MҌ*.�9f3���i\8'm��Jb?�p��6$��W6��,��֋����x��<p'��9 ��s�z�nvr\E��͓��K����o{�)���U����.c>=I��%��"p�&7��E��TZ���U]���OK!N�[}LK���;ny�Ӡi+�f$������0x-�=��7@��i_=X7��^�э@�I�4�>�ǭ�
�G�Cl��c�� *&���*S	��؋>�������T6.|�dЉ�>]�9JfMO���2�t���]|s�F�Cb�P�11�8��c�=k������-Q�W��ڱ�v�0�\.��3�j�+��)��\.�n�v˃,�B�>�T���3Sm�l,����ܮ�'���,1��r��upj�0	)4��cܝ{��8��~h������ڹ�� ����Rn�@W��О�L�v�U����mKk�T�=���\�U=�-���"AUJ[�Ä� ��ҟWO�̏,��s��!�l#�R��b�9y1:$	���x���v}Tk{����_S��u$�J�K(�n�ǉ)���Ӂ^�@�Jn����><�a:W&?���~F>0[]ȭ��suYIP߭��f1df�klN���@�1�y�ӄi�*��$L0g=�,�p��)�!D��ʐs�VnZh�k�V�������������F��bq���֞�>�.�Q�����O/�БP��g����Q=���_���o�6 ��;������+�Ur �wfh6��������5��"�%3a?�k�~��Z�ƀ�ȷ��i�!j�v�t��+��$ ����j�|�� ��o;���O�8�Ql*�~������q\��/sy�-��0�%��ekUm/va�9�ƾ���5Q��&�UǊ���4�5�{$��M�BH�'��!����� +�#_��Ĭ��TYP�
4^�Gq�l	$��"�op?&���:x�$#~�ɧ���ձHMu�SX�)��>�pUB�WYG�z��E�L�Ldvۯ;��?�D$���]�u���v;0��L{i��z�}d�G��Y�G�TE�q O�D3�KB���t1
�Z�E�U$����4���|�i(��K�2��Y��J�O7Q�F��HV�)?a��T��t�oc��	)�����B8�3f��ִDO��9�9A�*J�U u�.p �$����O}��``��@]�5��,&�����'H��c�*ܩ�ZJ��z��]&�4ȍ�zs_U�����R`���뜌hi�z����9��%��q�ZE
�!�hGκ�qֳ>�p�^���B���a�#�n��$!�QLv6*��~f���?��v�rd5�^=�R����i?��̤�8�5���f�����L�'�Ҷg�-�>� %]�hM�t�4���-vN%�!�%��h��D^��c�(�H�<f*9(A�hg�4�$%2��G�E��h6�xO�v>�Ƶi���F�vڀ�k)��A	���w�F4�àh%�@%<\�ɴY�����y�O+G}֯w�oؕ�8H�\+n��%yI>��屽1"�ڳ,��
�>[>��&@���D�g�7U1��s�'_�-�'5(zr�h:��%���,V-��}7�³ Y�2��Cdk����b�2ZVlC<=g_&pJ�yq��&c�H�3ސ�ք���\d�m23��3,�/�k��Wu����s*m�*���/J��$e09
,�l���@��j(���x����.V�O��20�d��Y��P�.�/O���P�WI�t*�<w���1����kjD; �Cm
өmk\d���n.M3���MOX��
��7�d�'��d�#�7-�	��n��@�땙��ne���a�Ju�B��K�(��?�B8�l(ZlQ���2������K�:َ�	��Ƽ �!ɤ�ʳ߃.k$e��{\�cT\C�=�����&�Q^<A���d�]��uaOl���^^�"K�P�׾:�/(��d$�@Г̡�&�n\�rW6����`���/�������~��������
��Eo���xsO�|�!��;���"�ȡw�0k5�V��Ir���\��0kj�rϴ��J;bܓ�N���z
}��nܒ��~���#�S-n[��w�p��<�!����n&":��j��3Ώ��;�hT�/{P�	yɣX�hˤ��A��|o�Z�-�(k#�T���ژcAß����1�].��^����1j�U�
���=$����=B��kIod��e�&?��t��+�X2��V����S,�[��p(�}�Ϥ}�F���W�YC_O�8|R�Z&+i��ߩ�d�5��:���O=�92�Ϧ��/V'���g56�T��M������i�j<n�Y�
.�q��@��xg>�4Ǟ����Q���g�ӣV���F�	��M��+�U��I����}��n/ﾗZѕu���-��O� ��s����9������0�/2[1�|���xC�r "���$����RG��tT���)����p���4��݃S�L����A�ޖ?���'^lA)�\���#Av:�rsZ�Jv=�Ռ_PN�Y�H��o�z[X�7"̏W$�����@N�?���b���|N���c[�����[(8w��ڇJ
N�\?�^�}
c�h���Z�����˪�ϱ�ڛOyu}
����Ǹ\�^4Gue�gP�2�R(3��M��{2�3������ֆg#��?,�TJ� ���>o=��%�!N�1���#�4D�֫�:�D������+L�r�-!��ʤ�Qfve}�� <!�v��s��f� h���:�A��W-����I�\"]�8�y<�!]�	�H/������_��ˡ�)C~���n�uֹu�V�Z��56���=�_���o�#|��2N�7���&q����k �� 8�U۷��:�����WDge}��cIO���,��slbp�0 �Cf	o�������w΍��s��FWx(����,��@~Y-å���?��	M�	���L��ް�|���"HM����9��[]���,�9��oe ��KJ�u�ݞ�����M��A��b��H�ۧkv6���/�o��H��N��kr��I@�X٦�u�{Sz�k\?r9���2�/�ܱ#-�1+�숏֕|�^��F$l��AK���g�%7����F�0�� f��I �� �cZ��N�Ԧ3.g��C�}�6:S�2;�835ˑ���/\\�:���߈&}�G�� t���eK$⸩�H�b�ckr[@�fG_|�2�6~��j&�9���M��˔��1�0�W̖͛+D�:���H��S������w���@�Ud00�A����b鶻�B�	�6:�6p^�s��@�wrT
ʈH]�Ʀ���,�v:�����
ℇ�|-�K�z�y�p�d�+L��F�����8>�n�������"�?Y���m��Ĕ3�c훜]�$�ɶ�P����
�1�F�]}4�sz�m��9 %2_n!�����.BI)��&҅��^9#7��}���I��J�n�i�����=hf�}�ÿƤn�>�b�+���{���ٚ��4�f*s��/�f9_���2J7��8�/�ZJ�*c�1��۫^\T��H�֎j�8q;=o	|�>���t
�|2+�/�F/q�W�Rʓ2�fq��fՆ@�/�*W=g�ގ��t�3�b�-��z�U��y��Z\h�<��Ac������	rwSy#�f���O!f%��j��q��9	�X�rƌ6�;鋠��T�\b-!���-z�y���	���EU+�cxu.��Z��zyGAإ��pv�t�P�wr\Z����ʸg�Ͻ��5���/��%g��+�x݀l�KQ=${W�|��Y9�0����+��RO�q_���cv}\��^���"*><Pu9�X�}1��v�󹣅���7y'���*"��D�N�y
��V��tG�=�}�;����:*ܠ�gNn�,�[1z���Rx��j8�.#���=�F-��	IY�3҇|F?�,Ǻ�(�#Ac���
�r+l�GC����!�!�ΫA�DM
1b���5�8N�L�k���դe?��B�_�T�܃����H��f��J++6N�+�%? `�T4G)lS˶�~<W�/�Czpw k�"��K�2x��C�˸,($޸S�.4E.��k���1GG�s?Ә��H~}��(¤����p=�[!��FA�L��)�:���"�g���e�Ҥ⫴�IH���"��$-H����u&o��%m���9A<b�;�`VF��=�Z����2�e��]�p�6�QQ`����ᦿ�R���iE�qXAyX�?h*2�%*YH۫��&oѓ��l J�8@U�	�� t��a7���Æ���)C��u�Z�f��Qh^ļ_ٖg�0��Xw֐=������'��㛈�-)�e����C�	�K>�ƛJ�逥��0�3����5�<��o�#�?l�I#���P/�L��֌2��7�U�$Pc��(W���.�B�d s�p�6S.��o�bޢ+��M`��i.� �M�;�c�8}�|�����22��m��8U�W�EM��r�x���ҝn9ךi�>Gb��F{����p����e3��c�``RlV�Z�Y��l���e��5/]\{%G�Բ�]΄���U����2n�ԫ����E?1�@�Ϙ�z��F��䮋urf�_�*l�~B(j~�w!��R;�
�T!
K�hVj'k4���x�fM���p���ZЕi�A���`2%X.H2��9�i���p\v���'�����[����b��S�죦��.���u�5T��fƾ�`e�X#��o�9#���R[���X�~��5h�������6�|�^��T�b���T9��z:��"���a<g�5�'Mo��'�J���"#ُ~�k��dǵ�g��*�{y>�����.g��^�����;�	�9�Vݮ�5�8v��鯘�)�f��T=��6���m��*w+y��O�OKm/*��N&�p�o���N^��NA1嵪 ._�x1C�
�kH�)kKӒ.Ƅ��F:vΈ`.&���k��W���˾�n3��!����V���?c��.��Q#�5�H���^�1i���4Ao���A !��%a�!��
Y������E��:]�U&W���f��D���My�s4G@,�yV9,@g@�w�|��t��?lQep��T1������3X\Z��k�� �6Ǖ��[UB�n�Z\���>l:>Wه���R�d-�]��;>{��`�g~{n��*g^��c^`X�)$���(��R���Y�b0��_��tN�C`�S~T+�b
��nX��+�;�X���O�v�6�׻�ƴ<�lu��ߕ�0��Ey� �h�#*��H���N�QCX#(Qu�A��rYy簝S��������}��z8��iȿ���~^:����W�Y>f{�]�w�?���zf��O���~���B
w��x���7#��:#��9c+'��h�5�ZJV��1&F�A�}��v:��B����]�,,i��A�]h����fG��f�B#ꑫZ�4�[��|N.��tAOWt�>w� v�׸Aa�l���G���8�������It�PrK0�隳]�-Ɂ;A����*Jd�#7���q�����d!���׏Y�F/#�V�Q7���Z$N�I�|*k�	;�OpV�B��Д�D��/45qZ%��)�n�6�Q���F���A�C���W�+��K�<�CN������UZ'��W~O����#�["dUZ >+HmUK�<C�Y+�{��}���o�{�Uw�ވm����AL)��Ou[z�.u���L	�g�2xI�P����SՔ�9������{�sE�C	���T�'Dɠ��������>@�es3$�]���\���@�^�����!�N�����v[k/�)�L7_e��+a�J���%�}�j8�b?΋tX��v/��O�K=��c.A�J!�F��dI[��X�UN�șx�)�]v{�%$��$Yu~G��t:ﳸ���40�� z��P"H]w|�O��<؋�D�� &Uo���~:�	����_~(�r/�
��w��K�x*K��pZ�+�+p�D+�0t�ދ3�YG����sW��a=�<�2�4ޑ(Y�y�����Ox���j��������0�٥F�_:�����_F�g�tJ3�f��=�ʻ�y�}�sؐ���f�`�^)$� N�@OZ�\paĨ�_ h��d����6���A{��+o��`c��Ɵ�_�8S�9�uթ&�>�t��[R�6rR��cp	21OD%��nE5 �������Q��Y�/n7C���l�ԓ�<&Z�j�����N�84Ȭ �6TE�+��4u�g�Hi���z��)�	F�p���~6���8���Z�1��/��^yn��\r����<"�Ѡ.�����
E��cM��ոr�%w�_2
�����ʹ��/�"�����+m����*I��"#�#v���I��W1�W�$����Ёb��S�������u����N����D+��%e?>��t�A�`j���t�A�C0It�׏a$���x_��AX8�L7�}�(&]<�ͯ]|z+u�e���뾌S|,��H��'c�Y�_|^��1������F~gL��n�;�ï^�uc�}�����py��U��q�U�������#�S�t�PT�N�Cn����P��$��\����<d���(��A�\/Ol�1��I$���]����ú�D&�a�Gq�Ȉ`�R��_Z ��"�N jiI�Wzj��w�p�}ʽ���D>�hD��F��X2K��a���prj��N�Ǧ`����5
��VnO���a��.��IAF.�W*R]�;�<t/��%��?��-XL�*!�[���D��8��D�:Ê195-�I�"�p&���w��H���ٔ�i�ꤗ[i-<0��D�A`_I�:z�T�٩o�o3`0[��<8�'�E�7�tg�KWYn�������b�ǝ� �nml�����!��!���wA��|Jx0��܈�(
8c�އ[I���8���ݼ�gm���C;R��n�TV�^��7�#�v)�g��L&M15�},;���"�V*��G�`�8�c���՚n���]��^�}5��³����f���u��f_�^�)ꮒ�H`�h����3���,������i`��Gᇈ������(��)��m�Bb�Y�|��/�3���^ܴ{�"u���oVL�a������J�2��Ԝ����Q���`���c0�Y�坿�г7��T;��7��~�׭���N���kQ�[�u6?�G'���@�������OA��+Z�C��a��T<!eyS���)G6��S`�g��28L���T�8�%�>���{��cv�=��~�Kg��Do�?w�Ţ�R!�[kX��uMv����S-<w5)������	I�[�":-����E�i�N�1�}�60gV���I�98Q�-6�%��M��q��=8S�PPܵ�*[�T`����Tc��G[<dS�iy&d|�Q���k�I�s0��b�0��.�{�(U"KM��X�@�������4��QM���ִ�r�8�Y�1�=}ѕwO�|��F`�����p���Ɣ6���/k�uw���+���gvi�����6(��[?�s.5L�z���S����ʾs�~%[Iꠀ$Cf���<%�G_7��5 ��*$�90��2��W7:�Uf�vYy����I$8k��ľ<��9%��G�X����y1�g������]�c�����Ǣ
�a�K�UTǄf'V���r���R{)�zؤ�\����D_���bcM���h�	? h��U(a/.RZ�B�?M�)7]{K/�f*� ���>6�c����gX.7�*٪�kn��Jb�"����Nqen#�.���U�Qb��O��[�H9aS��[��$�V��o�z����	���sgDv�����n��ō�Ug��}dB��:��H�u��n�@���P��9��x��O,g��J-�`�"�.��p�x��#r��weL���Z� ��mÜ��z(�}
O�\������� �e]�4��4ĠΊ&�^�]a�Xi)g��]M�gpY���@��aم�:x��/�+�G�fG�ߎ!�bl��.�̈�뵶6�n����*�{*�#�Y����uQա1U2���c�J7��-����T�,�d��L��i�:	��Ka!{P�@?N&;s�����yٻ�^�&�\�I�s��jl�6���)=�)>]e9�C�Or����$�'O ���n����}
B�~����A�᩺���[��%��� �u@�ăa��ܭ��}�(b���M�,�����U�؅���q�#��
zZĈ믅Ej�|*���;h��"��r{5������ߗ
�ȫi�{�{W�m%���7=�ZY ���+�)U]�Fp�2F 7q�����2�r_���&]Q��4�v'��O���:�i�P��� 㠚.	��1'?���?_�{Ձ���Wq�/���Ug"��cʏ�d�	����JN��Kt8*���<�{��#t���L6���Svk����iխ�������w�/��Ĉj���ݖ��M� �pX]k)��<6�|}���Hz������늂A����%��f���C����&̥����M�f$�|�����0J�thnG�����HPW�E�F��f�N;ɭ }�x�y�h�P�'E�s�,A���ő�B���w������>�˙�hj6�'��Y��r2�߶���t��p��4:�;�#؀�����"pԘ���I����,gsE�g&��e�PI�ĬJ%&��Ӽ�\	�S^s��fvp���"���OnǕ�d����iI�0~�m%=��gZ��Vf��#�(WW�R�w�^<ó�+
�"��+�?�*����)Tb�C,���@4 }�-CB�W��p�~���@�V�-9�'ź�L���"`3*�T�m�VKo�Y]k%9̒)���DN�z���� i�I?��m�}���櫁-P2�'�ZgiR[�ġ��V�1��� ���X����.ߥ�ή�W,��<�)(Zs�"�c�9(����E��>خ
Ej�"r�q�eX���F.2�'����ZQA	�BsM��7b��.;<�B<{ ��D[��<0��z����A����O�m���J\Q�JXVZC9'F��B,F.��>�gc�y�l���ɄHw��]˹6�)�i4V�⬁�LrG��'L �
遹�}�j��M�cF^�g�=LyR�u�P��YZ ���#���#�A��x���OUԝ-
����?��5Q6!rSG�<͐�ވ�_�$�풏�/̣��j�tfֻ��I�S���@����^���Mzfe2���7��%����Ј�G]hܟ��aN�:����b�Z�FD�c���xw�mF?"5�9��Ɋ*sJ���_��:a�4��&	s �˯��}Cʘb5g����II)DzQ?��Yi^_�l��N�$�So����.&p�5�'a��ZO��?��0d`D+��kų��ad4Bn�WA���$)�]��yE��ш�ղ~�؈�R���9����)�i8���+�`�E�&V�	V���P�6j��3������B���k����_��P���zxW�h:�hfr��p��_�0 �����3b��4���-�,E���\�X,Y�ԘO[��Q�Er�'/jkx�8;��
��3����F�8�W�D$�*�5�޷��Q2F�� Ug�^1���jF7n&8���l2s�3��4�����S�\�\�}�iRF�7�����$�b��z���{FmSZ/�/Y��.h�2eWI�Lz"1c{�#�s�2�D��ȄaOBJ@�L����dL,�~��T��N7��g�H~�@n���d1������Ac�h�[�6�H�0�!��d}ҝ`4���F��Yq�تj�P�v��.e�#��0j�������`�=�d�HCb-�8D	AV]��|Q�.�0hT�#��zt]ڵLo&\nW����ҵP�/�4���'B/g&���;طO�s���y1�.�0l�Z�ҞT�j�j�t�cx��Y�y�c�¤j�C�V��)~j�V敕��L����.������ފ#�LLL)��95+�]'�{�{���nd�,��K���>�:�g�,m�j]�qRh�}�I�MK���8�p^7��N��7]�r��
6&_y+��>zjX�W����'��AFdY%�1�o�e�)����4@�6�\]�&"�TZ�U���U9w�B��>ݷ
��_Vºb���(��ksZ�a��%��xa�\��d���l{��ta<J �M�?��e�Ե��gn�����7����%��Wp���o��2�M��R����z���{��5]I�S��T��ѾC`L��֎���DyD,�(p��� ��Ϯ�sЎRQ1.�p�i��/q�!��d�d�;��i׋}��1���W�
;�J��4*O���%ep��VJ1u
.���,�~c�a��̇���D�
�:4LA�/e��j�������4}�֩(��:��kKQY[�D�e�Ҩg����@���	���f\�ӑ�#-�ݠڮ���>�3/��k.�>:J��NE|�d㋇|�'�)��{�(�f�G�a�6;�>����>	����A�a�*��RBii\��*s�FC���;R�� ���?}�Q��'�Q�wn\����z�ʃ����'�Y3� �z��� �Q�UQT�b]-�1� �0�A$1�VOM na�
��O�L�`y��ޗ�]���4,���&ᆜ�"���\�	�U������wj������̗b�a!l�:]�=�/���$^���K4��*k�{
D�u�(�K\�)\5li� ����D�Y��w�WNM���&��.����y�F�>���=�͙��b���V��!;�xA�~����-�7����E�c�fL c*�:��]UL�I[}
�'�ǃ+GE��Z��3�����1/�=�y��S�:6Gt�'�]U���I��|vjԒ�W��F=N�3�)r{l�������{�T��q-�ؽu^d�rU��I#VϡA�-Vy}�]	�F���� j_� �>Q�ѓ߉����,�9Pl���v��ӌ�$;�`�,�(L?S�j���sJ�,���dR�7<uÒ=�ae���Q��P�Xr��g�
oMA��[��e��S!��m��q]��`(u�(J��K*@G�H��U��Wd�o�p��a?��$f���o�����lM��=���:;�:��1�oQ
i�Dq@�)x�&]��Nd>�E��v��7Q'mb�)W:J|M�x%h$yT>��	G?J@5K+'N�ܖ��%j��'��[%�U.�[VX�p�cNbo��1����-�0�x
�ͷ�W+�����k�ƿ�a���L4�w�V��P7�$��o�x��m#k��r���I_W��9~:[4u�]ciJ�1%���톥LϿ_�^Vs��M]�=���Q��Oր��.l��P���g�n���X(�]a�8,�5f?G��m����~�/σ�L����3ȷs�Ƣ��m�˻�`$����~�UQ(F�OQZ��,gV���ՕI{���y���^��O���pz�Z�� �/Dm�W��||`jȑ����ѐ�HY�k'��o^�&6�❑l�G����؀������]�����@��,�,�*��x�3x���A���+���ˆ��1�V#�$[��6 ���Z��I�K��g����ʹ�BΖ��2JY�x'v2�����sr���9�A����d�D���-����}�J�ܝ��Š^��<��v�O�/{�G{si�2W���.1
�F���"_�eϬ���w���? !�d(��]F��9�o#�m(��[����ƨ֦��/x���f袮)Q���3�I��"7�
�TX{I'�C���g�y�H�{��ʩe�}�ZO�s +���y0��QV
oK�~{�摈�2�K��9��m�B�`qMVę"�B��BJ�U>`���ܶ�F�}�	����,vN�l����r�Sf�L���j�V0=� �F�u�����1�m�
��稙L�F��<2�ڜW��2p�{����߈���b}I�X.���]KyC~�v��	Y�F�=sD�1'�V�5'��耎kQ���3N{�_Jq�B6LE7�B�|����d%Wd⃸���o��R�ʮ��pM�0�+"�Wprwde�f���O)���bm��?�Ύw�e*{Ѥ��𧍶,(�����6&8�Kˈ�Y�sb�t�d�l��$q��UKL�ūǽDv��W�㱯9G�`�(L*p�=!4���{�,�ժQ��Q�}����� ���3+p.��A&��L2���	��}���C��Ha���A@w����]L��EI�`�ޗ�C��<��w5�E���r��6z���Rp��FF�L�����i����cP(��R�1<��&Fp��]<���K����|�	�X7y��$����z��bh��t�x�}��	=���&���N1��d�U/u�����~%R��N�=�E���D[���ۿ+i���RZ�7����x���V�q���y+�M{� �t�D8�5�B	�x�ց�KϠ�C?��|�2�XA��;�8���s�wB�D;T1fk5<�����"?>BC
�Z\�����~�N���t�QQ��]W���r^Hp�[G��u�qH�&�z���)�7��*����m/��=��%9�([�/��0��L���i�-2�)7~	��D��̈�
��3H0�l'�}�m���UQ}�Nh]�q�1D\o1 �Lx�g�*s�.x�(�Jvf��X -u���C�R@.���l��ifW!5Y������3�� ]���"Q٘�8Jl+���v''�j��������9�ʧ
��ʍb�C`A0�ԊŒ���}�.X��\_E�IR�(�l.��F�Bj
Nz���$ⓥ���<8���r�j-���A�"��.�۳������>�X��J�ʦ��N��8]Y��<!v\㣏��}��#����"p��ͻL`lً���'�?KW�P|��?����*��[���ZA�GQwC�~S챋�o 0���2#��)���^�?xl�ׇ�v�!����\�߮��"�T�y�ב�(�5N��!�汄N�j��G\~��� Zyl
���İ����=�f�w4�.0�p���S&����n`��D�9��@�Yv�J�mދ<�&��{ӊgXT�G����[릭��Ȑ,�t����c���5��^H�h�N$S�*����$ a�h�͏��w;Lcɨ�����%B+�yMU�`���������w�j�|oZ��������͚~���"T�yh��W�~����y뛄-'@{]��@���x�{K�)i2٤�����BlE�h��^LY���E�K����i������h�[�>.Y����M!��Ͳ��+�UyT���O������W�|�}k:��ُO���";A���ƈ �l�-.�]�vZ�v���8����RĊ5�aG9�Q��Mz.E6fE��b($OD�4�u���<�(Gu�2�>"v�I�C"�Ǟ �{�*S�M���C-;�����[v�ҢU3��$��|�(?+e_�%h;�1;��&�Q�x<�;*x(%8�%^���S#pO[�� 餱�S�;^F��z���f@���z��eB���x��Q�0��_&���`i;̟�&��۽'. �d(�G�w�!HM�dd����>(�	��'D���#������X�K�.@��`ę�r*1��VF����: ����4�ȋP��s��v�p�(T+�ݡp�,�g�4�{��[L'��]#�c��Y�F���4�ʑ#�U�G)8X���a+�wX��㭜~%d��Z��0�������ys��f����z��l=R�h�%ٽY��ϰ��q�f�ʴj��Xa��h�:Y���壢SQ
��Hl��Ɯ�Y�I�3�r��4_iNu��G%�4��񛁚�-|�S~0d\Lu� �	�6���N�D����!?������E-E�|��F��/b;���^����A+���	D����������l5\t˸��f<�������Y�N�T��o���<ԳS @}(x��J��hJ��.��"����FRb�21T[��c�Cȟ�b���m���1B�2a�7�ۺm���+�c��e4�ϫr�G�귘#�u�a[G �

y���1(������-�d��4�>-������:�@�c����R���.w����������
�13�	�73K�a�z��q8%��4���Ԥ�pl���iq�=q�&=�iާ3�u���S�e�l;� ���f�@e��B|hN��$���C��~"�7���D��j�^�XvU��$+��[ V�F0���t3L�N�x������U ������G�����Y���c��dH&�P�HpC�ªD��CU}.A'�W���MT��U����fbDG0h9^=Z�|]�1o��nnڗ	�X���;,,�w�s&K�e���f��9
%����n���w������h4�|C�����Ѿ��@�>٧B`��J�-8C� �ނ���<kgD,�����0V쾸)�j����oD��,�C�N8�+�����������M�%��[u~qP���`�ڍQ��y4��cַ.2�A_<w�v��m�~���JD�b���Z��+64�5ݴse�ٸ!�Ԋ���.��ù�������:��DU/�y����4����s�Դ�Y�ħ���g�(ڣf�l�^��"���)%t��P���]ȯ;^_)���B\=��!
*�U���A�az-_e�-'���P�k?~І-f���_�1�˦��A���0��;�� �=$f(� �q>���>�;�A���|J'��9��k����`��@��/�K�������{lI���4�Su��83ć���Xm���7���������UCU�>�ٮl}l������O�-�,��~V�ml�WX<F(!�o�޽d��*�=���6K�C�&�Y��N� mk9{ܯw�۱(V��������o&���a[v	n-���;����H�g	?>�����ч#��Y����gk�D%���O��\Z^�@�=���q��k/�bN��#}�H�~��a���Rt��*���H*M����3?��}-�8��s��Q!W��v�����v��m걄�1R��Ȫ�Q�q�G%x(�롭e�4��Nf���8E��X�=�c�ሦ�\����7oϰ�'���7�gڂ�@�e�CHH�P��]W��Bi��?�YQTH�'�i�uNu�A�ɻ���z��2i:�p� ����!j�L�M����8C1-�3��aU����I�MG��[�^�k��_�Z	~��W��JP�z��k��)�pB��%����e��6����ᇮ���¹g܅��H�֬��z5��B�v1�c�[�>{��3e��Էb���X���J},����W/5�KJ�KՌ5��0r<��
cR)�/b.� ����$�^c*U�:z�	?%j�+F�W�p��v�r��Y�>T>�p�����f+����ݺ��UkT7��t���-3�z���WU�ڮ1ը=��h7��ie���|���1?���25"�4'w�;��NFQͲQ�I������4@Gʕå�b�ы������KD���>��}��Jt���ϳk��Q�1�p{�����	#�D4��3+�WD���铛�8�V)tB�濂	��t�4r��)�e+�oO}~�R1�U@
�<`v���O68�<t)�-y;��ɶbS���*9�&a���ީ竎��?v����Ѳ{I�hS�>��48
M�A�1)j��"H�D%�\�h�;�ᔙRX��R&gh�1�E�}�c�#�mD���V���?nǷ\�#���� ��N�E�~�PCq\R����������r�h:WtkI!�~z{��bY	s�,�֟K�%�K�(bC����{$���~��
B�.@������E��(�c��N��T�����v�؛�3�,83���F��Xu���pֿ��㥠8�������ͳ :�C���ҧs=�DN1��iH�@�Q�RZ�ѥ�Y3��?��ܫ�����9#(��q
hm^Z���uv�U,�Hq>ǌ�dru��h�[:A!`h�Vd��{����6�X�$#D!f�S"�;ު��%��~q�kOKx��6�'@8���7��_��[JX���i�����4��A���"dn��"s6���F�u�͗w���C٢q���O������Opy�\|Es Q���\ªF�J@r�k��f��4}�MS��'J�Ld��v���E�b˄����W��
���<���~ڑ��+*����>uRT$����'���9Y@�Z�PoNEe���^�4�~������{���{!�z�.l���S�nTHj� �C�=�U�3s���`��@��!n���!26�+����]�v��qږ��4L{�S����j���Ȯo�+�!z��Jv/K�-�FK�<�W�Bs���8n�Wϼ��
���X�'��i;�yvFw�Ø�^�	!��+h����Z��׎�<	��%_��V��;xޮ�,=����흿��^�h:�)�x�`��?Sd���V`�����Ϻ�]�!vM�r
N����F3<��ĵ��#�$�Di�ۊI�$����X����D�Ұ~�L0�=IWA��=e�;r�4t=�YMyD�/T�qVEى���B�j���F�Se���ё�B��`�Ĩ�/M�_]�b���ۑ�1�����|�ZԠ�
�y��F܅p�G�VV��( ��bC$Q_�Qk�s��p���y$s��Ğ�OE�, vs���0S��NE��t��O.��.�;�z���(�~�݃���تdy�E^�:4��GP�YRe�|T�4т�� ^�A�(�1�@O�.�ԞP��B��^��˖��I�H�|7�䠺��-9�Qee	���v�O�B��ϖ�Jq��kC��	4�n�}����~-�K��Ij�SW�:��������ڔ0k)��x��,�rkBo�i�ͯ�����d���f��Re1�
�8[�C��.�rE�7�ٵR<t��-��{!D6���B�]X�ao��y	�脒��a#0c�-�e�����q&�Ω�3�[�~t#"S+���HH���X�����DV!Y_���^��J�G))�>�/D��S�~�&2�$�G`�� �� ��e��x4���{������^m"��38,!ab��jG��ή�RMo&�
������R"�f���qG���P�魌���[�<�/xy����`r8�B��p��X�ҝ�"��LL[P*�@C~E�+�Ϯ�S��M���)�2�V'�МZ �1�!X~#}M��!=Sü�/��믊'�ut�x��>���.�	�}��t�j�4)�lݽ�� ֻ��R9wo��z!���i�/��k�/����`܃�����ڿvxT�L��߈3�3M�!�n����;��|j{�Lg����К#����H�0�>Qs��߭��ω��REI��[�l��n���f�<�b��a��|\�����CE�ps���t���=:}0o���pI*�� ��9g����������b٪.EJ�+ឫ�%�`'��K-��ۦC�6h�@HGkR��wѶ2��a��ZQ��PƋ�;��}0@P/����R	 -��Gnӯ1^>��9�]�<�Ą��ѶA��I�
0A3oT'��A}�9�tA��G��l����.w��G>�ul��ј"�6�"����OUb/���@�_#[P���1�A!���&S=ػ�mV[y�k�8+ז�U�,#h�����i1J�����#�� x%�U��
�o�\(�>7]-�M��X��DS��jV�D�B�}*wM˶��widfc��X'�gg�����n1`��Ϣߧ���hM�,��C�2���׆�k��΢�3j�-MU���ó`�����N�c�Se	Jl������!9��M۽���p�t�D��NzC5n�]zMi��<�����q�L���\d墱-�RԺ�<������3�~�i'2��vFy[�P�gs<��f��;��ø�w�K�M�AIļÊ�������ut�W�̫�;�����t�%�rQ��KB���Ń�&eғ ��UѬ-h��E�+B[*����+@j[e ����>����)�%�en��Y^G�Mvg�u�d�Y�" ��p����J��}5[�6�I��5�ւw�)�Q���hK�ї�
�6zWX��C�`���6����S8�.�t��\�H�����/�!�ʅ�2� .�������F���.�EE�;�GCP^Gi�A\��8�e���FR��kV��&mt��t"�?W�Ra^J�ۊ�g�x��(q�	�Q����+���'JVY����^�^1
W+B�����ڸ����C9�w�Pg�tM�H\G���SjY���Jn��.h�H/����њ�P�m�ޟ�,���}EJ uK�F��+��b)�+d�lׯ�mú�N��XG�LǷ�8�����&�9�
��HMH�Z��*�����@�"Ֆ�ɞ��C_�	1��y����3On\!��R�Dq�������τ$������B���ZsW��;���֝8�����|,y��F�Sv����؞��yR�\�����X�~M�z�&�-N�opW�!q���@���2�˕+�s�����fi{�k�����>����;g�Ƽ��qC��8~5ԓ�(��2���l}o�;�t](te��":��%�iR�H�8�W��XO�@�v5P�AL`�t��Ɖ	F*t�c5���`"�y6��
�+	����p]e�����w��9��e�wx�5�>�5��F�qm�~����O��?}�\ZTR���u��j~��!��u���%����غJ�B���v �H�p�YNFN��:y �c��|~ʘ㪓�&b�Z
�x��������ThӴ%�*���?\��{�n��ĸ��N���P�G�p�M�4Oز\�t���@6��z�$���q<h�C�7Q�j��5�
�m�D�$����k>�)w68��6��=ɸc�U$
�0[�%���p��3��9���-IO��������~�¤�k�h�%�ɱ���Z�9��pu��W�덾��fS�}s�JXޢf8]�[<YNV�؈��F�׮As�w�b�}5g���Z�u�]���s-�@��[�;�J������f�R��<]#L�f�7��`���A:��_����r�䦰q�ԯ7������ M����U�J��CĪ�R2����`�m�s�ڴ
����2$l`��:���T��Z��S�X�����x�F�4J�T'&��#8Y�w�E0_��U���P$	�����5�L�������D���R}Ey �0��J�҄$Kq��+KÝc!lw`6p�?y����'��v�ʬ}(�'�x���\�|���P{�Ӏ���C�eU���	�`'���'� �*�n`�s��M<I"��Y��kN����Q$)Pz�Z��`}�q�k(��.$>��� �vi���.6� z�a�����B�\��zX��A����4z��9xN��~��
_@��N�}N`��2���|������ms?d�� ��/8��r{=4}���xr�D�ò��*x�~�wAHl�F:Iel�I�Q���{��kl�0���b ��G"f �8t�i�!C�D��9����l�aVws��IT'̞fV@;�vo� 3�F����AnҡHұON"��j�."ƥ��+Z}�:�p�z+ȴ���3���ᓮSEv3�Ku�l��t�}P��^d1ikc(��֥�K�EÚ�x����*a��@��c�$B[<�(='2�ui;�i@��$��S�@�$�-��]- �܆����ޡ��X�;����j�� H�|��ؾ�g�aͬ��9�S���[VC�H��i	���J`��p~:[���3�_���$�&:Y�llg7��a9gm}*��E����Ж��Ȥ>��G���/��c��}:l�B���ojbTc4���(H�/�l?95z�SG���5p�M����nO����^ͲG��1����L�Nz˲)'e�]O�,�iJ�nI���b-�bc���b2���ܕlv:5T%t�-j;n?�R�_$���5�|���B���
�����g�N���}@�ģIT�Ⳃs��@�8�X,3ID��-�X�G��$�9[#hdq���Q4�m�v�G��j{��֏����P�Uu�־��N��9�n��)�瓎L��c)�)��T���zpܚqi�Rc-��e���O�Q�߶niw�ߓ�u7�"yPk/���Xd'����!�ʴ�XB��1\��d&a�;���8��e
>���I�hJi-���-v4S3,`a��
@ �x���c��8�8����㫧
b�UAU�U�j�p�
Υ�d7�����9=�أ�$1�!����s��鍻���jب[�jS_�L�r�Z�� ���]����Vm�8��>��R�^@�$N&��hk�a$����Te�h�C-��W.�,��c���#TO�bߩY��T_�L3�g�:�����7`�6A�C��i��Ҭ�k�+��J�lT���rV<و@�� b4��Sy���j�G�*i	Ʉ�ò�g�VTݪ����.
["L����tp*��*m$��q1F�G��6�^d dJՋ�n��d\�?��	�,bb?��B'�ڮ�8M��x_�q���ٽPKZǴr_��� ���V9��@����YF���S-_!Z-I/,J�u}�Ѿ
�����:��>�V~E�؜�ן�b��+=9�=�~12;�Q��^X��WT2 �J<��B6lh�V*Zd�'��v�`�r�M��SS��눇*�o��ޅ��`F�%y��w�gH�Č����83+���!톰B?�rR�v�رJh��U� ��TpĤµ�4!�CY;M\��=ܯ���TNE૸"D������XB����HwDq:�A�ŁJ���2�o����%�h�B���`s�y�����jl*�!k
�H1Ж���J�IGv	mk���Q�6��PG ѿ5:�O ;<����T��C��G�yP��6D2�O�?�ke��7��X/U�s�A���Z��~��p�a�a!�ȠE*�d�40���7���u2ROl�J��)x?e��*g���,Q�D�������2�%~扇�,��*��'�W.tl`As��?���i>/�B�ey����Fӽ���&4F�ŝ͐)ڹ���������žYf��A�y�$Q%��q�$}}&C�� 賀�|Ş=�����s�#�h��C�����̻+.�Z���l��IRQO��?r�͠SU�޵.�����?B�c�S�0·#>��e#,Km P[s����&�F�hߡ���yR	�)�o�ٿ']K��U,�ak�����b{�Ħ8�b�Xw;f7�
��a�)�F�,T���Il���J ~')h�&W�=M�����|a��j��3m��~nbY4S	2RB���R&���ځ_���Ɂ�7�*!��t�H��V��7�j��������"ڌ�:��Jv?oѮ"��P��?,_�8�4dv�����gO�E8�?.E`�w�]�|��h�N�d��uMp�m"�L���Q&�f�{|�x���? _����>uRl��hDCgI�t<S�h��{���Ex]�9s��c�hQ�C�5f��;:z'm�E��	���!Y�n�(V4�G��t������e�(�r��A:0���_��˞��ʾ�(�DN����L��¤��Hۣ�tDzY�'�~EZޜ�k�z�T��]��_�)���{�D\�d�-.�&/���̕�+�u���G|����/�V�ئ�05�5u��&l�uc��݁E!�o!]��2ӑH2��5K�x������}��d�B��/:��*��������B�3�hfQ�fh�G����ٙQ9<�K-*��n"3��UHl^���89�l�i�'|��G����w�P�k���&Q8�`��U����8���� ��<ٿ�`�z�_N�4 	��O������ױ�Y�Ǉլ�잘!�9"��-�g��X�%[�������9b͡�������G�!�����	[j���	>��,�.Q���b��$��/���u�	����x'��=��癪;&�>�2dr�P.^��Q�),h��7�
2]�Ip������{/�B�����)cקf����|���}����cww����~��-ꃡ���x,�ހ?�f]EN����A��0&%�R.��
�Z�7�E��@ �h5�wS�r�]:b���]LޥV|��"(�9��z�J�ߍ"F����G�@�Xɻ�H+�c��ʹ�&�P�up-Ϗ_������s��հ��g�j2��(l (�؟85����S�S���i FÂF�V�t�9��tB~���P�������a��d�c� 'ɱ����upQeK�!L�JM��;(�f�u�F�쑯S�R���$?��MM���?$L�GA]��eG�[pw�F�01�O�������r��2��r�B8��2��⦌m���8���o�r�w�C���"����by��/�PaQ����.]z�X��������6Q&6���v'F�މ�ٴ8IX�򫾊� u:n?��=��~�-ug5����$���9�-���87;i�1D.+�<��B�\��N.��j��1�X�O��Cf��1��A�x �o�n�3?0��1 ����YM?�#A���(޻�|����-���4%���:\g'J��F��#:�w����H�,ҔW!	M�"ˡ�ʁ������Tm��C��	q+�-yW��6ٰL:�؄��<�}
L9�2�>U\r�y��Kwӻ�t�؈6+r������E�|�˸��Ee2��h��3D�HE %@��L�r5t~�.c.z��Q�XA�����F�3��Z&�=����m]w�W���k��b\I3MxpzBcSv��܁Ҋ�1�t�>�[�p���e*�3�_*�/G�������/V�1�Pݢ�l�l)��RcQ&s%�nF*��F8�AvI,?H�h@���D�l8����0W�0�U����輗��Q�83~��j@���"øKɈJB�MG����@��S��LM���㦃�3YsF��Y��H>�V����G��*�7H��+-"OR��t����S���gt�I��A�h��cF�yn���ٽ쌸���VV٩���&�oX���H�h�%98[Y&��Z7n�(�t�J�jc�lܶ�}�>A{iGc�`=��a�9G�+\'y�м��ĵ�zO�C���-�Ӱ��m�u"M�l�6mh�q�d���i	q6��1nv���UB�>�I	���n?�5�d� �lp�j�"�)T��~��>���II{镡�g���	�t�l�FzW��E�k���~W��I�M��!u��<�Հ�D��oz�R�H�1?�ly�b���k�J�᥶�5"k�]��u
k���D����式=ɝF~��)T� �R� b�'	˱����Io���X5+9k� ����������x@d;��أ�V��L���*˔"~��!��`,��)C�k2�a>�#
8���a95w�ڍ|\��_��Ļ���Xʎ�'�g�d�Q��9��#�m�qc���(���c�}��P>cུzs�E�S�U"?���Rv$'�`��.`���]Rc���5�󶥥Lq��#���̾�
�����t��ک�6�6�N��f����Q�v��.����,U�ۯg�Ԇ��񂟣����q�%/�d��C�B�ҡkŐ��*�����*
��uT����%`
hH@�,���n�7$TT�0%g�6����p	֕g�=�\�ԮG��m1VAA�[E�{�b�R��q� �8����aB;�K	��ƶ Xi��x'r��h���Z��������m��hE!;:���!�61jF?}0����"Ǌ���D.* ��*����rAś[���h�-xd]reTd�B��U�k�'��tW��!{��tk�tʄЖ��}ϊ�,N���Ʌ-�����ˍq0�Q��#_~s�Lx���c�����d�VU�+�>�1�`�,�z�Zlk7�6���r��w�5�E�m����g��Z��b�����sȅ7�\0e�.�"�q�s+���(>t:37�`ey׼�<YA������x�m�q�{��>�x��w�oN���f��e���X�v�>�7;�6U��^[C���>��
v[��$�G<�������H�����n�I|�Sj�^A#�\�>����V���zN�1'��d��;�u����aF�pͅW<�cЏo����7���z't����Y������������ǆ�ה&�Ќ�h��{���,��3ʺqixZ��+xT*'�b-O��C�i�@����FYZ�R�1��ǥ�:������"��(�r[�+5��h{{{�Y�#��i� P��Z$�<�#o)Ϣ-�n� .��[8u\>���~�A/ �(M7����ȳ-W7��{����ݨtΕ'1�zpW{'��S"i,�����ΩB��*�� �lI\�V_C�ZqZ�jgRy40�qP����ޔ��δ�L���3_+@���䀍I4p�:�#�Q.��ЮY�E&J�σ�79�xV�'��w�t��������C���������Si�����K����[�=�xt��q8�����E��u�ޮ�ReV�������	$+�[���w^BMp��*���{Pb뜔��}��݉A��j?wZ��p{x4#�s�:qx{2,CFi7R��ʳ��<B�]K���̎
1��2�V����{�C��"v6y�9B�]�UD�wN��T�p�S�ި��fh�M	ƣ~��@5oƩeF�Aņ�A5/e���׾��v݁�Y�cQ��L5(KJ�d��NA+��؍��fN��$i5o��Y`����B@����j>d:��B�SH�PۭT1U�>�	����>�s�u���&����� O�p��y!�@6�R!+i�6�����[ٜ�,��p։kh\x�p�Q���:v!h
��7�ų�i�|�
��2���{�}����;*� ��Ϡq�/�D�Ͱ#+ӵU�����1ֵE��Y"+û%�����ow4� �)�*F�?ix�;i�-WX��'3���wAT���h~㼖�14Y�T�_�z���poG����+��խ���g����{��ݸ9=w�@|ɣ�x��u�Wh��'���E�>��
�Q�䡅��d��9�}d_��	^ٵ�)��}B�hQ.���2�"�$J��ࡾϪ���7n�o�EAƶ[���m�A9�&}	9�%���m���F�u�>H�$F~�}}A��Б#���;�g��@`SaS�%���	'/Q����������Lǈ}g7��B��M0��b�G5�6��Zq<sm�G��7C����^.>>�i�b�
�k�}(/��47b�/E|Eq|��Jȯ���� ������?�Ί`S�� ��. u
|�5kw�l�Zx�
HBiH�yy���6�-���=Hde�TV7:�h�������[�R������� �h`�_��K����8#L�a6�h��=W�4��y��4�{�/�p��\o �<�O~��t�j7�/�g��Ptâ�T�h�j���� ��Uާ�Y~�ۭf.ir��&�B,h(�Q�3�)�E'Yv����Oa�6����Ą�l��u�b%)�f��Bĩ�L+?K~z %�9�*��-�ѪF��C���_,e݃����r��u���Vf���j;�U5��Ou�;_�	���S�B�[�{S�
��0TrsQ/�栣�W6S�ۢ�PG����I�������G*0����Z��{��TD��!O5�V���+��}2�n��3Q2�>s{��S���� y��"o� 'ĂLK���Q�����p+J��S��J�E�"Q���P�	�H�%]���;��_�F6�Õ#�0��Q�$�B4y�3e�o��~�Oۄ��g�.ˢFg2z�O�g�-ت=X�_N���%�&�<+�F��aAb'�H�&����?.����p��Л�΀'\���m���,�>�(s`k�Ġ�c�d+�^���,t��2�Md��_Ȅ�bI�"c�6|�Hx���G����~���e'����N�252>G���;�e0K�e�����Z�B�0%_�����'m���U�x�]E���{#�����5���|pd.�b��j:�+�j��f�'�������7�ڥĆY�ʸ����=|B�L�5�ĝ:�|1���ܔl�p?��:�z&�|���3�3L�j��'V��I����t�p��蘆�N:�.����NJ��:�c�5��ɿ��/	re�"�F�p7��X�����1�u��8PU�;��0���Xks4Uu�E!ߍ0d�M��G�6��6�d��P?P��W���Ɲ\�Cl����lc�A��t��L<
 p嬄��l_նp��EuC��n]�1����	W��Q����q^)ʏo1�eGXML���[XT����yǇ���2��ڝ4�����T��e�E0[��m�B��5���5�H'92a�/�tk^�Z��x�y|���$��Tɻ�]�L��߶?k=��p�� B�3E	��ȿ^KA�կ�>���V����Э�V�z.��������.��Ɲ8�	F�Ճ���bˑ��U���-��nT�_x����fQ�%�1�������?K��zw�����/�蓇u
�mz�$�������W�@DH�y.SH��ndP	/�5���Ur����-��h�R9~�Wt(i����?�>��n>�86Cq[���UVA�e�B�O�j�����%�I�sh�Yx��iw��̦������ 4D�Ni�2f��Y�3@���T�m_�y�O�Ս#�E��=�P��Pz�=��r"�q泏�J�|{��8թ,�2h<���WATSs�>�9}jL#�)����bV���:si�鲭�y���sH��uY����Iݶ�r�в�����IЎ�&	�@�-�R�Н)��`�/:`��|M�Gv>����
� �gv�R��]�	o�tOM�2{�'Q$*��)�=�k�P����7S�)��c4Z��8$%�LS�@z�H�^c�/}�N�+�g.1àì\�u���K��3H��E���U�a
����^Tpl*��z���􁴽����c�[I��� r��[�&1�j�~�$ĉ��O=���L�d�$���刘
��5��˳Y3z���&?D��4nS��4>i�{�
M-���B��Z�K1�gS���MtV%�8��c/�&j�5�W�Y�<�Л�)b��Z:�����YqY���R��/L�[,R����hxj��@K"�����B$'��ȼ��ci7-��@xm�sBZ6�[<�o�ed��g���2�|�����}�����.^dW����g>U��ʷM��c[���SK>憎���Ȱ\S[�`#�}�X�<,Ү�Tn�C��a�<R)�[+��Qu� �AF�|$�Ə+"�U�%��C~�rfr]9��Щ5b,q��9ن�-� �-)3J�Zo	�1)e����}���L�[J�W����(y=��\�(�wi�TI�v�݂�ʧle�&ő'�^�����64z���5���WV<���l��Q\�P�s#R�����4��*�O�NH��JRB밪y�k�,F�>0*�	W�`�^�55�����yփ�.S�9h0�Rte�Ւ��?S����8��9�c�D�/[.�W&�{Z�>1���/	��+��0���'+oD�����P'�w����F���φ\th�$��$�_�!�.Ճ��Y<�o��>��7�"U��&�
�Pe#���ۃ0;�$@�`�$n�̓���X��d�k}����_�#�;L�d�rd�<݋�3j܀��9am6���-â�-��{����>����P��K��H���o��Iz\�Uc�'��d��HG��������\D��L��7������t��(wi�Byzb�GՅZxZ;#����<��γ�����ۓ�5m�g���*F�\:����&B"Q������b��-0��)Hq����98:�ZpJ^2R�5-D?�3
��\
G�<�C�ܗi�����5Y� !Aj��6 ��9k�"�'���`�$o�6�����-9�[�2I*��\$�~K�U������KV�"!�l�?v�#�Y�CP������N�㹝��ե�����+@���A������dh❅�}���;���{�/�q�!�{p��:���2�?de�̓ψ����C���}�)L\��x#D��*�L$�6�O��hn�%�0��.K0N!�.��M�qP���肤�p�M��'r\��-���TI��!ܦs�"Q^����u9����ՆQ�ZpujĕEg��m������g�8��'�%��J��D����-��)P�.��ܧ���?ދz�DmL��AOЌ�?)�J��spOT��m-���L���l�~Ց�L�I�x�Ϝu�׊P�sH�W��t.KĪ�>�׶�� ����Ͼ=IP�4�2 7���e]�Y�u���X� �a��LM�6�c6ĳK��.��Z4�b�'ڠ�]�r�C�VJ6|���TU�A��'�/�g�^e�F�(��h[�ʡ7�� � ���& ��(3�8�j�	1�U?��b�*��p��9{�����̗H3Z4�h��"1�N��ZG�'m�qZy�%+UvC�"�`&���[p"��c��Oi%�� �� F��0'�ӂ`OB�q��=at݌@x�G���/�S�&�oS�������!&}�[EP���Do߄9R���҇b�t��|ɟ�J���m\���W���}����0l�@>G{�e'��l��u^�k�Imv��N3����z���/$l������'n�`���z&Z	3��x]��2"�9')�環��g�Mƅ���X���9���ľ-�l�5��!�	�K��P %WJ��}�{��������ݾ_=+?_"ᰒǬ9�ߛ<-bRA�����5H� �d7�R�E��)-3��"�̔���2Q���t�['&����T��O�9z�xw]����@��a�(�Ыqsj�"�@v��ca�Mx������ö�H�@�GfZ)���Y���l�~�V�CA��f2sy_+e*(i1�?r���$��|�Q?�����&���8�{�wH�^`��l8��\?^L �>P馥mg�(��Ѯ	y���r�#U��G/�Hr	���:���6���}�e�U����Oa��\DH����o�R=ցqrW�á���q�F����C��U��`Wyqx��6��V6��Un4Ȝ��o�|ꏄ� ��g5�7S�s~6UY�����h����?\h��i���+V�8D/�4T"�U4�t���!&$L���܏9��c�ݥ4�_�	@F��ڠ'��K��8�L��+�(����r�.���$^<��u���Lm�&Dt�����^�vU�������\`��R��R\�
q�B����3R�*�$�)��ΗK�;y�)mO���"
W��=z�8��r>s��vFރ�>��?˯Cj��K����r=�� l�޼��6�Z�!y�,�e�o}� ��_F�B8��A�#@�`
H�,�a�cA(�P�2ؓ'[�g�\s,۵p85���sQ�-�Tipl������=/Y9�%.h����U.+�q�Ï)�X��#�Atp���� �i6% ��/�t *�;�P�f��d��G2M�4�2Byy����`{j�6ev�R=N�q��UD�n-fR��<��я�D�����L�ٜ�ATZ�߆�>�s������fz3�� ��M-���J��
b�9����+y@���e�|�N���u��@�'5�MP�7�� �\qTl֕hL<3��<����Lb�!�TAVP)!�Y��p����g�\�ܞe��i�a����pZ��}^�9���k�����&i��]����$�U�'�{n|]��d'E_�$��)wG�9�nZ��v6�� �oY7"�	
X�V"�wZ�@s�D��}nre��z�34ms�8]=�2}2�:+˦k���$��`��_�����8<�
m^^1���ڷ��Ĵ:l���E��}��{4EH�D���!\�NM]E��G�u�{�d���oY���D� ������v;N456]ȃ�XT����	�I�Jg*6��q�=�"���y�ap!���%��+B���R�����}F��bDd�&���͌�#�j���Gg�O㪤���k̾A����1+�
����+������E��eZ;V��F1�+�L����H���Y�Dۧ5l~d	 �����^@k��Q<�BĹ a�d������4�4�QR�hદ<h���+�E���s��D���b�@����O���f���\!�K�-XT{�(:(��]������D	V��Qz�ؾ�?/2{~v� ?���?3��%�I�\pM:���{���ͤ+OJ�*p�5	�!�o�����.�O�mR��d��XD'�:����A�{�:f��XbP&�9��1��4�e@b�U.��E$�{K;�}����B�']���+R2��y�����t���"�[a��[������Yq�,���U=,�������PS֫����.�߳iI&k�L�.��f& :tZU�*�h���Y�9��DOv���U^	�����]����4Q=Z���l��X�^g���Y��Y�m��� +�&9��e�C-�0��{�@�(ٺəG���X_��.cԋ������;����Ҫ��������+�c|1FL�} yr�����C���`����ȡ��CU�2y�I7��g��-l3���F"tC��R��ir��ĵ���W�:w�Y?��0ҥi).=__E2^��ە������=LCwՇt����͝��k ��������cQ���.ڬl�,���Ϝ35���M�����6�ٿ�d�IV��.P��:0x�8F-Qi�l�7R��kO"��.s?8�ҧ�"�Zgܒ�R�HJ��;4�	�`1�'�� lX��q��XW��n+���Ҕ�=��>����X�:��}�=�� ������˥�(2�Fcǝ��(�n�^A��:0_�ɋ
���f���U3���D�i@����1|$L������j��^�j0�Ä�4;�.���v|� ��`J�ˡ�7v`�h�$�Ǫ�*�`H�*[S��
/c�GC�T��S���ym(�M��7D@�`���E��,c�2|�g%Dk�;�QG���V$1.�����8>Hq�;��܄g�)ClcF�D���n���楇��^T�,e������W-u_�6��_�Nl��u˯��RŮ�틱��-�� �3@�5-{;x�*ǎ���~���ܽP�L׺nnj�,:
��A�)g[���b�6 S�	k�+��T������O�3ni�J����Ŷ�)��3] ��"�ޟ"
[7�>f�����&��9@Y�>��:β+���0I���C�Jc��F�`)�;�NU:6V�W4�t�Q�u-�?����"�}��G��Ѹ�ų�չ�����KO����� ������@�bwG �
`��OL�$[��V�T�	�H����"	[Ѭ����mo$�.�nK������ߑ�F-;{��&uI�F~���z[p��l���ל�a����X�	�H�3���#��g Iѹ�om��k��Pኁ�+���E,�����א�g�^��M�LH�n暮��P���:@��#��^�"���������9������+���H����d�؋�x��kJa��Mn �*�6��k�Ib�L�]/x=x��C%��>�<y�[P�.�J჉�f���}և�zݨ�-X�3��hƬ~9�����c��?X3e��U���8^�"x"DG5~=`���J��p�p��2<�y�o����x6ʌk�f;���<�S
ō�S/o)�T��g;
��f�3.�q�J�D">͵��ա�6H��Y�Ty$�����E3�k�2/l�g�p���h�'d��$�s�@<|n}��p�d|<�����AnVw�u8zSrU�΅s�N법��_O��'������=����~_�Z���ߗDa~8�k�4������nJ�Gu*��0S�s�G����?=� �,@�@��lO��s٢����[#���?��,	p(�t/��4�c�[�^���5�V���8�T��1���?%��K��7��ƭ8Q6_�d;)ع�ھ ^E
��r�����$���t�9�I�6dh����q_Y���+v*ʃk���rb�-c�k[L��j8ys�-o��Eu�[��o�Q��T���j��i��n�FTز�5��V�����C�þ}y;<΀��`ir����*AGrkG�9����^�783B�����`�o���qwI����<ʳ�Q������������t~=/�Sk�|�sLe܌"��f"�l����-~��%� <��F�e"@T_{�boc�D�4���ڈ�~�c�C�����m�M��7%ѕ0X��d����n�3x��}_H��"}�F&����͚��g1�r/e�N��e��[N���ӈ�r%>�PA�	@��
��<e���KNt;����SL�QΝP�F$�Iq��!r��PO#c� GZ�R�PV���4;���-���['��/v�8lԕ�MC\��M$�����gL��Hvsa��l��!�?l�OiY�'+�@Q�?H�{ItL|����7��u˼b�U����Um��Lۗ��Ƿ��,ӈ�Tm���vC��Cw�
2{�@%��BM[��G�J�OS���-ܷ��s=SEZr�Z�
|�$/vɢ�t5� l+��^?��]ƈ����<�[ٺ7�;�UApOT�r�����˺����ݖCC�fȅ����_$w�Ǥkw��	��Ю�����"d\�����}�>�;� ��!�n�QJ �jC��
zb��ZdX9@Oc�1����CJ�%;��/D��Ԩ�/�H�_��w+�t#Ci#�O,�F�C���H@[��`��M�M��,�N�D4,؊Y�9����G�����V�����v�Xd�󨽜_�(Ml��_#j�A�~[���~��/H��h���Y4��Ժ'l��#HW�I,��{�M)��7A����F�����.�v�Ck�m*~��j��L K�c2�6m�?�#~���I�ufX�� asg�4�������Oh�w�	j��D����^7�9�U!�����݇���:�IiU�owIt�Z�oΚ�}>�V�j�z���=� {C�s(Bm5:1r�G Pp�#�4�<�)>+#O�^�j'�~�9��D<	����K�úr�#	X�*�FY11� �=�����(?����T�*Q�8�����i�}���=��&�=�>u˳V����[�4���J�g���DZ��a�i@ŉH�̔d�ۺC�j,�a`��!5�� ����H�P���d�������8(ݖ���WTĸƁG�J��wN��?,m��o�`���u�PkOsc6���E�#t<��=6*`̔��6P&Ò���'��Z%}���څ�xڀE�S���*J�A�EGg
�6Z�S�<V��r�E�`eU~�C�hy@�b&mV�������� �Ъ	c':Z�s�&�Q�� o����R����M�~��G�uI��.˿�ØϚ=��s;�L�
�2ѹQM���w��.�UL�1tM$��_F�k�*K������s$���CX���^��mbū������Q=��>���B�Z	z"g	㝘��YE�����ַ��E�j�Qu�jK|/�ԋ*գCg�+4�<`��C�$��q������N`g{��/���J��o�{*	
������$4��|\��5��|%O4�vCn�3�|\�`I��;#Q���9�ia@���)���Avi�r��2��;9�|uGfW^�T�����I����M{r=��'��]t!�!��]D�q	�{�c��5�@�2���J�ne�/g`��2�y>-(��	"�",U����)�dm-����삲f�KA里�=<¾�@�_6�.>�~]B�;�+��.�&���Z�52	X>�!'k@W��r7p�&��O��]� ���m�g��.wy�xY}��^����j=U�\���˅�@��n�b�-oU�&�(1��Ȼ��|%�C�B��?[��}Y�£R}$�?����p�S�7C�4���	�4��rF�M
8�8#��q�l����܇�X��#��h�HNF==����&���6�M��	�J|�4~{��-z�`��l��O�l���\��v�B�s�.�cxW��@l��X�e�5�~]v���Q�������o���_���+=Q�ێ͵�k�X�x����!ˋ{[����2�vI����-qW�^�����/����9lS�)�~���ԏ�� �5�̽�"��19�ø��Zg�
�Y2�kr��\r}�l��C, @����������b���jDVX�J?'�0��Ql_r��A��LyV�Et_Σ�O�81�2+lT��m�=u1��^}2dtJe�#d���X=�,5�r����(�Z�F~�[9���E��&ػj!�:z�ph�����<`K��xD)�IHi� ���9�(��N<��-|��W�hSk���a�T/:F%�n���rl�:��׏Z�l���%�p�ο��S�������B��
�/�a���.Ȍ���'+�[_1�p��U�������&���L�j�a�����ȍ.�}	��?cyozԸ�ż�Fk��@�^}	?0ף),
OJu��)M�[La��4�����p$���}�,���-�V�o~��VD]�b�*�	���]��S�V[#�$�������F0�1�7�P�̽�`1~��N�4*iG�	q�����ث���%��"�-�oK��`B��	��&Z�\dmF)�Z�|��R"��P,:
a$?vqh�F/���@4f`�[��o�57��J�(���	�FkO�)P�n�U�ة�KG4�%9]@�4�V�V�*����z�0/(�-�����2$�_ ��5�x-AȾ�}�1��A�,�-� $���q����jG7��/R��Q�4�(R�m+c`�-���zt\ì���i��Zv��+�e���ƿ����8v��<K:��W���㱮�7#U��2^�y+���Xzc���-�F�@h��v� ��}�k^S[�V�O.  ���i�V�@��,K�Y������"��.�z�PX��":�ўz��Ŵj���1�G62�L
o�O�K�kC�@m_�a�8��Sy@9���!��cm����w�L)�:�YIZRiM��~	�"�����.�:0�O/�Ѭa$~����8s����uI�����/{�Q/ʊq����H,cC�oI�k>!�+Z���q�^��h�^�K��"�qE�Hx�7������=�Xf
!0]Ѥ�D�c�B+d�������P�H	����x�<��?-�A�i���)���5p���;)�)-��1������c�����&��C�Y��8~x]�O�'.K�j�X���	]��6F}$,��W��r���`��_Oˏ9��jmjy��G�8�����Z/W���w�f�i��<H�,n��qGl�:�B�m'�*�t�8�aDZ1�I���L'ZJ��c��v�ɥ���c�Ku2t�u�$�!��;�W�n��29}�@l7�8�CV�#H(�O�ta�H+a3>�s�m��6��u_2�ۉ0�|��~A\�V��J�B��Է�ӯ�crZD�y~ A��_�^�e�g�ws����l�<[K���[.�����~������Ϸ������O���Y�2�s@9�:?�gB�	]�����t
�;6e�?���Ĭ�������<u��RJ��na;Z�$ �^���gU��r�o)��8�N���J�'���oE�F���\`NU-��;���-�pM��~�5�|P��ǍBۖ�C��N�R��#}YǼ=�#��}/¢N@*\�􀮱������2���~����^q���fj��B�2��$��?ӈ��d��?���@�Vi<S�?�҄�a��17w �k..�R����5Dw�OX��n}��+-��y�G�]�%<w�Yu�3L����pl���R?rl>��D�.� k[��3h��x��Vٲ[F��@�����+<m����Zʩݭ�u����Z9x��5"���Ƈv,��3�v�]�ikf�b�(�i{�)��@��NzK�,�̵\vDX��5E�4��cEC \��eV-	��!��k8�@C$-��D������R'�h���PAt�1P�	Wb�2�
LHY�2�yۢ��,����$�_��"��1�N;RnB��]����>�+�#�p��RbD� �ͬ�M���IӤʜ_D�� d�La�K���LvP�����1l[6����~�CW#�)	����c�Xn�
e�8$ӳ<I�������*�X�H�ݴ�d����6$�t*�����x��4o�~ت��.�
��-d���q�]<�D]��n��O���Y�ӎ�O57�NY����KO%���Q��ةH���]	���"xc���<X���W�!���.��:ww#*k��ط_8�<�F�f.-�'�L�i���b�nJ��C'/��ܻ��R�χ!j^<�?Y��'�b�cG0�
������,Ip��/���t�-����=�oR׬�V�{�p�%������]:浭���-�U��g�B�s�����T�����gh6έ��������`v�L��B� �����1#Bd�z
��ωZ��կ�B.ŊLoJ���^V���J	Z�n�~���[m���a:ͫ��y�u�78d�@�7�����*.L`�_���$ՋE�\��9��I����X5��"��g��a�%���^�I�_���rx��"xJ��Zy}����i�d�ΔJ�K���a�����&ɂ���c�
-�����ՠ�_��ci�	쪉�h�4V,��_�7@�s,��J|���)����plk�K��~��	B�:N���J�27� =t(���8���<|񖙊�f.M�9��������/\�yGu�2(�^n��ȕ�s�nF��������Z:X">��sl*����R�l(y��3��k���<\�p]mQ>�q;�p�jv�V56v�{����K3}P���2oo���я1��#�� ��WW#����V̆&(*� ���S��(��76AW�PsK>��W&�
���m�6}����X��v�u��hc�S�W�ԧ?��q�����zY�K�h7��y¯9$��R��ˠ���?�%Q0tr�[���������4�ch���0��6aA�I��|�c��A=�KA�Pm�>���1XZʹC��}���2f�"	�ӜD?�Wrt�{�6ƛ\�i���F#�lһX��+�츕@7�`�6v ���B�C���~e�?�xX7,���
�=�����'��e�\��:tn�KL;|ǰ	(-Y����Ϸm��ƴ������־��f�٪�D"��NmOt�T��VOY�f>"�Yj.)>�9j���I�#�lH�ćOC3e�. .YF#��B �G�h�K���t��/	t�T��<D\ �V}��H)�Ɵ�%���k�w���\-��g�(N�y�1��ŉ�����SRmU=�f�b7D�XZVkߓ�i;�aL?�u���w���b�| �_�*�����L�*ԁ�4�ӟ�#��+�,NK��<÷z+���x�3�[`��Sn��������Y��a{��������{f l���.B%���l����
�;va=��\�h�gW�u^��������pR�[Bm[9OBbx��B<|Q�	~[4�q��+r!���Z$=_)����ָm���胊��]�\AEx�V;S�@��8T�x|*�,�6��c�o���m�?�s��6���ֹ��x>"�[x�ع��zxx�t�ZAd�"Q3��֖���[o�� Џ�~�s����AMR�KK�ڒ�Z=�����p����	q���+ӳ�ީ��u�����`���["AgS��VΓY�A
Q��?�4���fp*�$�������6p񟩢dT��᎑fP����$�9s~҃�ܶ�;r�5�N��	������;�O�����)�V����P �n��t���K��P8p����9#n'��$Ym\�.t�?!`بj�\�A�%�*�Oݪp���3z )ǒ����B�]��~z�7Sn%[��	�$�en�( ����Ӡr@B�R���8�O+���yB�Fk���l� �܄�
����Sr8���H��q^:rsy�W���zø�������t(�wW�I]��S?��P��Prk6e��jsf��,���q��@�d7p����hT)(�ĺ{�˸5�v�Y:����7�òN
��[͎k��2ab�Zv}Y�^�ikP��3B�^�1��j���qu����Ə*-u�dB\�(�����ӣɥL=*�M{��`�f����|�r����Q���sA��p��S��:�ҹ��(���%Gg9�{a��3�if��rl9���J�f7=!�ꎹ'k�W\��.�������� ��Q�����0��^P%@������b+�n/a�	�Y�Ucv|��(� �y�f�`�-��i�l�\?�c<�V�4�O�'� �ϟ�d3�;����9J�k-�+1�ִּ�k��gdA h@0�![�!$
?��C���ų����I���詀���$kV.�!e+�+r�Gp�t������"�l�-uvX;�Lk�	�{�K"7�-��^-E��N�}�0�U��\R]��\lk�jS��W�ݖ�LM�~L��C#�Ǆ��"�C������ �e �T��xM����tɬ������y6>��Q^C4�/�6���j�Z0���b��Ӑ�3�T9�^*aX��	D�m�q�A�Oe�����6���w�X)��oA��L�G�9�H��O"b�7a=ĩlC�>����A���ۢ�d�YJD'�!���7@�M;'L�"ud�ޖkǚ�<5�$x��W�֧{��o ���O�����X1ڨ<�k,�R�ב֙���^�����U��t`ԕhC�4i�o�ap���/F�qs����IQ�
�[��Q��'l�ͯQ3Sش�C�������hGQ�TÜ�{W��%��79p�WH6�H�Rvi��NB]�RDJ����ف�J�Ԉ:�`1d�����$���g;�z���Jm�t��p�d��tZ�^s����rl�9
��=�U!�~]6��|'�Nb�.�]�H���U�܌[���u���p���^�u����4$B�v�^GƎ,@{��eqj=�~"��\���Pqyi�sq�
��v�$C�� ̋{���1���LgnnT��7_��ph*D�L{!Xg������.'��dy �2UL�%�n�ĭ��op�׈�H�
�Dv^�����\��h	$K<��S)�t��.�Uqq��f%�Q��4E���a�d�� ~M�4����v	��C������Z�]X���Ɨ��V�e�l<���K�V&�
x�1<%RW��ĽlPu�o{���$���.��%-v�X��pmx�+!�����<�T��_AI�T�U׋%��|�5W�9�<���0��+���B�}����%b)�b|4�jJ,W{�;�P�����B��6����Iw��S�;�,#i4�`U�C���Ȱ/��4�ې�����c>L�V
��G^�U+���6�(��pK����6�&8a�b˔����(1����
�<��ݣ֬)��h):��ƠC�T{	�a�:F�����Ѿ�\�8�_�#�?m�_�H�0���1ΰ:?�;���u5&G*�}7�Ģ��#N��0���2�%��=����,�]_:���e���c�m�d4�d-a`R�55��pN����9���\���Iǟp.��:K�Z���]/"�����zd\�<q�)C�;ɂ"X��&�=1O,#�)��sހ�&�b:}}�x��(�K�Wg��w��pݥf"2d���aS�Y��-9_�D0$����pΨ�N����R������B�P�7d�&�O��)��V���O�FT=��,�?��݄��X�颈u��ˠ�!Z����0G\J��*��_�x�ܜ>.�[��K���i�EP��H����X�YQ-4u9Z�i1���v�_O�"ͬ.�G3m�͎ʺ �$����A]2���=�?!�Lߡg뙠���4>8�ыWGe3��)E�#�j�A��J�#��7rMV�����i�Ľ&��C��y�$.��Rx�
@�2�� ��*������t��>�ո����O*^o
ڽ�_��G���h���'��b[ˈ���Ď�֤�m����R>a�2u`0����ȕ��5�@K��}0M�l�@��@�c4�����~��*�)B+߳����y���r�7f:�[��k�f�؈m���f�;x�9��ͧ�A��H>sb���#P��"F��aFK߷���ZDU!��`"��:�53��n�x&7�|�j���|��/�����㛀��2n�φ�笅=d�i;j�ס�8��P����'��P��PU�}�i�J����֮�2A)l]�F�&-bx�$�2Tu�H���#t�N��HW��ZeB8�Dt�s��m���S������fP�Y &¨��IM}Y��)�M��q-�;��3s�\-FW2˃�ÍX�`���L�Y[}���X�Z��4�h��l1��خ�=��.�������K ��C�
��jLa�)� -<���J+��.���;k�S�G
L�:�C�2&n
ڈWB޵(�՝�0WH'�p����Ŗ��p�t�ᔱW������dç�.�A�K�J���Xu˛�Q��ߋ�'���(;�z@�o�;*?�rH
�o�K��h�k%��f�`U�l���J�cm^�����"H��C9�Q���y᏶^fA�)(���s-j`��ƀ����k�~]2�m�A�[������ӳP22E��k�w��raN�Y�������f�����#}���:�dN��$��n�G)C��K�KI�Aj�m���kK�kH������T{B���,M;�k"zГ4:lq�>Ч[��pTF�Jq����+߁U��dN��x��ɿ
����N�0���n�d9�[H�ؕ]��т#�c��aĂ�ȓ �����=ǯ#4�̆��@��¶�{��]�����!���U�������囗������U@�H��JvDxq� )���ۗTP)Q���#*��&����a�o���9�{W2v̞'B��z�#��E4'���	��}.·�XkF�����DS��)8�� AwL%�̇D�aw/������5��n����4�tY�$�>ET�2��!�x(~�G!� g�4$�I�YR�����Bg��4�4:�� R��L�pn�K�����j{"�aK(@	���A@�t��OG
y��/: '���j;<���/���!RW|����� �;� �ټ����Ayу��s|-��"�>z�[���R5{�T	�TK �a\��(O���o�d3���xv$Y��#6�A��q�G�A�H���y�G�|
T귡Ư�څvs�M��W���(�h�5SS�lu����ׂ���	��kI}Cڥ,��U�������� �T�>LIi��B�Oh�֐H�J�d<�۵<���jf:Hր��JqNv�rC������]W�Ϊ�-	���$X���`b�]��Q�3ivqox�-�4#��1q�"��]B�|������K���nN8���R��C.?���!1�=r=
A�o�,�4����떇v�0a�OO2�"�o]՗N�n��-�~&x��lA,��ʹg��$�'�h�+/cZw�˘�5�jnx�u<,X���U�*R�)�n��u���d�21%#C5z���
��A}�[_��{�G���	�V�#��`M�s�2BhH��Q�����p+�t�@o����q������GoQ�zy�+]�G$��/�.�z�Z�ud�#[�2���Д�@�@� � �</.NR�K�[M�1�P�[ �k:�(���qaf?n��c���QW�`E�D1W<��m��9J3m�n�:a�����o�:ˏ�
�=X]��1�|�ծ�=�� _#�#���'�r�Bg[��I}��I�>���x���T ��g�AJ��G�A}h��PtJ
���d�D9;���뚹F��k7��pI��f�`l�L�,Q�Vi����LȬƒ���zCTV^߷�� �K
��{I�2&�rB�Z�!�Ȩ�-v[�A�1V��֋a�f��"#�sw�-�%|��J���ֺ|nH�o�������+k�w�RW���
�� Eq��_Fc�g�T��/4�RnN֕�@��J5�{���΀p�+
�)���VeYGh;�h[�<�_:����ʶ��[�S�ϝ~e.va'ո��b�$+��e(w�4�T��3�U·��+5]i��O`����%(p��0����^�$,։p�:ۂ0p��ר�P�#J�m��A;�`c��n��z?�YU�AIV�e3@�%�LM`VD���5/o��|\}$5)s �3*)�H0!��s6M9C��M�AI$�)��)��6��:�O������&����U4�f4WYc)���(/g6,5��������t-�yK���O����ʌ�#g�N X��Bn)�Qk�D!���M�g0��? 3� �Y�����^O0r�DBoM��U���:�VSΠ��lT����R��
�0R���n18HnG�r�X�W��	f�ө�^јcY-0�<�/+�850����T��
��M�%&��iYV��o3E��2j�Y�e�)� �xp�d��dT}���Q`��� ���W �%D�H[���ٯe�g���E�e��:G���M��,���R[�;�[M�����_���i~�K��w�5IGt﵉n; 0��d� �=WQlx��b�qǤWYj�P��R��������/+p.��[�C8@m�}�E�*{rD���es�)P���y�ۤ3�L��x�"S���g�$�Tڼ��R8�H�}����<�0��ª��aA�<�;ǣ��^3Ա@�RFW����O+bb �� �.�JM�KJ��K� [_�G`�5K�0��;�!� n��(8�9�F'(K�;�ub.s���8,(�0A��,�R5��mg ۰Q���,j*���&R }�fBJ}z�wP�)Y���t���_x�㣋Fu/[yt�)��*L*�?��5��FT�3�쿞�ЌP#v�l�O;u�7����W�{���O�窛ڢ�����K{=wlT7]Z_P�����
�	q�8��*Cf>}H�*'��qhPP��]h�c1��]�N�(d"��J�  Gq�Rv\s5F�M�5d�� g7�C�x��r��[�.�f���0O�_��J�G�X���x���L��~\!p��Hjnc��1��R��j䥓e��ԗ��4_/Z�
��:Y��e��X��Nj0� ƙ���jV��N�Cd����'3*)r+�s��4�5�*HN��N�Ȩ�J278��!z���b2OdDk���������H��&�l�����^",0�l�`�7���G޵�w�|b��-�E�B-�^ y�@���a>��&�7�[�Y2qa8�
80�Q��N���:��Ԝ%��]}iY�O	��Ҽ����"�o<�'�d1ߦ�b>R�b"F��=(ӱǁ{��b�;���04�����7ь<�������?���$Os�Ϟj}욾��  ^i�ߙ|�ޞ�0���V��r�T茙��yÜ��b�
���絖4��R$n9qv"
Xx���S!��Z�|�3���g�@e�XJ��9�-�M�j\g�Ytd-���_o�;�e�M�A�qR����Oϋ4��W�W�p�֜8�vpI�5�3p�nĴ�i��I&&�{��}pw2d��=�4�����R�x�I6`�f�ԑ�[��}M�1�3go��#X@C�rFŲ������EbtG#%С�vh IR��!�}Z�u�p9J�oK�I�n��-$�����Dȗm�h��3��3�^�#�rV1���7�O�Wa������ ��mͽ���3�=Y�y�S%��1(��]$�i��.�@����K��B���,�p��1/�<����k)�o��Hy��������r@
/t�}qjY*1u*4��^S(	�胄B�/_wj\<	<��ή�j��0��Q:��1�h�J��8��e�zf&!�Po���nd�[� Á��]����[��D�����^ T��n���`&��D7������/�>��
��I�T'�Ta=UR8��o���?#SC�1WuCI�z ����>�3j�ڤ�����1���IB%���F� �#�Mk����^�h(o�uĦBV�Z�fz�T+�E�W^r��>Iu8VWiU�^����b��P :���,֋��E2��N�������ȯ����S���>=ٛ��=���4FB�ё5�Z'})� �މT͡^eJ��P�B:'\Z�p���di�`!�@���Қw$���=D���	�Q2KFr%S԰z1�9�Og�h�h��]�0���a�pT�����c���.�
�~ \*�iu�����M�G�%���t8�{�0����(�����V�u|:X׫%g�7�%�'2�u�(s	b��p'(��d�PJ�Efެ��������4q�Bz
�X�}�~�Xբu9&���L���B���BR�j�{ �j8�을�%O�ʯq.�~�*\�چ��[�h��2��73�����3�<�i��/͝��(�V66y���R]M��c±���T�G%�;̖ˢ�h�#�'r����Mn�sʌ���k2�X�i?��)�']
�7�\�=K�9�ݠ�c����D5Xf��<����2 =6\��w��ኣ:@j�^@^R���7Y'���-dQ�#R�e�9��.�>�7Jx �_�%v���k `����%V!���m��|[���]��al����ɧF�fn0���x������!�d���֙k�̈�����F��G\F�bu�ը��Oct�1 �x#���r(c���͑ 8�{P�p�D5���7����n1<4�����U�ގ����X�o$����+�΅G�k�7�b�:������á:��t�%�N�}xq�\�,�'�� ��K� Ij��Ts� �v_!��{�K�Id��R�yK7~"����#1Y�l��Ƶ�K��1.S��X�RB� �w^��Q�R�̙�1x��h�F<o���������A��g}���|����(C}��Md��D���Pf��F�^�C��d��I0a[�@yd�8-D�{���d>F��g�M*�&�����,��(XG4�曋��XV�!����ºwf{�~��ѱ��a�'�i��,��!��n�����i�n�(e�:�)�mDDo�~ru��AM~u�Ø�,6	;r�aգ����jL�'��7�U�x��o�W|/� $ ����Q@���&E�L_хIU���l@�i�)�w&ްn�4�S+i�T��ԟ5	�כ��e������q�w������h�ֽ�d%/��!ƅ��.E�ߓB:�,?�ѪQ��������'�C��z�n����Aap��5�uD7�h������辣U�����|~d	p�2��3�UL�J����ހc�µv�kK.>�m�ȫL%$�������9
/����D�d��UW"l_�_����Ȑ[An��6�Y�H<�f:��?%����e�p�f���o��H�iC�-�{��ֿ���?hE��+*h�u�;�������z@�R�Ȍ���������g�Y�x�����X��`E����.��E�Mύ�Mvܞ��d�����(��5bq\r>E����^h��x�so�k��	ʺ�5e�MJuj!j�����*Wq�5ߡS�M �G�_E�ꯢ�O�.�ٖ��&[R�m��Ͱl�|w�y���ܣ���v�vz���28^d�w�^͗�����}���zg�:��;E�"�=$�<���l���0XoU���_u��0���4֙,�1A�+B���A������ �ekO�3��ebL:��U�͝%�"ȽU�&J�4&*�\�N����?�bޥ�8t�6&#`e^��U�6B)J���ii���5�\mrT��}�8̸4>�$b0О���y��z�KC�Enҫ����Y�NV���� 7��}��Ӡ�{�
%��ZI�L�x@��5g����h��w��j�7(���bLB�����_�xul:!֊��Cu��i-�A��·f~��[����M�,�}�.��k%�����"%3��R�L����-x\��h$*_J���T��ӽ�JoyJ,b�g�s�d[�F	��J�N#5-9c� ��v0��]�-�O|�^ �1�:$X�e,��߾���f�%����l"���X�s�k|�BBqx��"��B���k9l�����?�Υf=QՍuq��7�d1�QxR�\���֟��#�9-��3�Y
Ҽ�g�}��,L@�cV�z;	,*�TU�D�J.0s�ӌ쩉���s�#�dYD��SY�;��B/������(	�1�8-��� ��G:�����M���Ǎ��߆�ô7�4�LR}�Wu٬Zo��Յ�f}��à?���a�	�C�M�qk��w�/^�J�3��l��R^��<�_F%PK#��7�rC�Ґ����������v���TI�0Kز�p������z�2��N���#�4 ������v����������TK�V�=y�m�s�!�g����^���-l�g�X�I(�����g�m�
%qˢ-�2૪>������X��	n�U;Đ�13�n_�3�@),Ԣ�����>�Q�:�Ol��P<�j���;��q�@"3ॣ9�;�ED|�]�f��8�v�cwz�m�8e��#>B��o��*8�,a5�=ۿ��$�����g�X��D�[_�ڔ2V"�7���mty��9.��)�J{W:�|I��`
�U1�
X7�7qې���1��k-�u_�<9���OUr�xalWs�1���!E�KG��K���}��]�ǘ)�J���6�xnW�t<1#U'��7Kvk%{n��O�:ѓ)cM}�""	m��"ykx�C���e�[|#VW*�	S3�u9бd����gl�ka4���ǅD�a�����g`k�2D1�ԕ��>��J�9���S������?2.�`���H��k�	���u%�@�����yP#+!k�r�"��y?Q�}.R!���вo�O�?>����/��`��v�<��ѡ��Hq��^fe��s>޾P|d���)�(�6r�+��ڷ�V�e��ٓ�.�p����g��M@���'E�zI6	f@��T��a��ٍW/՜�aD���D���.��S�vcS�y�3�"�ݩ\���R��X����w���8D��@7M(�a`ڦ��
���E�shD3d;��2)�@=��a\�L����¼�c��̪I�2�c����'}4~c�Qu�*@�����ɥ��7��y�Ŝb�]>�/���[�H��*�q1����3N~h.��*�^;����k��M[�	d, P�Ŋh��C�@cj4��s��W	4!C	���A�mͥ�l�Ӕ_p���h!�V��h.>������tL�0�i�\��$.E3gR�wM��op���k�u�Mӫ��o�>��W������y4��/As��>�v #p�2��[�F-ED��z:fÁޤZU�l�Tp;Qv���t�W|~�>'}�S�!/:���:���T���؃������/��<�?O}"�e4`m-�1ͷCm�oL}(�`J*X�w7��u�{�Q������Ƒ���]�a��P��9Ý�;�m��X'� p�x��~�9&94dP�W!���2q|���TBQ��� �P5Zz��A��; <p�ok9oz��p�?<���Rޕs�;�zf�r��%�@h�3��C@,�萂3�e�R`�ֺ���-�5�`ܠC����5շ�{�7��R��(������e#���q��k� Y�Z�i��z?*�s��
}�Q��L�?�����ߒ��S�m=�o������=ʁb�������h=���h&�3�"��~0c��)��b�_m���m���Nw�����D�2ݢq٢֢���l���8Np`��p'��/��ޤN���K�ԄIs��ox恢uaq�뾫�v��_���G�\�t"e$�Y��������j0�W�6+$W���jڰ݆�����&�Y�Ǘ�!ֵů�Ew��}|r��������"2�ЭWK��s�\@�a,��	aAW�e�V�#m�}.�kM\P7��H�=ߪ�p�"M<�����|f����{uj]���f~1T��d����O��������J�PDR� uG �"ƲFǖʪvd����J���Kso9�iY�Lj�?�2��c"�@+}	�dݹ?v&�X��r
>����|�bb�iP��]j$��9Y����)�5��Ȫ�p�|x�y�� �jD=I�w���
�ag���'���<�i��10@�'��x��l�A|j�F��]�:9*� ��I4��|W�/�t�9��*��g���+� H�$K���������~/�R_v�I�ps\�V>���X�M}��g�}P[�k��V;�j*h,��SҤ�Q{O&��s��� ���1]�d�~��_h66:_�sq�*��MO_��+1q�����^^�v�ި���c��gU����Ti�"���z�Bf��l�v;<Τ��j�ڕ�f죯�+@vmXo�k����6D�ql�F�㹽���q���o�ą�K�vu��ᅽhG�^�GK�$�k����2{l����/'X���f6>� v�Б���L�m,c�{ AG���RW���b/�gi��3k�4���W^Q ���f��d؄&��Q���G�5'����E��\����&���|K���������"0�z|�������\!q��v�4�G|�-c0S��TV��m��=��^#�~ᆔ�u�>�*�q=��<�
/ua]��/�o]��"�N�#�T���dXɿ�0v��&l�>�;h0�}-OY!h^ſ�L���:��VS9|H%�9��
�Y�`>�Y�Kŷf1���YqȌ�Uf8���P(�novk��m��Cb:)��k'��g���J3�&D�C�=X-b���e�kA��ٖL�1�%��[�7uG�7L�s�o�IC�#6�SF5��#�Ų(b�R��ƼP�u��#4�����Oϝ����!��s��}����3��z���i�)�bK����]Ѷ�ڌ��,ٽG��|Ж����h�a)��=B���޵?
a7m�X0�F��R f<츪���W�"g�kF۩� �S�|�/��� $�;Smx����ϱ��&k�l��ݍE]�)6 �{"�/
�N�Q���i��L�, H�bDGdH:݃t S�Ѽ�5_8�I���y��S�&�vS[Y�zq9��Mڮ߅�����`a�N"���ZA�{��kT�cK
��g>䐅�*2�Z[�}^� `,�?���Պ[��Y����t��0�T�\�Y���@����A�V7��N����i�b���/�?3+�9���o �������QB����e��D�YB��򰇐ŎI~��Jڀ)��q��y�	F��R�:]$�¿{�����B����~)�{j�����@!�̪'ꂾ	�F���C'ye�2s�`�F{��Bb<�̟�\T��"�4D��:>Y�X��kW0lF����j^!�>�ё]Ź��	�SY�S�9G��n����v}Zʈ͍ʌD���L$�M0�fW��q�tJ��w��ډ�IO,Q�p�tiJ�c*�V���	
��q;(M_������C)���$���$�;�K�[~T��e���}����W;�Ga��s](1H0�^^�Ί�W�1dD^\����͒��2�܋贞�=�c�;r������˸lb1��z� ����v!-��B<��hó��dW�����%qH�E�D����j{�;7������B���`4��\/�O|>�*%��_c[J�|8�=ļ��M����`Ӝ�ڴ��3�{˩��o���T<7J�ˊr_Bv|y|/h��SRJ$p�V �mYp	zd$�dw��H#�K��S6��v��2%W1��Tm��u<��L��\�����Њ�=p���V`:�*p���PV�~=���+���O������R���]�+��E�^��ͧ����
\> V�3h�ނ�n29▌b����>�:�;�m��W��/zg;1v������29T���{�9>p9��a�x�?@��dz% &]',qˤ����܅��Ã��P]��Y���С{�S%3�$���3~1�_z2_��}�NQp�~�R�9j;�Ĥ��Y��'��^�4ѓ���ya�>Y��[g;_�>	ޛ���3��>�<rM��)na�T��*��U���,�d�+S��/��j���'2�hrQ
%�~����[��g�@X X̕��nq'�)�T�2a�⮚K1�O��6��ؔ���C���# 42�Cw5[��PS�f/]���u���1POl����q������P�lCΠ���Ip����{M���~���-5�.W��
Gѵ5Y�B1�?d�ZJ�'?�c��h�	�uƓ	�n����$�G���O�XT�зK�g��Z�����71S;����Y�Ĭ/�_#
m���K+�jSch�7����������ڔ������Ŷ[�M����j�t���0���}�s`��ӄg�[��L�[|S\ys��֌����7ϕ�.y~I��!��p��E�qg�r?�́�?3^1A��Ѩ��j��r$������;+{���
��s񸔂�v��.�;,�oLLp��W�Uylz�����H���g�^��./�
�ӂ���uX�zM�s&�6��G��E�����l���ra�(R((�b���3ly�{�
�/��%�0#��9
̴�? �~�O�1��<��q�	��K����;�!�4���2�����:�������C:���ւ��������H�ʍ��*=��R)��2�Ġ|�- oSŴ��X+��g�=�=�Ь'eR����Vs����~��P���(;���'�}	+���v�n�)�K&��o捅��\L�)��wz��?�z%�KJG=�v�� ��A0#���cQ��]�A�"B7�=�}G��n�Dg�ͨ�z�¸��f����t�&F�d*�Pj�^������M�� ĕ���G���������@#Y,_�A~^����ض���Ѽ_�'siu�"�:��7<�`����8��f����˯��Kmra�*��>�6S�4���ۻt�c��a�z����Mq	P
�T���1��� {�T¦���-�c�@����ʼ�@P�U�uܮ�h�s��Dt�
�����xӏ��8��j��te��T�%�U�JZ�ɑ�Z�15�5EA�&�v�>֥w��8���Y	[��L��y��/��Fn�7���p�kT�퐲2�5.W�i�.�U��tH�},�v�>��aMf_�h�OG��9�pZ����4T���ɵ�ߟ�k�ѿ�V����E@��f�{Q#d���֫�j�4�Y�%�J5�Av�Ǹ��^�NV�7�U�.@�]���E�z��5��`ֱ�&懑G�!����}%�ݠ?�f��v��M��}� Qvn��VOƹ7�G�
��`�)�M#�,�~��q�<o�p�¯P�!'�	�	�g��:qLQ?{� ��{���^`��U(?ӛ7�J���T�wU������w"ECJp��猸Z@H��:F� ���dv�[	�L�ߨ4���j5~.��Pd��Px'i;%�n�3���_>"n��H������;���*Wu���d��3�9��؏��7�Dnk)c�RJ���4����R����/V�Z)��V�Ex��<K�N���7��$OD�M�Y$�Rtm�Uq�l�����Q�|��^���W�����TY�Ϛ�Gy��@����[�9'���RCea皋��A�8E�wIՀ�h� kl�w:ֲ���	���:2GC�Zr�H~�L���&ҧ�
��%�x�uQA�fX��J>ݔ�s%͎�_pU,.BR,D�h��;�̔Z��P��x��L�@=�7��.)+�5QN�ڇ��Գ��ǆ�5�L9��':8�� ��7���� �� ��V��m!:=�w��oB�L�i|�
�<�i��l�"�C�4&"�:v�U͟�	�JT���]h� X���u{��~����<_����:w��"W�o����o� V4@��rj;�q/ϕ{E���g\��i��@��
Fw<���+|���i>=��9����Ψ[~u
�����,Z��dc�P���^:9m�C(�qB�C�r��S��Z����<#2��ǮDP����.�AS�}��Y���y&�.ݴ*�~[t����v㔜C���f��:�����?��(��,=[`���
"�M,�f�k�#��j�D����a@��V4��
�!~�l���{��w	у�mr�Jo��N��ԧu���t��5]Jf�V��❇���	�v�s�H�x��W��-����ͯX���S�i�ؔ��[t�o�s��J���m��]���I��7b�]���_Jx�n}�kc����uc�nO���i
���O�ө)��̮
�aAx�u,�1i_��*��PXD
��߭����`�?p	R VOV���s^�z�N��c�:�����&�8�߮҉g>�:HKM�wZddQ`���v�5�Ӭ�02�05JݿL���h��+�8$Q�70�h_�ss�+ڭ�ݓNإ�Q\/N�̱8*��l������ʢ��޺�c\R<�����V���+ ^���X`p< �'�Tb]��eI� ��"�~Ae��sy7d��p��t�����n����2�ڿ��جHr���*H�כ9��{<� ��K����Ѻ8L�GB���V���%Lř���p��Y��kk��f�qDY��I5�̌XŢZ�2��u� ��w�ja���rw���F�9��lTu-�q����+0h1�t�����	L��}s��[���-�իq�o]�yWmT�J�w�0�k�cHg��d�`��W��)Wi�Ͷ�I�kVΎ8�72��b���,y� z��C��yr��15���9\J=�ò�i�+��v���}�+N�E0�,T㪏���ɐ5�] x���ʓ�gAlܷ��_�����e�~�#��J�WRIp|l���5�Pq�c��}����SPs�`LA�g�y�-�t?^d7v���:�z7�M��h�����f�ˠ<±��yF�q��������}�q�z��G*�f�ӥ�3EK�δ�k�#�4�cl�!Q�V�č�����*gQ�'ȕ%փ۫\��JH8���G�3��+ܼc���A�/ߺ��05���p��޼�ٴ�ﴑ"/[�ǡ�^:�eMi�������bb��}S+�[�x%�o�3��K���ɢ<�l|��F�܇�#s
�޾��{:le������c����Z�n�婮�lG߀S�ü���S ��n�s�������4%�@4�M��U2�@��.e�b���E)�Mudh���@q�i0��uPd�֞�5�EӐ���4k�&��&+����A|�uxI�Ş/����ک�x�~��=Y�cHX�<�aW��%��*�iG��f�&p��H���L6i�������a�X|'�C��/����(�i+��3�N����j��Ȅ����Z,Rc��i�oL7ZŖ���f��-}�D0��.׃Q��$���^kt\�JG��/�]�$dW�a" �=���{=�l�v����Z`��L�v�y��� ����H�� ����/nq�c�p�ˢ�Bu��TG6�K(mHJ^X�I����!�a9��`����Z��~��j_O(4z�ɶ�n+V����~����Z�a�^�2��S(�&-�����Yő��=̗4���+v�{����u�uw>�������W�����UL_�3ϛ�h��݈��2��&{�{�9�3ł?Cb�|7rQj!�@G��w�.q����z!�8�c�եfY�i���R�+8J�|�F*!�C$�EĴa=_��O6Nm�&�
 �o�Iu
��pzq�ߕ�s�u.��VQh����gf&A���n��5�na������{n!ĒiHNl�&r뫟��P���hc�*�Xb�R=��n��(��\;U^���	��Jb�µ��ӡ���Һ�p��)�Qbǎq��s�b"Sh�'3�x��y]��-��?���(R��+]��n��a�VF�+�".�O�����cZ�j��еW��r{�8syz%.S��[����^
���;��S����`�Ac
����l'/ek
���a,Wm����Mq먎^Y[~�nsZy�vqU���|�]�6jϷd����]��e2�:g-��Za�����\yEJS��d�,7*y���.�Ai��A�g�_	e��bc�e�x���c��'��]������ : ���W���/D�Ԑ��gkwz:Zd=y�P�#n���{���X"	���"��7EA_��z f�c�[�Ú	k�Ƌ�tpc+6:��"��{�$��Û�r�h�|6S8�%}�8�?V� \8����[3������gȉU:�KL|O�,;��3r�8G^��n<����C�Tw�&��5����og�;�3�ͷ�����/���"
����1��0��3��wSw�(�~c&d[�(<S��.Q�X(���}]$��`:sH\��.�ld%8N"Qq�ACz�j$0�	���a���\*S�h��n����%�a�+C�]<�)�Â��֌_c�gl:Wn��hD��B)��K@�A��{>�S�N񏋆IW�k��.ŻC����_3����/�]��4����x�����+�������ǽ��Ӱ���H�j���O��M?�3��'�o2jS׹�e>�EYc�F�'H̉��Sd�6���X��pEf`otTN�ɷI�������0n+;�!�H����{�E,_�QO���D,Ȫ�l$��$�B�����[y�($��2%�BR,
�#���D�k=�sT	���v)��Ϊ�;�m�P3P$�N�D���`a(�e�艹G�0�G�����]���$b�T)�K[�،|��d;F*��;��{@�h��t�rMq���TT!�c�������02�������\�⌷lӊF�;9J�IrW��=�26LУ��"�
�!���fK�V��j�k%�XCꀛ\�ٔe뷊�ҏ=1Q��S�A�< 0�w����tYOU�K��<Qk�g-M�����O��0V
���jc�%�s
`��[�%�O������J:e�H\��8�h��@�K��,�[���ҿվ�6����	�{0�SwT��@8��3E�� 2��:��+�sD7E�lg2e���"	�UP�`-�z.�u�&��bHL��L����D_g�"�p�N���tZ����n�%J����&��k8�K܎�	:��-�!��J?V�U��$�IU (�T3W��Ȉ:�6X׃���E�5܋h�@N`~7�.��\?{�j�0T�߁�Z��/{�����S�L���3�K��Z����imW����
I�8���Q8_��S��z�?�e���	������V5�.z����"o��崠���}�jE���\-e?�xh��x�9�O�߀ga�`�Azn�2tZ�͂�	K����>�<]66u�l��D�QX�90ۦ{����/���[�U�6�k�^~���
�$�ݐK��2�;�e(7��3���J)!y���fe�gh�3����W����$�C��ó�Jb.���T���=����B.B�;�2%�1��X�p�|��[� T���Ge���a�W3ڶ�q�@�u#^�%�,�7T��v�+d���#PZ����?�XϏMOx��<!�>�V�5�!���AyW��d�x�m�dB]` �g0�����A�ާ�M��c�T��I�KF�ZF������p
vY+J�Ԓ�O&�Be�"��A�O�
I�����V'׵�pU�V��jTӵM�a�����KW	!���e����Yf���@���=�� O���8v{ha9 Љ����iI&}a�B�+u��"=_���0�L�vN�|
Z�.��~?��S��Uʗ"�^,���Z�����i|L �U�$�'?ak�[�{������g?����D�á\Q�QU�0��!�z��g���u�֢�t��ܜ7Р��U���@��G^]��������H�X��H��3/��D mÜ���~�Qї���(�*�Yuڶ8Q�,��B����Q(*4�0A^� ���_֧mp���.��"B�<���c'���p� T��D�l��T ��N��T����5WwZ���S��fũ$9�M�6�J,��n��#�J^��KI�$�3_��*x�J�>���Hi�������A��r!(ٽ�9��M��=��|<�#�����$�ƞ�/�.�~ִ`sfY��a**	�ԙ���rP�5I��Ȭ�⢆�W�@��N�"��f�F�2�(/��x��h��׎�5o�%�Gq���aH4�(bO��osPK���d�:��4J=H(��~Ms��%�~RP��U�z�6k/��"�b���裕��o�%p�7�{��Z�?"��<oF�#O�Y�Q��`*	�4�!_D��v,��cp�4��˭�?c�k����;k0�ܺ����~u�v��}�AY���/@1�0~��8�h6n�@Ca��=hO�~����Y/`����m~W ���\Dx3���甠�q���s���zQ�0G�WWE�1Ћ5U��!FZ�10��h͑�aeJ�Y8�(5��3�@���_�>rm����U�K��qn˝��+ c����o�@��!D�x+l��Qm��ch����V`E*D\f�ߟ'�۠u�Ԭ��OEV�j�s��:6;�+����jѣ�g;��J��k������8q��jO�py!!����PX�F���J�ɪ���kU b��L��l,����pNr
�B�oE�T.��ޭl�z�R	�SU2�.c��a���k�214%~șw�zmm���ٖ���{��^�d*�>�R�;��?��֍���-�iOJ��.�iɿ*n� /VŠ�Bsн�14q��)Ȼ�E�V�;i�R��'��W3�j]�V�	/ذ%//v�{=Am:���7v�UzF|��[����ݼζ:$GRӷxރ�g��V��P�LU�i�(=]O;����*ԫ���!�\����	�>e�V�z�$V��� �����'q�-`߆cF�� Ʈm��`W��
%�6�z��6�A���LӇ��!�4]���|h@�6K�����/�`��ݵ����OG���O1����y`�;����1���$���Ú+�6��`B�r�d`�C���Ո,�<,��/q�\�LupZ�ck�uwN�-ctg��J�F�d3�Q�?v_��-IK;���:��_��XuV�A�
}�x�I��p�"Vr��Ѿ��k �Ȍ�b�&�%�H�)�65}�S���0t2X��f�i�T�D��'14�Y�Mu�^���Eji�[?�ع'�I`��UP��}/��E��d�} ��Ay����d��H͟��_k�ޔ��UE�K4k���@�& U�o�>�Y��(����S�LU�n�P����h�:�'�ġR`��x3t��A����x��64��j����R)�^��D;y����>*w-�]�g9@L��;p�4W�Tc�t�&Ƌ�/?�4k �(y��,�Ru�laÒl�zȜ�]I�Ppq�j�E��3qܱ������is	�d"���;0tՖ��땫��x1Еjj0@{��"�H!�=�H$$�_r{S�O`���b�8�-p(��d����gq D�.���<E�4*1�Vo����e��e������&>~ʍ�yid�W�<�`Guk]��Sv}�c�e�L]'02����;||ks�H�o�������[:2�+��0p�lG��s<w�w��]��A����m2��YJ����'wB!��i`�A*1fz樐��������|�E�n:`����)/o22����j�,�ą�5��S{f�{����\�p��{�\�n�`I�G΃@�ԛP����z�? 	��iF?�t�vT|���\�\L����c��e�B&�<����VYF�����z~�����$u5ڏ�>DuR���`����/�B���J��Ԋ�@��&�$���i��t�{"gr;x��P�?��v��|D��c���P�����e#���~f�r�;�qX����*L�{�]5�?����qz�Ʈ�y�x���9#\�!.d\��a�`�g���������ہy�H��F�u�Uv�r�5��\Z��S�
|��E���zo;Ј��%b8��1��Z���Q�_��y��1}hVx�:���a��5O65��>�ce�2�������1*��v'��������"�y��*b��� �)I���7b�����GK���Y����L�fj����i�&�ln�X�j_"���9teRC3��F�51��RG_K/�q�����5��  )x��>��1^�1��ʠGϫ�2:OEA/X:���|^���ĈMGy+D�×Al8�.l�))��/g����ݸ�$ྠ������	mSQX��7y�'��aԋ���Z�)?�5�u�vu�K��n�1G�_��Zi������}�%*+�%�,��z����U�Pj��~��g��a��}���δ��xw�`�s��(��kT}3��������ά֣c�N�K}�!����Y@MܞU(��q�F�5P�)V���pR	�=��H�&�#��j���� .��.:D�l$����[���ulC)!�:-��d���[�ݫ2�#�����҈����iT�A�V5e�/xQE�d�(7ʳ�-���^�Vy%_\@�8������=N;Bݦ�w���
Q����O(\gP+~�T�A�E`����<�3�C�I�띅��P���,���ࠏ��5���Ϳ�����u��.�J&[��e/Y)�1J:h)��R{�S*�oƒq{�,��1H�V�mn�=��l�F'�`!=�~�_#��ę��ȥU#4eYM>0�3�D��zB��M	��ykQ�?�]�p��b�����2r�γ�	Q#�����
���O�+�Vd��L�1�p�ѧ�� B��h���������{��P�AcԾj�\�3������oK�)$���*�h���7w�!�6Y.-oPy����z�*�ـ��;�g�ơ���r�<s5w�$fY̤�x2*�����W��T���l��Yk�@bN=ܻ�;�⤬>�y�ڋN�Φt�i�c��5Նc�N`iԤ�EcX��OW��/��&~���
�^�tkZ���?"�b�VVW7�_^åm�d+<�f-M�s��;ٖt�3�����H�g�~D�7��N�؅\��R	�A�;�+?�Œ�9����c��*۰b�z�L�O��b�}��G5��ˑ���\�}�#����juLe�Yg�/�@}/�j,�!�Y�I��'"��W��Y��fu1�x8���1.'S1��4d��z�`��ɜF�9���I���_�Q���8q~5��gXp3=���4�k���6��r����7=�(w����B��dc%VK�"-�HV�Q2z��<of��������F�hy�((ik��0g�M�P4tx��F�B���uڻ�A#p�x��nP��T�s������ �xrf��k8�8�m�#���8�I���L� C���O kyY�>7���?�XyB.�QX50g,ӽ( �m�&�����i�L��ؽ�s@��T�j��!)���ǈ#�2�=�� ��D���q$�1̥J����w]��K��'�7��T~���?��@8�d����&�\�+����m��]2	������⛑L|���ᶷTj�I���E��ث�����e�!�����ڀJ%
�1s�B|�������IP'������q
�c~M�tl�n���-������^����⢝H}��Ҍ���,���B�:�o�8xY��+o�-|��`���7 H��_������-{�/<�ք��/"�Br���[�⽜�1uӒW���{�%��p�0B��<,V���m����iDE(0��ܱ��A�8�6�g�]p��}�ߖ~O��������bXS��)���ĳ�W��S��}��q($��-��@�8oA)dœ��.+��b�sΆ8����3����#~(��Q��z�=R�bz�*�P�����absE(�y���E��l��z�y��M��Z�/�L<=�ri�� �8@���f-(*���WF��aX��{�0�����-
(QR�j�718
3N�2B��,+k#Y����l���BGr�$I��w*I,K�Ev(�؈d��NN䥵B/H
��	� " ��F%'���Z��������1P�iQ��st���/��F�P[1�!j�6�O�eq�Q��?ˎ_UAV��|�͇��|�>���c�v>* �BF�:��P��[l� �o����A��}��7�`�$�+F�4�mA*�x*'�}��Z(�K�=J�y����7�,I��a+�`�I��
�g�,�+}t���l���>.[y��e�����pI�;p ��&o����ɳ�v1n`�������F��(0f1z7=��w��r�|�f2�M�'��7�6V&�"�@�<��Dd�$�d���*3��#�X>�}n�V��RLN���x�xL]�Ƚ�GGs�J�M ��O��ﺊ|��2�����jcW�>��83��3 ��s��)���5�n�)�,�:ɠy)T���0��/|+:�<9=5���O;�ij
AƸ���2Z�ot��F��6
���8&���o4�����X#y6�N4]�*=�4��P</�ؤy98ޚ6���7σFVR7+�i�7����T��-76Ӵ��-R?�93�wo�*fo�#mݬ��a� \������8�
�_��j���vL/��ty�-(���ݦ�������/���X���~-�8\#�鑉\G�TI���J�-O.�����Am�D�d_T��P��5�M95J�-��ʱ+���*��S �vRBZ�Pq�B��!O�
����l�0��&��P]����'0��Pg�'vlT̉]h�±{��B�<���Cf���퉚gײ�̽w�.G��|�M�v�n5���^H|��g(!��S�:�A����s�f���1O�P��%�\��h84�И�8��+Ēm�H���=Q2�� ���-]_���|����ö8  ��h�IbqӮ5Qdsh
}�j%4a,l|�;�E��r�5N��exǞΑ������x���2�f*�J�Q�������1`Ke����J�ɴѤ,�Z���X6u���{�XB��$��h��q}%�1a��,���9�(�`ݡ@Y.9�I�̵�f ���,u���j+xSE�R*�nPh�O�.��Gw�9]ٛ��C+6��ꏪ���G�I��y���c�%�N�!Vs���$6�{_3�57�48 ��D����m���Bp�j�>P���'�o��kq�T�?*�,�d��ϩQ��_A��ՙj ȫ���
WO�������s|�r�U$?�ݽM�dږ�ڗ^��	��3�^_]�(��La9��� ؆��E�8	�L]}Q��T|�k8qR����VF�ݞ�X|ũ �h��%���[��G��jgð��%@�z��Ânh��
L��3��E)dSk���2
h�~�Z$@xa�T�,�	\Y
�5���Q����o�2Ϸ{���߂[�hDT j��-ՠI�Q-䖬�к����h��|Ԙ����'�1���� {%Cʟ�!�!���?P,�V���go. +&�y=\���4>H�����?�tM.�q��|�����d���&kԆD ������f�/�[�K�H�w����J���D\!�X�f���x������)�����"��5�K�(�u�$��މi�QZ&�M���"�B)4ٔ�(0*�x(]��0���J�^	]]/VJ��S��@�{a�w�~�Z��� ��b	߳���x���9��2K�� 8�����c��x���?�)f��9�j������2^������nۖ��BWo�w��HW&�������Q�[`��%�;���*�t�,���G8f����</	,O��Y����mFg>�D'
�I[��3�l�2��V�50d��0��"�Mw��<IN���3�Y%��M߾�4K�c��B�O������k���jD�&Q����f�%wd,Q>�� ɼ(c>��1-ȕ:���0%zx0�HTy�4\��[���<��٥�Ͽ�v0�P��m��ҟj��(՝����ϼ���x�s���O�������-a���c=51���æ�Kx����-K�h�W����rAm�@fDA3�����~i�,��|$�YCY���鶿/ޤ�bd�^~��� *�b����ο�x^a��ڸ�n�wn����>}V!]]@�i���]@�b1o�a���}LY�.�v�@������� ~���v(�fIiF��Dlsd� ~Ft�td�I�ć	R&u�3y��˳f�-�����l6��w{�Z�*8V�I(��  ��0�Y�r��F���FK[ܹ��*�ÍM��.7o�V��p3�����x ͼCWD�X6Ӿ��]�rer񈑯s��3b�G>�T���^��m�4���n���Vm�1���{���jK:�Z������I��V�W�|صhj���C/Nd��ht�#b-X��D��F��*���,�e|���&7O�P_;��.�'a�Aj�iɓ�0�]r�E!�kɛ���pz�*�<xꉟ�5͇iWC�a<o��ܠb2���@Ix����1�������1a�St�큍��JB�pȎ�$l���.�;ߠ��[�i��~��q����d�_Tb2)djm "��c�`N	x]�g��8c�t굗�ď���a��z�u"�0Uz���+O�Y�^�JY�F�HH���*���Op�(�3_|���+d�n��a=��?k�����x������
��d��O��7���K��푪��F&+��R� 5���9��c�����⳯ġB���2	��ͷs�:�L�Mq�Q���j�����>3^�D=�	O�+&%�b:j�/�����u���]]��� ���P����L����x���/@�۱!�Ϛ/��� �����%��+�:�ሰ1��9c� L��E�f ����%W�*^�� K�3HDhl���Mv�Q���B/�Zv  R��o�$�����Xwf�ԨԮE�3L����|��-h�Q�	��5�ؔ�dS�R���gך��/(�LI��<r��6)(7���5oS�9*r�M?@��Po`.�p�ROT"w��wGd�3��+Գ�p����pLU�R�|�{կ�	�>7DL����r�I�7o�QP�<���z�>����#y$L\9���ѵ?��s��G*H-��`��hc�G�c}	�U7cP�lC*��lWU�9FWV����	DB�qst }�<o�c5���J��Ӧ~��l�� _�o���ش�f����x�4��
:|�=�f��4lET}���J��8����1�x%��z�]C�����!<zy
��;	+a���IE\FN��4n�PEʿ�����p�y��Ɲ?���7n�����`J�^M����Ò���|�%Y$�ٚ����b_Ň7 �u�A��D)פ�Q��)�*Ċ+��B����5Q��-�Y�+]F��u&��K��ds<EX1^xշ�ѱ���Yz�&�e�^t�e<:CW	ۭvq�YDgw1�H�h�)_7gW����WW%����f�Y��U��՗���N��fs�n��f���k{���C3��d����at��iX,$'w=��G�J�v�=�y�����V�a��4��uN���Mỵ̄Uo��A�?���
�᷵�'��M���~z
N�sFs�3�w �:Qh[�}�-���ܤ���N��<��OR�L�^����d�<��RZ���㜏:b�8F��&dN��? �Y��z�;�' ��zX�oς�-\��jraFAmH64a�cG���Lʹ�S�bJػ��P�,��r�s�xqk�?ۀƵ�3�X��\w�^�T,��{Re��G<����Z�Rd��6T'��y�g+�yE�$f�'�jp;�׌�K����4qH�U���?��b�C�Y*m��I�Aܯ���e^���䅠��s�)���,}Ǡ�@�д�|��P�o$�sdD�R�9E��.	�
����(����6]nH��&W|�_6~��4^��4��#��,`9^o.;n��}s*��zylѵۀ ڧU��Q&@��W���
q��T�nNF�-��3�����1��Hת{��c���-wA�M�-��Fe�@t}��"��Х�_��y<G)#�� ��k"ג�UU�(O���W��]��b j�a�T`}fm=骛 R�1�C��nE��P�l�{�9u7���0r�2��G�*>��9��߮�J�ڼ)j)���BZ���Fp��� T|���A���"PE�x��7�߳p��#�{6`��/%�h�ꖜ�Sć����;�T�^�(d���En�ˊg���q�"�����eQC�؄��'k���Y�'L1(����h�AG�����V�^�n+.c���&h=-0D8�͍���D��10o3�l�R��ۤ���'�A��®X[>R5^��?+8K[O_�<r!BL���Y�븦��l2ͩ[:�*�D�W��V~ݨ7%l�zj�̓Y�՞##p�nkʰt���ۚ�D��T%���s��0N6s!�4�������-���p����tA�U���
Xʧ��� �t|�e��n|�OMf�;����~�l��w��U
4Pm?��Y�X0oU���K�Mz��$J΃�v��
��z�tX1:�*��.��d��[!X2��jY�q|�Q\�b�S�?'�2;q���%�ԓ���'���qDv����}oL=��A�`�e;uzf��2r2E�Á#-�� o���=])��Q"��2ݛ�K�<ө�����-y[Uf���a��1��H���$���gpRa�<�=b��]����y<#�j�ʑ��H��B��~	끈r����Բ���p��?�=��!��A�&���<&��kں%��z�Aa��5x2�p9�԰g�g��٬}ͣt-9=q��ыUiI�;)��S0��^��N�X�כ�f�15�~���i�{�O�{��3����mv��Q�S��@*���W�pH*2���q��#d��	n�xD�9������U��AD����\]?'�� �I�r���3��C��^M���'`!�c�Y�&bi�i��S����s��ց��d��K=��]�:�]�t���l��߁�c�3����iom��ӈ�Mq�Ղ��@���j�����Iz9f�V��Ĉ[f�&Ʋ�|�m� �8��ME �Ir��hn�m>�Q�l<�5<Wg�-ד�dd�c�����;������;�� ���	�o�]9B��P�W�ճ�k�煓9�0E��k�pU�+��^�L>�|��l6�ԃ�-��Sti6�q#y��imC-�4h5_�V�P8����E"f>�d������E*^�V�Y�G^햬��R~ʗг����x�5���C�d����7j�������j[�;	t^�r�W��q���e���tߝfr
3�{�;�ৼ:��Alg�ŷ�?�����Tj2{a {U~�֢z=O���	��k�T��Q|�7���e7x��?���C�z[Ll,�k ���D�36���,�.��n�X��nN�,xHoU`l�?b���\_W�)�<�|�)zJ�۲'*n����-�f�;��&��	�I#��j�����	��V��r�[0z�N�b{�9�D��4����FE�4�_�S�B��J�`��k�
�W��������a�k���;��:���H���;����7e�p�2�����$p�?�]5�0��{���|���
��C�sAyh�jG:�v�1J�Oc�lg��q��g���;�w�q\c����*(d�j�W8��4%��#�(&��2w�L�S���Y׫Ժ�^�� nRˀ�gg����}X��U/}��0j�t�"�����`�y)!�8;��f�#2-?���l+� ��A�שa:u�wW�r!e��������#	5J�v���ktf��yt��?��	<`6r�ಐ�0���W�o��z�����N����*Z��Ժ
>9�;To:��Ӓ�*� �&��`�Γ(�-5v4�'[��ן׼m<��a.7���go�f&�����H�uq��t���|6�OK������,܉��-�إwL�_�s�y;��@�����2��^�X)��8���F`,dE٦F�X	gu�K�3ȵ�̝�y˅~8�f��־I��;2vV��M>S#8#��V�������	0��r�
�]asb�r�ra��w���x��^����lo��ZZ�ދ?E+m�)�_���S0�����O"��iH��X���^fB�+�툗Yhk��W�?g��1��8���U�fA	��>̌���o(�� @H=��Ķ��8C�o��a�c%��ד(�)Y~/����m�������`�qJ�h:���`��f�0�(܊�)��D�8���X ڿ�&@Y�mt6����+v��ߟ'���#�
+�Y��ג
�r�c@�?`�̕�IL��#�eA��F�����px�(��i5]�I�n炈�X M�������[Q,e�����o�� �B�@���+�������'�\Ɣ��&hx0b��(^�5VW�Y7s/�r��iX�Oi�y�� >��X��Yb%r�Eh/�������K�C�w��'�0��u�x�b���ouon��*�����&�R!�c���;�0�������]�u�`R���@�,6V�XL��w=��M�n�K�h����
�c�]��&4놡�X�2��%LN���rd��1��,��#ߡ���č47��p��j6TID�v�d�HC��A�
����/ö���@����l��K)潳�#�8B�����Q���Ѵ�+	��-���'!����^��减���s�	���F�GJB�?�d��vևs�U�Bݣe�2�s:��v_�� �ap]�W��K7�O�"N�������|7 P�1hg�F�A��?�������u����h�c}��py��#�d�p�S�oJ��#A1���������q͘�?8?��g'�7�Q��lȟ^ن MFq�+�������x����n�@.fϿ�sOUg������W��؜��������M�a�)U��m���A2Dٳ�C�k�\��)�-�`جpD�������U�����{7����\���wɮ����L�oR�L���A�`����_x��� ��Td��I�5���Q{]��`�Zu�;�or����`u�6���7�HS�;�l��Xi�Ԝ+��$z��M�mz榵e�'�Gc+�����]e�
�G,�ur���&d"۩ж�q�"l�7�P���er�|E�a�!a����)t�h7�m���l���V͘a�^^5��n����m�ㅱ]졥Y�7��) �����H�V���;�yB��DT�
4e�Z����T�T�\<�مvw������1���#���㿌����r1��~�s� � ��,��B��h�[ų�x�O޾�p���1�a����~T1�[M������4*"�����Q���l'W�ggh�3�5%�"��E3�}�>��T��La�.e}��Y1��[\��� ��/���d��r�P�X���zQ�fe��#Ӫ��-ґI���:#���UB>�H˵l�z(W�؄\���0b��COB�`�]�&t�9ߡ@��X]�����@��p�%��2pU�Ra7ͥ��_� j���e�����^)��7�����";�����]w23�9|2�v���
���\��RR;���*j,]H/0Zl�u�oqU9�e@ k|8��Y�ވ�ח!	,��훾���Agn��|E�jt:�U(@Ǻ��j���t���'�YJ���]H�)��/�'^Fx�Z@�?�+��2ԇ��?���T�,Ez�=�̓�M�f�Ku~�|k���^�e(���#YE�W67�䰎�O������3i4:�`�*��=jmazV����u�u%V�/�2k@ޓ.��6a4|�fa�����A��E�8��f���#O.x|	e�];!���[\��(7���K�!E�ԋ�.��� xRcN����<�S3S{`o�Z����B��eKH�H`��ܙ��1�������];�L1�Ӊ������~�G�lr�R��E��*q]�V���܀�)�M�}굴N�?�}�lЭ���f�I^u^i���ñP9Xc��Z��r'�/��~�m��q��E~^��J�he�֤�l��&�K��f5�k�ș��D��hP���FQ��G�r �^���Z6��v��v�����"�ǀ���Җ�jS�`��X�u]�
�w�����z��T�Cd������9���ks0�/-�ᰩn�Z̈́�f�&Ԉ%kK��G���M���՟�����`=�M�&���r�&�(#� ��xRhA�_䑄?���f��!L&��a�Ɵ�#Q+z9����u���gڹ�ǇG�#����F�E<O}�s�<č{�s�m'�۝���J�I��A�̅Lm/?���P�:����~W�Y�~��B����Љ������:KQ���i6z���Eq��	��@���HF��TU����`�v��G9��ڸ�M�X��Ͳa2�(�:��#md��A��63j֓"zԳ��T�bMna��t*�6h�`Fơ��4��mޡ�GT��
	���;��R�7B�=���(�^y02�X��.
0j�;����α����C��l��8��q������]G������HT�����C6+>?t�Tut6���E
�f-�l�/% ���1�)�EkݲW��tv��,��X��c�o^��۵B���z�ٝ�忤��B�<���xk��`�
���<f'������#��Rϧ�c�ý?u6�d.Y��b�3�����lz|X�f}�*N��
<�+�)b��d�˔�����k���32�T�~0�ΟVD�J��1���\|��-�L�k	'�(�m��ѕd�W��h��AM��W%��h�C�����Y��=�h�ܜ��|�qH\VFٖ��w���eВ|E������l=T\�<�Q������l��=��{��î����d�A��`��vG/Y�N�%������B`Z�tK�CM5�F�L��ʂK��,\�kO�d�xe�6�Kj��v\æ�<0��o\��)�C�� �l�_�����q�w4�����Ji���w�
�ad��z~`���j��2xLb�����-wB}�kx�(�T�~Z��J�2�����adM����J��|���4z��>�3����ʔݳ#�м'1)Kr��$�ը35^a��� 8hhM�R�Rӻ����P|�2��N�q�j�m�mgR�}�Ez?4==�nݒ1ۇDE������m�A<浥Ʊ#��)J-��y�d�n�E�h/��)��:���!����KBsp�nͭH�N���5�m̘�%��\)���B3Uw���϶�-;R�ݣ�΃�;L�WzL+h<Ÿ��d4�j�+.8�"�@P���:�V"F�:z��]�����Z�]K�� ��T�wy#�����ɰX��>������v��L����Ց�v{�Hh����l6�CGx6�V"a�P���n��?���&
��{��1�ď ���-�U��rE�A ��m�@1>3L�kY��B0U��C���1�0* +I^���S�LU�{��<ǕҌ�Da���r�l������<d�VV?Ҽ��������(�콯�ç>�,<���R��>2��ӹ4<)2������(	)n�:)!�)��PKDp�u@���qQ�(�vV�B��в�:�m�<"%��v,	L�tE�;�U+2�A넧�^`��_Z��c^��
3���#\.�S�f ��&w�BZ�	�Ӓp�i�P0_�o��S��؈�A#��6,��9��4��L;�z=4q�FZ"�"/�y�>����/��J��������(������K��h!�\�3Γ�A"�(>$�Ա�0��EFR�������0=�(�u	�%0�-*�[�m�P�b��S�ˤp �k�T�u�A�=�9�H%l�/�ѽ�j��l�;W��ρ��:�	�7�6�T5IR�2)"L�ޢP�'!���/���;�AU������Xj� X_��	Lm��PEGv2.f6����{qğ��*|��Pj��[M���l}��7�Βxx�N!����UWޖ�i �����ε�e�� |��s���H��r���G����b�	>D=b//�����J����������\Db��R�Z��w�p�d���W�ew)E�L�_"�w��P��T�ԉ�Of��F���?J��4�օ2�������|NiG�oV����q7�o9�+o��9��N������ٳ�^N��v�?�	�57��L��r�Y:�� S��g�o{訾@C�y�6�����߷�{�O�8r�V��@��2[��ƳhU����_��h���%�.�g'.N(���$����u���l$iv��+ŵǑ/Qg�^��>v�FQU�Mi�ƣE\�P�;
k�|�x׵�Ǔ~��dN�!S�)��g��Z�*�G���;����Y��1��\�5
'4�s����Z��i�Փ}3���>t4�д��lJ@81+�t{�<^1י�'�٦��û6k���
���0F�Zٗ��h��/�.:"t�'E�ą`��_~p�ҕ�8$w�4j��|bi3k:-��>�lv:�A��3��OXDj~g�������n�&�����%V�Ks��/tHk�_^�6�Ov�Gz�TR��:�?>�=\MH�j��δ1�m��Nx[�k���(�[�� �Ze�{�>���5�q�W��i�	�9,\]��`��!P+%�Q�\ɽ���d��C�^+q�h�	�n�#��  ��`���+�ͥ�w��P��%���z(�׊��`��2�W	b4�"毪���#g�<ߥ[�'�>��K���Pڬ�1�AB��S=ͽj9%�R�e�4ӊS	(?E�̘������ʹ�ލ�M�J1��QS]���Y���c�ʦ�D��i��Ձ�j�f��������@3T]����|����J�9��]�`�x���e�MYc��rt�DkUn�A�A�`5H*��!a
���c1~��)�lp��'.��Pq 3���A��+dU��h~s����U�I0�0l�E�2Ubj�l��.(j�ZT��'�N�%�P��+��b�>Oi:s�5ƻb��%+I�_�����)�{�Y!�g���]/���EQe����2ߵ�d��c8!��f.$�����{��qBwI����6,B�v/��I�v��W՗�"2�}0��2����Vf���I�.b�4s:+2J;�����$�)�g�h���y���~"��+����4�Ϝ�{�O
U�WF�~����ˉ�W7������O.�hx�֐�I�w��W#�M�E���������>�=���/>�A�	����1Ǉ��bqZ�O��*���]v^B=Xf��Z��,J�u�#� �|����AJ�R����9�s@`���f`��w!#�.�r�>��ꈻ�mw�c�����|�;���3���\����J���FB-�`�}�Bg�Y�~�Ɍ��#�֤7�u��iض���D���m���Gu��K=�7@u������@��R�R
T4��wd��*�V�ׂ����c��G`9���ݜ1y�)-o���&�K�`]&�^���@���)O��P�5�t�%2֮Tq���'ǪA�����/<��邈�M���a\�s�Ē��� V��7ן �s��e����$�5��dۿݙG������Z����Q�$�6./ŕ(J5�矜�s*��2��
�2�>M�>��*뿉NqB�$>��;p��"ߓ�C(��7]X��̃$�P�f��{m��Y�ʎ]�}\g�N����8o�������w���`(�~��)��Y���z`�-��s ��7'�|i�¸AO$N�vQ�Z�36h������gs�,���@{˄(��q�N��˭�EƓ�`6׬���-���]kw�x}٘-�܁���.ιv�Y���t�:��cW!�<�����`�Sc�C�J���b�\��M3��5��d�?�%���x5\K��?�䂗+0���0.�>δ�,�9��/y��x�-�րe5�P�e����X��R
9��3�D�+�JS���GK/P
� ���s\)��.�S^� k|;��-�B���T���G4��>��R�,R�"5M�#u	��r��#�\�` ڕ�$�2"�X�P���ھ�^�s�,B��*�GA��������/+������%ĳ�FC�z^͒�������5i��� �P9)Ϯ`G
�krE��-��(g;ǾR���ٗ����F�T-)���f�U�U��>�n���|ʣ�z�+��I$+SI�J�ݨ�+rR3�A4�Ԅ1�������X�[:�dP����I�2����	�o�͠r�M1�Z�@G�2^�=O�,�y�ߐs9zq�(G\̔B�¶��Վ�qu��&��\�6�t��O�^Ll?+�Q�AE,�n6v����Ѣ l����eLe���4.Z^\��x�5��/;�]wsAR�I�00Ԅ�fBUX������'��C�9�Z8_� �k_��ë�\���Ģ8�f+�Λ�^�[���p�S�!e��L��c� %�X:��������EI��3�wk4�Vy�p��?6hH���u=p��u1�=㎬�~�O�����$,&e����9-�Lӊ�'��:��r� ���u�FV`5�*Bb�/�×S�z�����Z!�jWp���S����3����A�P�kA���Ƅ�C9j���)����?�`./�7vXPvZ��+O�xlA�r����Cz�� k��SF=��K�b5~���5��1m��%�;{�WjHe
��nD'��f����:NT�0���g�
J�=3F����7�ØR��~�Iw���?vx�F�����LZ��x�n�G�"��&lL#/;A�.���wL�ͯu��E�ŀIq�:|�^���z�� Tm��Oߒ�I�"���T���t4V�
e?�Ha��8�����L[ې���`
m�v�X�χ-�?���X�ٖMo��헲�����'��}����-��"���Y@iF�^��$����IraZ\X@1�iń��T�>��Q��d�W�	���^&9�*טּ�*9��"�vԭ��T+��c��p���jB
a+�H���|g�ɦ��|_��Ad�|�+�K�e���t�]�����Ȗ4�0@/V2I����X˂b��� 8��9;h���Y˓�p�A�?�3�w�o����@������jp���	�tS��Il4}��b�Lz���a�%���%�UC"84�JԶDAv��'N��䐁U�5"����v��BI���:h!s[{���!��Q�;������@��A �y�r�{p&އ�a�G1�;��~ږJk�7�XI�}���ܕ���D���6`��^OW�R�ʙ�0�����-J`jN�?$����_�{l$�Nyt*��*���; [�/%�\�*��0*��W�h�L�~�P�A�X���qkky2.˳2T��Kn`�����#�3;ڃ�޺��D�9��մ?�έ�Opm��;��?�TM�MT�î�ni�dR���=n�{θ������ �W��O	��cf%/7}f�����&d``ϗ�*l�����o`���C��X�\��r�d�Iڲ�W��[Z��f�$�@�����8I��b�0�XQ���?��`P�9D/�u��j��O&��HN�:�o�	��t��UY|PȤ��Ԃ��
r��EW�iaӓI�,,�!p= ���2��ѐ�*hõE_^���?�p���S�#D�1��`Ҳ�+��`MN�ķ�	�����m�&����>2��jЌCo�N7��Q�t6�_�E=P����kNs����U�xnľ���c�Z�!$]
�-1�k����?Ǭn��Q�M�hza�d�s�fiN�v��������}`�S4��D�>��`�	�@��vƷǘ�Ҩ�H�N����2ݥ�0"���VW��i��K��qhF���+��6l��H�A-O�./�YY��Dd�Ӂ�2W��g�䕤O���L��8�e�f�y�Kz�����Ɍ�w����@G觅����+ǽ��#[S��:r�Y��}��g@jz�"�:���5᧋���\,�a���5�l�)�ٮ�������'�.l8��)FL��j1�7���45�T}7U�3�2��:K�9��v�(�x}�Z�$:'��XI�I� S�b͂*���vW�gk�q�zB���aɽ6!��)t���=�+�a�~sR���Uc'��4s�I{1�;1�v��t��q�5*�TW�x���Be�t a9��K{�⇿�鰓�϶�"����!��D�����P�P��E��V�Od]uЊ8	�#��'����w6Ing>(3��Q�N�'��	UT���yD>��B-:L&��4�o��� W�c_�����/x"���m��ط ����ܟ��3i=A���X�O� 'p��	.@�'~+:W����h�NG �?P�z72=n(��N�V�fd��G$x�>ۚ�@�Y��6WإK��(b����&y�N�b'l�\�"��P�O}�X"���O9j�E����8���Lj�^+*ĵ���d�<��	6��U�G����OW��9�O$N��Y�.����-�~D�7a��	�������ȭ���#��o)��#.�9��>�}-��%G7�pNu'��C������-��z7���0�7�I95i���ibyP�٣,--��SR�Ӓ�U��*�Mo������d��%���|����^�*�z��B�ذ5�����6���3n��d�#�b�4κ؆بY�_�t��`�R�E&�w�w��ƺ|?�h[�ŬFO�Q=���2
�!�8%	�Ұ���>6|U���J|ۇqo.SЈ�[��1�F�rK,��V�އS{:����.��9��N�mFE���� ��o%��&�JV��$��	���wA����o��+�Ls��uߙ������-���yȮG�""�j	^��^���Z�yd�c�q�L'�`b�!Ex��|ಟ���KU̖.���~rt�T�ؤ^���.���q[]�ݤ�՗�{��uX<���D��j��*
�u޾������S.�3����|��s�V%tcx�����8���~����CK(��f��:ϡ�(4����x_�G�������͏(��[^�h�[��5A|��+��םs��U��Å�c���A��?�T�f�����2�#� �%%�<4����!쪟��z�Cȋ��)����gi�f��)�߄��
>���X��(e�JP��B�!��վ�7�Z���3�J��ϲD�����+��D �Su�DI�T9a��i��Lz*����Ǜ�N��z�"�@�'
�o�jY�p|��]�L˔�Qm�(k�����w��o�yP�F���(���9� %�LQ]$�`;���yY���I:Q���0�������m��c���G����^����'xY��pL2v��s�p�gJJ��蘞tL�N�D���N9E�K1&��Z���g�-A��ɜ�*.f��d�+�x�vK�,�
zh�+��#�i���:�E��7P�+Z
d���9�7�׊�n�J��G+C&y��Ɗ��5n�w�>�Kx�Ր|j�6K�,l����X�T���̋!��\9�$�F�1�$�F�����S*����k�Z�~�hO������Oj�&�30-<�C��,�A�0K��_Hӷ�3�7�Ո�j	�m�.f�t�Ȱ���ER����`�%�ؕ����P�5-z��;t��fa\C�s�1G
y�~\���0u�/ղ��7Eт��z�3�Nϖ
���w��n�����s����+�e�u���|��`���v�!EFN�|CR��IB���{�aG3E�-��<���p�z�Re�Y'��Vi����	�",�Ĳ�Ę��� @��κ�	$�B���5�Z(����/c�r���'f�V��	'��^iq��5ݠ��z�A������#�-��$�
���L������T���C�M��2N%ܔ�C�c�5���*\4������,���u��S�hO	d�{��n6����jv%0w����O�����M'e�''��n�b��ck�`!�Y�ûT�P���+%�����7��!�ӯN~�bѾr�jC��ߛP�Ss��
�$I��'ne�g�}��}Vq��]Lq1�v�e� F}�,�=��������q0�%	@f�W�^r�@t,70�@Q:����!U�à� �\�}�?Ϲ�j.��V�n����L*�)S_�L�>�*ތ(m�ku��>�T2#�7Z�=UB��P�1Q�U�������jLaΐ� "棯��f�ގ���S�E/b~�'�Yφ�@��X��*:Kl��tv^�y~��H){������A�z�.�a�d~�1U�҃
$k\���D��b���f�l����`������I��Iү"ؼء�4pHe�V�`�2�!�'�t�FOJ��E�X��̴��MD���X�+�?i�T��Wޜ#�OK[��Ր5�W"S��:�3/{����^�M����=��)��6��
K�:�Ŀ?�t�qv��8�ML�� ��f�vG�{�s�/�l^�M�=ISc�h�fpv1�I���6.F���#������v��'���9�_bceZv��\�h��S���!Ȯ��-��ʹx�J:vڗ-쵔�Ʒ7Y�9�c���e���KH�*��
��y̲0xݺ�a/ߕ��ZAt��L���]�!�.�`��ߦs4w�n�^|k)��0���]4�dt����m	�7����,�R=ְ�^�j]�î��+�|����98�c���I��<��JOjl��貀i7���z���R�i�ܝ�h#�f~�J��ܳ)���UH�	!;��DO�S�W��h���tp�Ł9�*��V��e{�y� j�g����:�M$�%}7F>P�;I��l��~�t�6`/�9�GO��9v�M��e���%�(\�e��ˍ�����'/��^�g?E�D�u��Aءo/5i+%��W�s��^>R6w
Ѽ�p��L3�� �WU�C�{��t-�X�[�Ӣg������2��.���j�A�8$��جW�'�߾\��؁�o�_�W�_����f����W,	�(1I�/���E8��DX���N<&��L�k�@r�����Y�))Q�	�I���I��m]��Z�:��ú�P%� ��U��/r���N��!��qZ�0��>��Z�G.��HC`�?��<�B��Z`��i�Q�?��I��⑩��!��a�+�ZѰi�{��#�)ef��*R��2��XB�>u��/41,��M��6o|�_�l[�Mj�V XR<��.������U�@Ֆ�[h�1�!��v�:�E#��k\�n�K���ͳ�@{�`aS+a�4N�r�� J������̸��ɸ6�#=�&�{av(��Y!M��ű$R�ڜ���5"V����Vs��E���#�v��`����1	�vv�Q5��R��P~9���N"ݘ�\Rx�:&�á���"�R�{K˅���Ux7��rV���db]��r�r�F��E`^'�j�om�1�wuu,��vt|Z�:sAR*-]2F{�(�����<RQ����O�R&��d�H@���y��`Pl�j\/�=�|?J��u���yG�	n�T������%�_<SlY�(���_����������`Zdt ��៩%�
!-M��������^�;�I�B|�HZ]U�~oY�	Ђ	x���͕�!�e�40&���V`��(�aϮ �qv��J�Z�&�b?�VPH�v���nj��ؠFDW!l�&������U�x�o"2�������D\8�7Ƃ��6�@��2��e�0��r
GQ��$����^c����F���$��I���\��K�%vv,��9w��fm�����]�j�d�����cg���������G�m�x�cWte�����A��!q,�Fv#�5���..���|ʐ2�3��w��:��p�0i�$�Ԣͱoe1��V;%`\+Z���	%�A��hԑ�J����9n>>U���R�B���%R(�UE>A�,�6C�K~6Ý0���7�Y�O���hs�-@����/ǰ��yM�rL��M ��ȁ<�`�o�	�o7ʸ�fQO���4?̤��?)�7Wz���;�Hd���..�l�#�K=�D������,�^o͕��Sl�jM�ŉQB�n���C�Y>K���!Zz�U�(*�r7�b`lw�I@Ca-QY�x�Ǘ�]Z:��۳""��U���;"���>�?�{������C1������~7
�^������!�'�P��D���)º����A�
Y�h�o�Ty
&yEg��No���:8��ؗ���u{� ��_O=f�t��}l%�e�6�i�	�AП������	0&�k�rN�BHB�����Q���3)Bx�\�9�=� �H��B
Y��
��(��Z">��X�$�[�VDF�S� 3I�����i�-	{�ih�1�Ð�� ?�1���-�(�ĺۤϺz+)¼Wi���b�Y������(����)�W<��X���y�!K�x!N�c/��������Ń��(�	ڻl��u��0 ��F�z���]��E����d��I����M(�ύ����V1��8C���0���YU���$%��t��L>�^A�^$�q��\��6�gӏ!�-lS*���.�D,`������	<����U�TA=uѐ�B�V��Ӹ�wDJ٨��/K:M��:h��hGZ�cu��	��l�KV�w=��I�:\��	�
{R�r}Gǘ���y���&��^U�vt�X����)C�kM�9�� Y���7Y���g���(�vT"��n�F�&
+;3n~H�n���O�,f�uX�'����1(g�y��bx�l �d�i���I�R�㷣%�c���K8OYSG
}����E�ryV��Ʒc��>�h��QK�xi���l�s�S5�d�U��8z����Y�"�%��X� '����'S���md۠]i<Z�ԵC����{�}!}�]�l_�v�j!��4�U���T�s��ӝ=:�,RㆭjɜF����#��Y.��x�J�T�=1n�۰0�)�C$�S�տY�_P���Bu������}�Ħ���֭h]�-�g(=���Ry�����!䄹����&CԜFFxϻs4�'���`�%y�b���-
#�@�K[��*�M���^>:�an��<�S�!4��p[[��s�ǜ�P���gQ�[�jǵ�?\W��1'ȩ���Z�@�}� ��9�՞�$�e�������p�x~I��v7$;��M�~��6���H"�J,}�&��.���X�`�쓽��&Je�#�f*d �ȅ?Y��N�eM�1�ȤIu�Iz���w�..kzH��=#7�i�1�nXv�� 셬^Sg�ȚԯHi����.u��jp�t�*���;2_��믎�`�8�x\��N�K�����;���^p�M���S9].�@3��F���?�͞��6��?C8�T��77�Q��2gD�o�n�5B�md�|����:�C�.k�Ț^�����:jJ7X��l�跘�4�1��ANs0����`ԫ����]�����ĨJ�׉�qDJ�p	Qr9�E_QJ�t�}L�m0.a��q�
=K
��Ŕ�ごu`~��xStW��{���Q��� {�9�j����:{t�%!}���L��â��.C;\IV ������8�d��'a����>b.Gp�XF��b^�䏧�``�~@L(_�dV� ���X�B�2�m��BP���N���`��3�O@#��������q�>�&���G`�æo.��A��53LUd!��Dwb�H�	pz���Γ[�~�mn�(w��e�G	�?���յk��.�q'�j�F���>Ӑ�؝�s�W�@Qt�E� �HQS���s���;ֵ��d�ɹ�U��|�t:�qu��Հ��Qt�����$`���=���=TU���-�O
U!�S�pJ�nSϋ	�ф�E�Bx¹��^�5��Y�s�BV\��.��F�c8��m� l<��R�m*X�� ��A��~�Z���/u����-u.J��{��g�9\����y;����~��_)�-�c�)�:��P>�t�[�C�k���VOk)�w�9В�	���]��po�;�����*gVq����Ұͦ��m�u� Cc����c�c����i�����
(�PW�΀/���j�r���>z����t���؜���y[G�1Vk~�mU�唐�Fa�́�%1o�fq�H�Rn>��]`L�+��v�f�7�&v��7Aڣ�)n1�Ϳl9�����{��f�h_�"���)��eS	�,	���V�L��O����)����^����Ԗ?�vB�/2͙72jm�����'T��Eg��|�3�z�/��(�2*5荒��1�x@�"���Z;,�/+�~��R��z\ ��Nvp��x�C�����k`6o_���M��O1n,M�s�,/s�mgk>�g�?u�3y*!�?>)y���4t@����+��9K���n��� ��6A8�$�1��E�1�$�YUh��s3u�C��N�k�&����J�Bx-�W�%M�S��.�i
h�� �O�z|:��+���x�b2��?䠱���� �	��
��F,(kU[��x_2zL{�T/�u7���<K�Ō�����%!��D�IX=����k�@V�������.��G{;H��n~�E'�yTI�=��"ї�c��r��D�f����xs��̡�dro� �I���^���������1�ݤ����w�!خ�ph�^m_7���P�:�#�h+��)D�������x�PG���ۊ-�6n��z�k:S��|5��Y&�vx�����Q�Έ���_/q�""F�t�t��!g���� k�[;�����j;(�J/@C��S<k�����j��s���*�O���5���\�S��BQv��
����1��*!p�G�Io�J"X4fs1I#�ĵ�ܗ��G� 5x2f0�1ɻK�/I�_�{Jsd"��8���wC�Rx�|_���R�qμsum���Q��ZL4�i���X�2��p��[H!υN*`(꾭�
+[ 8U��+2�bVա����M�-���c�q<-��Gt�/kF�O��L~���M����,�3��/B���qG�Te;�ǐL��wHj������XE�Ұ�Wd��K?<yH���!�@93�v�Q}^���U�,���ڢ����x�Y��d�D>���1Z~� a���*M�QA'�Nk����bD��ZL����
 ����#��:��S�7oXS���^��`��ċ�s���P�T-���I��>����5�4�Ӄ%��o@4�=�\�'��Z�����-t�F�[ӊ�އ>
랒V3��Y B��Q�0{B�6�8�j���B��_!Ō����ݞ�x9Ե �����E���z\����n�L8���Ȇ6��V�) =����qUYu�ő"t�u�0O��N�á��O�����*��O�I�J�p'�eݟN�4LXh��]ǜ8�.���������
����3
�1�ܧِ�5��D��7�u�h��a�e�F��d��8��&nŷש�\I�i�NH�ݔVv�ʇ��W8���ů	.�C�`>ܜ��5�ZX���z��I�X�G]��.��C&��U�Ƒ���͑����k�c�FU��<ݥ=�F���2��c�$g��:.�@�*���IzO�v��:����W"�p�bU)6m�(�D��������l�:�΁'c��ij�Yl�2����r�}���Q�Q�����ga;$�v~TL��uL��d.�^z?7<1~_3iᜉ}�+�c�湧���#s�zfr�0��:���l� ���aQ�=R�&j��cp� �܆�����!:8w�<��T���NH�?��3� ���(ڝpc�@[L."j�c��iČ
��V.�)	��ax��� +)T�$�����1{G���6^���o�,ha��-�"\)�%Ě�TN=ώg:��f��JP ]:AW�pQ���H��T7W&Mv��!��8�"��Qi�=)�:Y�q�Z��d�k�!;���/�(�G6�OcR��iN��K���:�8��3�X!!?='<,���_�+����-t�������zZ����R[��h�+��g��F|�FR����*}�V�s������d�^�+��f;2�c;��^���:4@��m1o��U�B��0ĭؕ�����*:r�m�*>��]|�_�9�Ihr�Ų��D��\MZ��C밂|��箼#Xع�X���0��\��9��S�GL���U  i���O���ݗ3)j�D/��QXJ��\"���*X�F{���+ ������T�m@�TJ���F�A��ռr�Ú�[�:�y��]UM���i��Kt��b�,��p�yD�vǊ��Do�E�����#�m*^0T�`��U�2��N�ɸ�o��UvA�Ï']��Z-
�O
 �ŭ���%��0N����&O����
Z�r���Xӳʴ�۞X�d�*]BF��s��y�w�4T6�A'v��C����]��ᛢ��ӭ���T��*/j-Z�3�~>�"�f�9zGPy5x�T���S��v�	V!����*��KL顂o�	���®,����.Y���
�����͸��%0o�ie�*���`�.G��D� �L�����qD�꫅y�$�m�gs���f�)%6.����k��͜�%��
�Z�XI<e5~�P�r�|B�D���j��Uj����&��/d)�xK3�c�2�(�`6�u-���uًy���jh+<8�s�	ty�=����a΄u-C�$��}P84��8���l�ۧ���P<�����D��LI���T#C��CG��u=(���r٧_�\=�|��`Q|\v@�ԇ����|�E�m�v�j�����伉� $ޛr&1zS��f����q��[o�R�R�I�f�b�Ţ�p� �|����.(�G!D*�v����R�ȭ!�����\ D r�iy���p[li�:��L�b)���7ִ4P2^����DR�I�c�����̻w� ?Je3�s[��f���#���VĔ{TI�J�^�ŗx����X�. �@p���Ԇ��\���.��f�����Q��;�,��Dj9<K2>�$������ni���e����27o���&k?Ӳ��wG��3W��K����,>l�&6菚�a1'�"�P���b��A%k��D�U���*G̯�smi�.��B*�ĥ���I�K�מ12��U����ߴ�Vɂ܅��'JWa�+IMl�w����o0p�y��Û��Hn�>6aF�L�Yq'��i(J�>"���}��2A��������Տ~��$���K�]�O��	d�7y��rU�t9�����r�����Vs�&����d�2�fD�&�,g�W�d�K�4��ʱ ɡ�Ҕ=E�{f���p��(���Rt��Z�Q�vm�T�#��2;#��0�9}�۳�o�x��z\��O�^��Ҝ:sU��ȕp,8�.��l5�J蘖��	A-h�h��Q%��WP�q�����&�#bG�/����xcSo��2}�#e�A�� >H8�s:��K��I�H6�k-N����j�B�[:"����7�N�r���,;�z�yКL��X;��Ov_Ue��q�=�HD��_T�E%�@�Wb"C��[�#}3�G_.)ee�
����:\a�S-��og:��#��!��v�������yM1�֝]e&�p��D����!�W~.�j� #}x���W�t��}n�X��ަ��wB�Ƹ��+\��}h�\O����/�),��~�M ���CV�\����,I�$tB�^���R�f[yJ(X�ۄ �����F����8���/��I./0�f�����Pm�K?��\�����1	F$X�G�����p��{.�|5e�Q����Ѩ*���-��VB�V���s>��r�
��l�+�mn�s�ݝǊ��K������������Gs�R��X�>5̻Q�F�hd���j�$a6?���#��DL���T(�ՁD�jɡ_��3�qA�c���><��D��"5��̓V;�{m�Ũw�������Z�����q⌮�0�k����3udK,?��RW�z�ؐ�PU�S��*�HVz~c���\��M��(gz:�{��n|���
���m��d��%�4��X��_ ��d���C��ЈM[�Y�;����@0�̓J�*�)����oK�B�����������a�W�]��b�j��j�R5j&�����0���}�U�4��,!\4h.�ī�ſ������hR��:G����|�vbf�L�������=^Uz��T@�7a�\��_�t� *���WK�m���*���1��VC�5Y���.O�p��n���=�A�p=]�.��������%Igm*�0��>�b'�u'��3��%/R�!^�S�C��Ԫ(�JM��5��~MZ� Y� �^�L���{�w��\��Ǧ̜&k�4��Sd9�|o*�X�������_$��`�0��`rr18�;#�qa)s��}�aq�l�z�ܻ�A���"�����[o�>�)*��I������6�N(��I���m��>����ۈ�,5�9mN�٧�m/s�����~L���;�/#�!� �=~�y�r���)N��g�q�f�G��&�,dZƹ�P�~�0��E�{>ߔ$����O�0��!N�ݹ�F_m�S
�K�G<%A~�R��ʅ~���� 7�(8�|�d|R�� !1���ݓ��?T����֡l����7�|���p����w�%]J��
< Q��[[FtoO| �2�O���J>��_u��8��!Zڅ[۵�j]���S<3��H�z油�7fb�GC��5��!dG���r�z��^=�b���ㄍ�ƌ�>"��q����/�}�q���u�Td�����ܴ�5�S�c.O0���Ql�+Aϡ�����}�N�.�I:�Ps�����o4�cm�8[8�@����n�����S�d]��2i�럕�41����\G٠'�Ɣ��/.�S~ws<�mEZ�w_�a�(�u�ǵ.�ӆ���C;�h3.��ŘYX)J<.���<?�%k��P.�w�w⛮?�=||j傄dB�����Q͎��O9��O��v���X�y��/�ZI�0h�7{��c.c!���ad�|���Yi"<q���Ɍ��)~�X����T�P�U�(a���K4i��$�[��j���;u[^sy$�#�'Kzk�A��mƐ��i�nnѤC-�`Ь]�_�%�RE�I$p�B��t�9-�Uz/����m�E�rOn�:�]n:}/	�G��8
��Vk쾲c#�m�K�H{�?j��=v�AN���o�n�`��y&ٜ��î��k��4/!2��S'v0���^p�Ҵ��e�7�������o(������_�l��1�E�֒0��a�~;����)$�R5�v⨦��kqNQX��r|��� nG+�|a�|]ǐ�����}s̼���%�:~�dn����=�V��7�Ȯ��Z����N�(�kC("�`(q I�qN��y,�{�%�9nP ৩�c�B3��h��CM\�T�j�x<x_��^z�Y���ޭ�E��kT����>c�C}��~GD�Jn�p���-�C�<L����<��-Ԛ����3F��C]R����bx����؀�꽲��DP��nפS�΢]jv���z��J�v�ؽ�D�Y�ӟf�MlL�8��U�+0�:,46%Fˠ�DT(DA�jۍҕ;����-���?P2��G�by��	rnI�~D�����Q��D/�����q4��Q�W����v���2�z��Q##�!������Qb���^�çP1q���oS� ���r;�������O0A �ak~��iDB�w���Q�x%<��{X�[�0�O.�O�*#�F��z�x�qx�����X�TqO�W�l�=�Qu[ԫI�Q���Sd�a�_MSl�e��d͔��_ '��X��ڦ+�wN����j��?����G��;��Vm;�i���X��(Ӯ ]�x#�"ֺ^�8�
cN@cy�Ve�v��{ο<G�:u-&��%���\�ۯٝ��G`4� ��ROD�Ko��{��2����s��IQ㚰�CI�s�;���?<�QhP��G�B��9�U�"=kǻ��TF �j�3@�� �L��-6����fC�KA N���3����'^Mbɬ�&�'_MVAx���� raD� ɵ�z5g��dVDD���-���Y���1�6GR��3�O^xX<������bS��,�Z��Wp�6Qw�]eԫ�F���N���]b��L��p���?��h���Y�Nv�6���Y���/��ZĿ���p����ć?���l0⦒BȑPZ=�~⧻?���砚��w(�n�z��G����GŝC�f���/Z�y��"��L	��'U,X�����[�h�Ⱦ,.�y�"d�	���i�`,����nи�0�@ˮp��"�u9KfLMg$�¼��t��ex�>�`6]��BSA} ���%��sQ�|��8��"PK�p��O�C.���q~ۼ�Z؉��ZDa>���<����.A���(ý���`߲�u͹B�i�0��š��v��,^zYD�����3"���\��2���)�~��`��<C������?�_6��(lƳ�����suf���6����: UY� �ݧ8�$�c����kh!%:e�V���k=CB��er�Ņ��<;���
��#��
9���
.�R�Uh�S���5B(�h�P]�*pgY�\���G�*���n�)dN6�O��L����rzP���'����}���C����k[�|[Q 3��E4q�MyCϽ��{?ۡ�خ�����o�A�&hw�&�j���/����F�`��E�V��J�>:��> �������J���\�%E7D-;����
Qv!��n�Ђ��e��(@w�U�;@b"v�� ��z��.��8�B��%�K�㖠�~��=r����I˯���X��8�G��7���f���2�0�uًWU���$���% �D���Qq�:i���ϟxd�,�/\4�J�xG�,y���P%Ӥ�ڑk\��1Uo��ML���gѠ�~�:����p�Y��/ɣ�[���:��+9Y48�����9�EkA-iXB�A�I@�Qb�H!���������ݻ�/�3"�P���)F�7Н��p�'���.{BE�W$m�慣S�m��)�Mn��]�y`q�;�\�_��Rf��zK���$�����
j g�vϥ�ޓ��<kŮy]�w�� I�9LN���H�Do1jR���(6Ù���ƞTV���;��}X� �d�D����N^�D0�`!�B��#>����ѥ~��[m��O�>zI�X��?�B>���=� ����cO��ɿ�S��!4��o䕺��w*~�i��v�)�N�'��a����_	K���g����|�HY��lms~�6,6<h�}r�[���%�Ml��H(>Fb�1jʬ�Z?hXC�_��z�U��d�*�e��j��T��줲�W���r����_eؕ�+����yqx���� ����b���
h-�,�'���j�����>Jl>�����b����r5��xa*C̱�V��$��"q�d.Vo��/��M&�
dS�����܀6�}B�$��Ci+H�\ a~eZ��3I��R�UJ��B�N�/5й��Sת���`:2��)f�H�@�aȯ1��#�K�
���a^�ŝt�"l��)"�W��i�ꙣ�s�C퓗^�U�!m�3Jv!x7`Cy���ڂ>��v3 /�Ԡ�5����J�[1�j���]s|�1�u���- fY* G=\رC¨���L73�d�����wL��E��H�|PaOU8Ó��>9�����F�k��|�L�4��J����D�,(��S���+�)W�U[TX'��N�O�̊I5�]s�G+�:�Y��ƪr�]���J��cRv��GCO�{Z���%c)���/��p���X���P]�Mo��8��0�m��6ˠ���湹����d$Q���-����iǿa���=��l���暥)��$�=��\�k� ���xL\�!���T�������h�΂.5� �����o�Yjyž,!��w��z4^�9t���7dv܎���ŋ���kuh�tS��5	A�6�;��,�sÐ�LNʬ`���h�Ϫ7<Š8\�~v������!�~Ҿ� �yp��JnU�げ���mԔ!��)��/�=v�+ui����_�P�}b�z.5��A$׽{M���z�SV��]\�G�(w�ts�{�œ���oF�y�5�¬�Z/���8��	���w��������6�"�`�<,���.��H�j�L-^S�v���[yr2�������mv�����oJ�!xU �>�������m��7@����U��	��Z>
Go\]���4��%�+D,й@J��:0�j��l~h������}/����Q1pg�[���|�,4S���5Oh�\�0
�zl{D����^'�S*�Bwƣ��y���S+[����c"_�6D�:m�&���*a��t��_�Yפ�}�57}vya�/��o�N������,�*�&��@��8� ��Ɋ[��Ku�����Y�B�ջ��^��[
6��u͌f�g������썖��I��E���&��X^�ؖ6n�@{�7]{�\���ݤ:P���..-�ل��b�_�\�Eꏔ`��h#����~��<��$�wRRk�"�Z"�W%	�FU����V�!��WA��>B;ˣz5��q�
���k��t��k�j�'΅E>�]�#����D�h��,����>���s��QP��1�0{������s'�W��Ƒy��v�#�9{	�L��8T��k)mF�tB'N�T���tT
&c��L4c���g:zS�?�/W�y_C�w���Hx���'��m�s\^�ê(/����A��]�p��D�>F�~%����]���ER��3�H87T��ߝ?Å@]z���Qk���	
��c%��A�D�<j}���b������4�F�k#��yvc�����䒻Gd�xąX��ś@/FH��������9����2A�\#{pw�[��,�_|\r�w#�_�ʻqD�@�=�����CZB�X�^��˫ћ]gV�׮t�4#�yTz��~�˅3u�7 ?)M0e�R�ܣ�|���~#��^�mci�ڸ�7r���G�8��e�7_�ďL�<	뿎(�O �yZ���f}z�c��v3��:K䔹��2�rң=���J�!��j�@5�B�>/n*;�����/��@y(D�)T�2;�B.����iӫ�4��+}Rkuc��q�N�8��.�(�f���w���kdv�}{)�l[���&9�x-f��L!1��CQ�#�^t������Jz�lH�jV^I_�	�CG|i'��9�ro�Cw��v�e�� ����`!���j�"Fk��N�]<��j��7��ẃG������0��s�s������0������S|�^�ʋ��Gug��P�����3d�s����^�È����m�}��]������Ed�ײ<;���� 5B�Q>݅bJ�B�%�DzQq�P�w�ǯ'B���:�!����1c�[�_/c�!��[]�Q����>���DX%��v����1��_�`y
���%�j����Α�p��&�5YU���T�����x�-`�Lc��H��q�Z��G�=Q�̃᪤��\T���PIc�r�i�X�3��]�����,�un*}L�}�`����K�����r�Q���-���G����u��Ii՘7�[��Oy��T7�����eB�f�o�HS�:5�S�wG^�ID�Yg�� B:H�GR\x�ǟFQ�����n�h]��rU �jp'a��{n�����~���#�:پ_�Ը�ʛ>&�a��T���xag�E#AЮ�!����~���Y���q��)�Iƣ^qүk�d�ѫ�ӳ�:��^�6ڵ��F+Lm �߹�8�=��;�lc�])�%Z�Yb!Q'\H�.�6R)������s�CU��<�^��\�w���Q|�;PO�lbˬ�&Y���$#8o귛W���#�z�)}��b̞t�e�=Y_�H F��W��޷��&X�N��P5:��s�xu����}攊.�
h�9y��]\��>��զ��xSPct��������~���v,!�E��":��ڛ��G���࣊�jʢ)5!�h�}YZ����#����uN{S�z��~{�5���䋮��mNi�782}M
�T�J���h�B�����[F����/Z[����'v�C}����-<��$r�u؇d��|8N䄤�b]^�h��l�+t�\=ݯ
3�|!��d���58<b����k�4W�
�nv`B���:ba�+�hu����H����O�a�G��l	 x^��m��*�.���:e-tTa0I-0���HIĸ�$����|$��2��5�č�n�Qp��5��Z��4tO��ɘ�?�h$䟲�T=?�d�� ԑKP�1��
���:8s����AG���	P�f3��J�F��(����$IPpD�VS=H�Ww�8�w���H3�
����H�<B�v���00��C�+�]
B�,8������Cq�D<��(F��DUyw�t�����|�t��f�~7�3*Dv�66��D�.x&�xS��w�B�B��f�B%hN�6����6	mm�߆����ؾ��|��x"5�b��z�k��*�����Y�@�	���R�]��d#	��ϠW��Ϸ��3Vn��Y����x[f$����z@�n��X�n�]OO�^�:n���<�l��j�Ĕ"	�E���<ZtH�M�B��˵�<�@�(OƷ�Z���0b;��� .Aq�4�.5}cцL|!ʹ �s*@K^[�!H�p��9>U(�
�h�h�s���lR�̻�.�i��˨̨9�8i �`/|=D&��ڥGq��~�+�~��̬�{���M0r�;�z����.k]&�g~�k8[�:]1K�`�	2Ü��QG�Z���J���{LM���L(���Al}�-J�V�WO���"�8�6�$'����bnk��!b�J5xi�s�J�uvS�A|2�W|v�����NHj�0��j�Nn��׼Gp��4�Y��T�B��}hp 8F39�[�eD��̦�� S��c���c�/���Li$�I���IH�!���wD�ڜP��.���k���i�qT>���W����3��^NO��*bp�޿��eT龔�/���Z��9����5��6����խ3
=��fx�"efZGsN�O5Ю%K-����F�/sKV��w���A&�:6k^A_3�=U8�O��;jS�잿��B�#�����b��� �l�9�~#l�D
x�`���n�@舾���WPY@!�IU]�PN��&|�,qԱƮO$�Oc�U��Ԅ�K_����y �0�����]]vX���"Ұ=�^�����Ǐ�XL�rrg�E/Б�n�Cp�|�v���W8�i�7�f12�ի�Ka ޝa���9��|�*���a8Q����RKOA�C�������_�l�A���^?�o5��YP-�J���ٲU�n��e��W���</uH��&O�'�J�W|��T$P�~����k��@[dg�b�.���ϝئ7~rʓO�$�=���]�����q�NZh�Vpi�Đ�����V�e�$F���w��.ȷ211T��X�)�狣��*����3K��=�+U8">����A�	� ��_��u��5-�<�?iΠHQ�"�J��`���=Q�%<kX?�wdL�s�b�M��I��㚃M�mB������1m�ָ�o�{���5���m!��q+����#�mԒ���b���)�6�]��'pֹ�?�O�5�z������p�R���<Y��`���B;ϯ~_�>�sGC3<����l=�&~9)%��`��ޓ���&���xU.�厶#iM���ڲ�n�E\����P��H��*ך����u��zF���K��f!�V@@{���;�x��U�%)���}��i�\��E,
�g�d�aޓN����d�?�{뮭l����3;m��N7��{^H�w`�D�(
SB�r�ס�Y�O*��R������.�"��Z��P-$��!m7��1�gj�azL�~��U�"���eX����.��!dx$L?�LH�&�J�x�r������qs�y{)oh�j����+TZ�狥A:M�Y�I��:��_(��`R7���g���#�Q<�A}����+<��˝���E^1<���8it��z�!%������ݲ�o�h}Vm��+o��0���ǟ����Q}�����}N-"����]x:��yv!b�Z�@O���AJwe�������|b2�2�O�k�a �r����8�;��T �� x M�6C�l�����VF�����,��/�N���ާ�`q�e�j���"�$!B �׋H6�)�����&�1>f��{��{E�K9-���.�%HJx*�T��U������"_r��en�,�����	�B�jvNBe�`��n'jé��	�s�8�%sC�Ӿ����<.t�s-�ۊq�N�IL��A���|������\�.��{u�1���w�R��/=��GHC_4P�����o辆���	C���l����er?3}ts��l(�+���w�˧����l��n�lV��B �(�b��X$ [d���z9>�b|EA{���O
R�I���P�\��	*JP	BO����~�^�N�.*��1�]A����J���u㑽"�$Xxߋ���^q�:�D��O5��J�ZoE^?��@w��Z����A:S}ka�]�ɓ'EDfn�d�/��o�W�?��\�f�ʏ��}ʩ/��:��Yj� E��QÇ����|�h��������m�|���}�gw��R\����jA����b����L�ܝ���W��E���wۯ3S�P6��^~�\#Lj��mM��O�0Y!;�����eT-��/��º���b<Ѓky�c�Y�=x��96Mʪ�NH�W���u ���5d����]��/{�ӆY-s��}Kn���ƍ��D��-i�W>���/�$gd��LYb��+���S]a��[F�D�0G��L�X�#�ʆK�Mg�ArI�ܗ�Y�p��������F�(�����
��h=�]���ߋ�~�����	�<;�Ul���N�\	� %�ݜ��޲�wG������P\Gi�|�[jP+���I�Ck�/u�Ofm���XzX�0�n ��(Τ�~٫�0q,�m�=pJ�.��.���n��^"���b���Z;���X�T4�*!k����Ԭ�<  b��?�k���5�����1O��n�4�S��]����Z����	�#��#�`��6i�����b�mQ{��;8*x*g��,�B����Xw9��Q��]t������'6q� D�ۇ�=��~ ����C���S
>���GIC7��v�^�������5ׁғ�������}q%`O�ߺ��/�V�l�ܶ�|��]p�)`P~M*ZǪY1!6v+���{��3�FH��a��L�kQ
+�Y�z��@�,�OL�+��r�,���d�˥f��4G�\�ޛ�!��k�0:w41�ae�X��=_8nC��q�^����T8|xy܏��O��e��)Ǥ��p�L�L�-+*\�H�D	,�Tf��k�5ك�e�I�d�;�ü� 3S/����Ύ�)��M��㤆�&�7W\�zS>�,�e
�*��`Wž����-mɭ�/@.����AA5CmA?�e�E�ypf���^E��K�����j���\mxeM��L�=�J�$�$��1$�ͩ�~�޿��w�uq%?@1##)��+0�T���6uI�m��P(�h�t���nX2�JW��y�2�x4oמ��S���Ҟ�#^����k3������$+N���cw!�"���QD�׹��>U�*s�p2��E\�.ɘ� ��Zs�[������Ȑ�A�(�L����"�q�� T/�m|����f�Ŋq
E�~_J(Ʃ���,�eٺ��"����g�Ե�/lD�c_��8�z�Oc�r;K3��~E�Tv��#�"�{�nm!je�l�w���y:����A���=�_
g9�#�hH���&���%��
��QR-!�#�6m�?�Q�D.gjD������ۅ��]�)!�Zߗ�5՛��n��g�ZS�a�3�֝<Et�O�����._�,�N�v��Ut���ü�bk/�ߵ�����%2Z��o5��g����C<�n�#�։��Ţ�X���&� z�����V ��uť�T��8���l����s��ɘe�z��8�:�Al+�܁f�j�5�@�9�l!s���r��C횑(g�?���@��_5<�����'a��aǧM���~�����8\[.b�R�T��t����K�t�i��i����΂X�E�8-+��q��g{E{���?.g(��Z�n�����5PC�y�
�� xld(-����r�t�u�YL�?"��er(Xrg*P����i;>%�v��D �΂��肁�s�h|�7�2|�j��9�wb��|���_<�:�*����5�'�.�|]l�Q�U;��U:s��d��Eh
=��	^L����j�|��*)Fn	�-�w��ѿ����z�y������)@f⣫x�G��Ki��H��
�5�{9]���w��ou��'�S�8�LeD�=pO��iIӁ��Hݡ�3��wR��f"���NڔNN0�q1X}���<�?�q$ך�檍�[����폧��ϐ�̯��dC?X�M��b�ԦP��+����b=�oC'� 8
��u��V�qȑ3oࠝ���d'�	�x�"��ː��s���"�#Qv_�vKS	v2@B�)�w���L���?�ˇ������^3Y���{�9�'���5Y�j�>��p:�+D��<�<VT��;�x�h~��-OB������tL$j
���2"�����t�<3�u����>�<���J�6�����[(��]&��� �mP[]�a�J8�9�D+s�<�ۨ�vʿ/��'�H�5�.CxME{lr����W���v�m�o@����q��� �NI.�o��a[�3��p+�-��C�F��tuA�^H�@84���v#  T�k�^a+q��&��l$;��3�I[�KbĴ��|R����|+'��MbGV�x"R�� $��{�!��KLF͛F��gٳ'��[���"��eX܀{#�¥`z6�2K]��D�ey|Xe�Ѓ��d���aW>u\�
<@�v����%�)j���'�G2��L1%�8VP_l$e�G<�^�;��ݭ�����l[t�R��0̾�Cy9��R� @���K���t�	�����Sj� �3o�743�s
,l�/����J�߮� ��TEE�W����<2dimS���W��J�
2|#v�`R�Gɧ�ۓۢ���~�x���YV_��3�-��v�����b��t�L�|��:�=�aZ@�0��"�����.��Z>1Y���W~�哚^��U����S�	h���q�xN�+C��i"*<������ǯ��ӦC�j4�8�2�ϸ:bN����b��2eCk�U^.0o�#URۚ�,z�S#�<����Y/$��kG�#e�pܼ�;^_�q�=�"��4HE��	T)*)�0�����Mޙlfo���;�P\o��Hɺж2]��]�R�I#�?�3��b8�!�Wdqu HKUA#x��o��Z�BoǺT��WQ	�e�B���%u����3������K�b�!��[��l��=I0B!`׌�p誽NIn��ޞ]]?Gy��]�KO8(���
?z�t����h.�R�=q|\�+�
Zg�m�/��-���5}��~+^m��1�S�áM��J���A��������bM�*�r��ͨ��g~a�SK>�l��;�� )�u�� �+�(�Y	����L ҁs[�(˹Uްv/�Q5�J;9�א�dU����~�B��OE���ᩞ�4�gl�Z�<��2�@�	�<�(m�Gf��/���Z$�5�6�'���&��Z��i��w�E���ׁ����Φ��"�'8Ƥh[�Y*b�w#��V|����"�3��5�G���G��i�T�&�۸�"���'�I��蔯|Qs��꧓�I���F��a��Y�X:���70�JB���Eo̴�Cg�.�U0���D����S��l�&?u\.�eֲv�.��J]"P�η��w���	��1�A�6^Ԣ�^Dh's/�N�N�4���_�~$�	��P���U�sո*�2�3(C�^�Dz��2%�� *t��f��=#Օ��ŕJ��Qܰ�Y3W�Pn�� � �t�4�l�buOE�nz�Ai\�/l8ܥ;�d�2���+���l���4��Y��*;�S��x� �Y[�©�ȼ�$c~Zv������9�=+���je�[Lh�JN$�C	�=�H���Pm���0.�1U�SW��	=�~t5rb�=�����m� �Ow�r~��>���=���CޓOA=q�G�l�KJ��!�d2��ySM*)u�F��h�$�&V�+'mpa7��@���l���ņ��IY���b�c�蚧�Q�<���BzRt�^����Y?Y�������\�ԙuT��ǬM���U�g��^�U��z�?���CVx��-Ǯ^��(��eLVU%�栙P)��$����rf�Mu ��퇓K���88%���� ��ȿc#�R��'���eU}�ï)d1:�#�G�B[�7,�Nж�r��UY��l�� ��ĵ����vQ���ƺ?�c2b?+�[;WK5��S�i������`�re'��y��zp<�Z��F�#�L�&01�l�[���Hܶ�Ɇ@�T����s����̆�t�� ���.y��]Q{P��G��/�q鉻��ġ�j��fj�W{�IDه�\@a��`^O��~J��F�&�@�B�a,OiȚ��p	���9uzzvv:�UO�a#4�9���3�nl��f	�V=�Ȧ���W�1�:�"]���z%�Za{	��Q_�iW���7�҃�	P��q7�����j��_��:��hczJ�B�=�6���_��^Ô�^���C1M�I�	����;�%����}Z�G��m�b?�.�����TO�(�>yR��c�i����R}�%���ˎ����úæ'K/����h{\9�0B7fQ�ed������M D���FRG]]��f���� n�m.����%�yл-᷽U��s`y�⓾:24/k�\>���
)��"��lZ�cm�bz�ӖOc���V�����'���1�S�.g���0�ߥMҟFr���9{�"u�Fv��Z��Y�����d<�j�HɃ&)�h7�2�r��A�Fݣk��	J�(��_6���4�[ھ���62:q����<�j}P�����Ynu_p�����9/��|(���Ƒ��O�	xT�y!���3�vh���U%g#������2G�/|y�I֌�$��l�6E�2�\���<����i�t��id�!��>�M~�[."駒�`�p�H^����l;�`e�lpQg'��5Vɟ�A�����Ol�Κ��ʏ�o�ӆ�.�<��J޽-i��煁%2'�Qn}�|^+Y�^���it����IH��ܫ��z��ug<8�ʶg��x�Μr��r^�8�>1�ֵ2ڃ�a�9G�����@��C?4t$�t臮sy��.��8r��z�V
7a��Mv�
�A�n��%C�K������!�73�;Q�r��a_{`9ۋ�����l���D������r�.�Le0���Uk����cB3�]*ʇ�\��\��� �s�$����²K�"�l�A��]߼G��<"uw��{Y�e���#�A�Yé/aK����2�}������0z�Y�W�zq�
����&���F�K�*�O�Qb�P5���. +�D��T=�b����*1b�vH�G�T�ϣ�)~��IT���X{t�#���iD�:m6+&�F��v1�qi-ۘ�����@c�h)Q�ɠ*CX[����T�)�?�Ǟۺ4�Id�NfJ D\��`�n93&� � (�>�MƯ�# :���$]S���g�E���!�6,J:n�r�׿��
uJ]s-�[ZH� ѯ�8`�������J�֫��m��8�Z�l|��d���1�M���LV~|{ ��!��פ�k#l��!��a:r:J��{R��L���n�rH���h��t��s���&(��w}"�$�1����6��2�c�E\���e��+M���0���|���ϥ�%ݐ���5��D�>"N��EP��G��Ǆv��W���w�m?2����s��q�;Pb�l�)��G�4}����h���+4�m�#S��[����%��y�)=F�Z���}���u�+��S�t�6���Ubf~IA1�m�bq��M��3�]�8�.���uL*�6tU;s��m(���k�2^@�#C��ͷ��4950R��er�+"|��9��@,�[��KH�MtF��O�&Xxd3�S�����<�L<HRLf�p+��u�y�d�xͦW�	U�C堚��E���C�'Y�>��>��V�V��o���������Xh+��W���ac�d �w H@[�QS(��rT<Ė�0��-(���w�(�[�A�~��M�m����d�y��ho��
[�Y&OSp3=�B���62����Ϧh���<��e=���ZC_V��je-L�r�o��a�F�e3t� "Mt&��U��N�PX���N�5;s��I �o�����i�S"k�h��VY^�.TΚ�*��I����]�&��kC�ݯ��"Bhm��t�#9�As"���a3�U����C��,���g��d��h�ȴ$�_��juY�W�眘�r��nw�i6��!��h�y)g�c�+�%�ǹRL�������Z�X��k�"���)�(�Pw!z5�e�<����R�t����R
=�LK������P����Ϣ�*�E�K�_���ut'�`|#�˔��z�����!`���mZS��V!.2����}��ϓ/��>3��uH����������D%B�)" _�S�h\, m���@ ��4-�F(�2C�.�����W����ԉt�,C	��/z!��-v���X�)fT��4������;1ǹ(^���)�j��\O �3D����15a	�m9��T� %�	3�kn.�Hv��u�"LxE]�*����z��Q$��	�r�dZ0l�F{Q�a��X�
qhr���V��������Kq�k����X���fu�¼ւHj�.K����k�&ķ>�)��.��3��BN�e�K���Q���f��m�͖6��r��r�1���4o�c���tĻ��[���� �vX2��ǖ�<x �@�M`+������q�q�L�=�Z^�a)`�4l�i�w(F����k��C�
�zoA�2�V,N�c�[���<���7���+�V �w�1���z��D�d>U�x%�q�f"s b��~���8�ɚ�Q��8�|@��i8o�2����^&%���}x�GnJ�ߔ����UV	gqc;�����N�~���ES7������[�z6���uJ�N!H�}�̇�e�:oЂ����[>��`&��qxG�	m�����X�2&l�Xx�v*�'�e�T�Vp�����2%E�T�2�g��i���!/L]��Fa�Q+���g���\���ܔ�GnI�w�Ļ�꼋;7�4"�辰II�_L<Js�g�����x�Pa��/r6��"���"���D��!j�E�rpl���i�Iϩ��J�e� ���s�5���m_=�UO%~���I�L��
c"��6>e2!y�E���C�d�lE�A�y��[8?�tܜH!jӛ?o�0LjY!$���ò�:\�eh�	�ל�����������`�?DY����<��Z"�f�a ���M?�Iy��8�`t0��与GߘwZ�����VbW�"�$4O`���ah���3��V���ԃ��}Q:8�L!R��x3�'�+�|�|g�g:�25#}��gi��9:z��o���������Ag.뫫������恏���p��L(�	T�͉�������]���s=6خT`�3	�o/"�}�8=i����� �l��,
UR:tӛq�Y;�#o�y�^M�!j���zAC����?�����ݧ�A�.�{H<�N�;j��� �%��U�8 ��Y�~�Ĭ�P�u���ro����\��0 y�tE�AF�ZX�U����Q�%�&�*5�9p��"�B���	��yџ�Xo�n2l��ɡ�2��F�FPy�_�>�m���տɏ�6�Э�nl9�~P�V����v3��w�@�'�s�\	�d���x�;_#S,J����Ť�R7L��#UFc�b��Y�D!Z�2�<͙Ww������͚��" PpU���r�-���#���h�R	��*�*,�G{0����� ���l��ZEv��Qc��wd��v#{(���<D?�$d��\D;�J�~H�R�n7k��h��2�*%�XAV�^׍R��Y�R7bE���7��B�6���\6�P?m�!��Q�KQk>2��?��3�a'Q��r΄��`�of.C�Đ��l���=-p�z�tT��-����2�0A*�d��Y��Y�ůW0�~��a�0Pߴ���zFQ�xyI��4�=�Њ ��&�r�&�zu�z��&ր~�PdxU`����t#h��sMț�� �BV;"[�?B��X�ʿ>a�d��VvP���|X^���B������/)�Z�j�V記�����S,�v����
�5c0�RX���7Pl�6�� q2��TeLo0�5~Q�J2�k�+�01�o �e����XD�i��K+�ů
�f.��k)r�բ��A�t|๋}��ug�0s��U):�o�00E4�e1u��i�P���3�Ψ˫��x��,�5�p|J�����6���ţ�hk[�?/�K����f�{Y��S$��pڊ�A�@{֯�,V����F̮1F��7p���I�av��Ȫ�쳎��� �)�gA rU�t[�on�DC��P����
�N��?����L�t7�����@��H�)R�����d�8x�8ĺ��Lㄗ*�¯n+����3?C�6-�R7�!�k�q��b��Ӽ���@<��%N��f���d\G�}~�L`���`��~p̊�f� u�&vB6�Q��s��U�Q�=�_4ԃ��~����I	���nU(Ԗ,�/Ɠ��x����;O~ɹM�$k*����c���'�W'+@`�CL�ߔE���W��Z{��-t��Q1�kJSE����ABA<qA��j�Z�m
������6�8��_����cn���6�B������&Ɵ�j���ڪ.dY�X��l`*7D����X0��^yW��[����Vfa51�O��p&`�=��Nz/󘴚�p�jZp �.��,)C[��I.��q=��W%/��:���h̦{��`�C���{K Pͣ 8��Oxl�'>��@83}_���a[7N��(C����[�	��(���L0M�g���>?H�3l�Vj�3��wXGx�p���xwf��'��,f�!��s�������Lnܣ�-Q��$�6u���㪫�xCY�R���aHFKc#c���S{�g~���PX�C�=;��1����Sz��zCw1W�d=�����*�sY�}e��ְմx�5�'��и`-Ef�h.U�_��v�R����|FwE%�ZXP-،�*L��E�`�fU|��AQ_��
-�-�d�~f��qԁS���|/˔������]j�B��2��������Ћ�C+��\��S0����r4_3�|���cЃ�o���>`Q����S�M��!Zc�H�2�n7Ki�҈v�RdR?�;���O�)�x|�^����x�-I�wYY8�=r̐��I�]�JH�k)D�^�Y�qv����E�3�Z���K2�]73s����|���l��讫�������P���z}X���w=��]��%�_O�Q7�nN�e�n��9}���T�C��4�X?�G7�Wr�E���%��rW�B����5x1��DmY�=�rT4�_vw.�}���^�!^>	~P�-S�ތ���s������~���>���ǋ������!'��n�"I�p�K�♞l"����J�l��*G�-Y�=�*�@�cq����O)��M}̥/d^�>��YH2��>$YA>��&���������&Q�>��/k�8�R�v�����]����d@���|������ N���jr����i�B��q��+b���{z�=#�p0.�+J���A�2�YX�_��Ex=u�w}	�/��y���2T���C�$�Z2e=�L
#�0�#�-���u�Yb�"��`c=������:��ŉC܅Y�p�.�g�B��c���:�T��&���}S��~h��*ᴇ�f��3tLO�^��;���a�U�ӂh��d�LD���]K�N�<��(���_�gQ;9���!�~��m�X��s��7斜9�j<L�j��.6��s\����v��O��>��w`�������)h]\u)G�Hpw��=�P
y���{�:�OO7���sx]�󣉀7���-���}��w�R����5Ȑ	��aq���]H���eTC��Gk����ĸ�Y�v�w�c��KS��}��)Rcҷʦ�߆���J���Q��Y��ۂ������T]&�G������졹>����	be1��,���Z�A�ݪ����a���
�����[��rd��96�eO���@�⣯��<�=��V7��0{�%$/��m3�<���{\A}�&���7�5���U,hXտ�HKv����n)+�W���Zl�)��߸��d9�N�jD�P�r��Z�e5���x��~U�����B���.����G~�Πx��׷���#
�^�|��Q���yU�(��0�VP�Ƌq2�*O����V��*]aX�]2:_�!XC�QL�œB?2zV�a5ȗO��ꝶ�+Z`���U��7��+��+����,������Ί^�g��0p5�=GUR�L�5k����̈tNB'"�$���8][���$��F�Ma��J�O�F��Х1.tG'�+�)fG'�ZLUS�V䍻�)�@��ʐ�ɜ<���5Dg��lD��]<��ã��B�Ч�r��8�t���"����lF�"pY��0ޘ�zq�!��sP�m��8��T�w��O��`UP\�t%˘��u�k�a<uStɽ�ϛh�;0��E�
{���i׵ɝ�C �w���+�P)�qM(�`Ʃ������=z�DFسN��"�
~����r����Y�`I�Cc��M���xk�|�1
�U��._*��4刵o�I5]�������)�M2� �ˮ���xE4_� ��0CRQ�%�	Έ�\<z;�Me�^����ۣ�P�mJ\n��SC��y��	�J�Z�i�(7k�/�������Gm�7��\%��b�������5�,xWXH��U�����s������A�W����
`��$1�� ���aC[j�� ��?�F9�`Ħ�ro���3�-�@-��#y_+>�}��xG�%��J�E�����������ï�|a�h�h)����;�}%��Ng�F�����x��;�Mb�Я�~�ev-,����V��l��!K�֔"0�n�P�������z󹱜��#�z�f_;���ܵ�ژv-M5O����Ѷ&ݺ�[�>ޓ�Yˉc����t[y��Y˔�)smm$�J�[�e�Ѹ�&z�*�Jڶ��ԛD�<�f�z��T;U',#�8&M3��yyQ2��,��!#��N�(��S��XJ��˫���E;��C\i�a�$r���њ�FVX)���M^�>���i^u�w3�p-8���Z��?J��Pf��*��{���~8M��R�̣t����q�L�*�^;���Kdx�
ż��ߌmP�1��1���nXB���g�Zm �S�%��?� ,{�4D#�#� �q9l���9-ዖ�9����y�ҦH�E�kC�6XUx�Ϩ��؏���M�N�xG�6F���[�U�DV��}7��F��ʍ4��%��!�C9���D.,K!-�8��s{��`)
/Kȋ���Bj�e`I�>�8� �`�4j���*��].�nM$?z��.P���������V�1�]Tj(<�����l!�ϳl��S����
�f%:/��Vr|���K���Է�n�$�V#o�֔��cnt�R��)�v�Qϝn��{$m�v%�>�lXѬ/1����V1����e�D��3]Vy��A[��h�q0��x.�?m���0�3���6T���7�ů\��º�o��˦v�t@��b=aA�����	�;Z.�!���)�Ꝏ��,a}����U/��xhW��x��X;8|$m��\˧�/L5��i^_�խy	�%C@��7�,M��;��5kb�w/d�s�8p-y���j�K���p?��sW\�%�s�8�eg�%%����� ܴ)���		�j[O�=s�6g˕Y�s1�<��c��,<������@�p��-�5�"�3!O�*h�<p/s�9+����z��<ߡJ�"
�S�h3,d��{���������e���l��.ͽ��a�����ĞT1?Jq��ЪJ� �T$ �KC�W�.�_KBb� ��T^�x�Є�\��놹��	�-�m=M9/�%����5*[n�(Td��/s04Y1[_q��o̚�<!8C�ak�k�1�ӈr^B�&�Q�\����?1K���\־r�<�D�9�#3�m������Թh�{��W|�r-v�91g��O�b�~�ܺ��v�(�d�4ؘ�����T��H��րvN;l�^���O^~��-��U�q�0O(f{�B~��FO((lw\���@z/���Rk���N��� �k��o�>  (�"�_���yV�c���m�O��mcڏ����#��ۭ��^:�ս�(��O��$ԣ(���by�gQ���kxM���e]�%|#1M%�	'V4�-x�m�{�����V�� QB�.�4`���wGI�K5|�����D�J�����A�J)���<R���Ƞ��U��$=�y*�Y�K=:�7Hs�Cn��Or�
�˘UR�q�J]yQ	��Mpq�W������S�V��ΡϾ����Oh��&�C��dG�,��oK1�?�
T;�"7�c)��~^����2�q�H���2:��:��>		F�&ͦ޺�Z�4��1ğ��'c��m���j�����C  ��4�qd)Xb�`nT������]��m/�=�pe�HO��)�+$Y�c������;�nS�CI?�&N�,��k�d"PɁ@e�V.w���!8i��v�� fu�LRcI���'|�P%΀ �&���&�aHgl��&������?�y����>1w�P0����`f��Kg''��)*�5���1%��LԷ�&2�����}\MT!����ǻ�d�GD����Y�9<�O��1�̾���PމX��D���OX��1c����Ϗ��Fwp�TK�Ȱ����'Xi�*s�G���^��R	�	�#M��%~��!%#Ѯ����6	���Q7�s����-dQKV �m�\�I�r���m�?Rn����+�	��F}�&f�/˘��ԕG|@�5��}4�ɜ�����U�`�z=G��1�e��J����	q���q��H1&�$��>�Ҿ�[�[&;)�"U���O���_���o�5{l<�l�;�&;RԪi�$�����X{��cy}R=����2�n>�R���0_�2q�����m�`��$@a敡����:��z�����J�]�F;P���CϑV(�en�1�Ld"P���V85���6��܋�w=7/�x 弤9���U�#c��nAn��SBEH�]���Gs9�x����<#g���XaF�!�*��cZ�W���!	{~�<m����y�3ɑ�����d�\���V)s��!��߮�=���0h�RX�I��b3ϴ��\[�7���EO��ے���?;WI!���	o56��>g,\��-Za���6�	С��}��kLh�'��k���nn����̈��b�)�Q���ˀ@P��aF����l;����L>����n$v�Q���!R�KQxr?^��9g��d�:����_��ׂ��8��A��!�\�Dʚ�^t]�*���H�� �RC�'ec��!���D3�&v���k�����8N�||�nfg�9;�Pt{��$�U;�I?i���&�n�S!Kc!��������m�8�*G�߆N�J��{x��)4Vv���&m㧵�sʾ7�X�n�����A9qݨ�o��-�C���<&����; ��l�v�����b�����)�Ӧ��q�@>��@$�)9����6f�k=�h�+(���2�����N�ăl�v瑆�mَ�PO��l��]�e������ʨx��7p��'G6<[�Qg�]0>��%�KyU�)�b��L�8�U�,˺�#fȵ�?�.�����j۲�˝Gv.T*�F.�4�z���,>�˛�v�P���6X2_a�� ��.��7*]oy��"y�(�9��� T��ᦥ!��s��$)��S���W�.-G��;q�--�'�gǀyX��?������?�d�Gp���:��ujD�>��m�5�LI�zG�AX���I�D�L�E�hCF=4�K�Ş~Ӷ�G�xC�x�Ǯ������`e���ֹ��M���&p�x`��L��ג�}�+�.4�GL�}�}�9ǉc�P�-��1|��lV������A���.D/@r�r��f�7ʹ������G�>�m@�Lb5��UX�$��Eܘ��E)��N�6�A�f �R���$�~��"[���:K>�8bj�M�eĻ�/cw$6SDU�у����b���=�e���9�5���d<�Mr�JrRfA����7TDs�ԀqU�Qx�F�ZB_�]#���-�����2<n\}��2�q�0~�S���>�������((�4��RVm�7�T\��\rS���tMJ�7f)W�@6�^���݊%�ꆼ+|g[b~��ݕ��."��	ܲ�"(4�p/�[����xl��3�3��"y�rhgCﺛ��EJ�k�ʷ��EԿ��Y8,�uЦl^X$ȉ��qЍ*.��2G4�uTpQh������a���T�RU|��Z$����|Lh���q̤F�ihbdr �]�A�#��w����ǯ�D$P�3j?3a�R+��Yo������?���=@D���B���"G�1�s�NփN�rx�������������>XsG��q'SG^���-��7Bf��F7�M���O)���8�8Vy�۟r񘛻�]>���N����8��-e��&C��+��7|ĲU��c�&�g�P���D{�����2I�!{=.�����p�E�y�WPF%Idg+)V� ҇�� �C�b#�7Z�� hbkqݥŰ��k�l�~S�)�s�L�Ϊ��}Y(�r�{]� �q@���j�4�n��v8R�
x�?�T<�^˹��X/�S���/�萿Xލ��3�˵�v�f�T��	�������`؛a��K9��$��o�u�mG�ɭ��׃1�����W7�� Q�Xq8�+C!���j�k�<�2S�,��q�2n��E�]K��Sl1�z�pŰ_���:�Q9B���N�����	��E:�0�v�_�Ӝ�6��� i7l�C�j`C+8h-�]0Lz��9��R�,���6/�����l�xvH-��L��*�-g�A0�EYQ�>��x����!"�J%� ��a�D5uzX�������Cv��ŕr2��yo�Q��,�		Gb��3^P��z��0��<��( ����(`8+t!>K�Η.ͨݍC�#E�۩�9��a�˶��Z���D��Iכև�9��?���j%Gc��Q,ѳ� ���V<�u$4��eʃ�xAb<���4��,�i��j��V��Mܹ:%0V�BQ�l�e�ф�؊��f�&y�@M�Yq+��[�*��!h�p�H 7i:���+�ґ���	B�Jo������(�����8���U�o)�e-g`CS���'��_���6񆂘e�����.�'����ds�5���<�N�@�$:��,`��){1�ǉ���J<S@��X�V�K�o�=�ry2�'��)֙�{. ><e��/n�8�����u|
���k���c�U?ru0{e����I}q*����K;I��^<�LD(��)a2���H��w���9�|���@ Wq�&�s�e����<���A���Y�z�7��c��7|}��h��]A�Q�Kֈ�躚�/kPb�&��I�0���O��
)��S���l�=ҁw�$�"� ��
�����I�_��;ʒ�9��(HHH�m���b��:�7��i�k_������p�zTt��$��t�����j!-�
K���(q.p�^�D҃��i :]*���ʐޥ�s~��n����`�ʬE[������|��k���޲�U;O���]�-\;�F��b`yZ�1�4)5r�h���(k�o�1�_�us@�iA���V�d�\УwU��Q��5e&q����^�|�%<��̺�Uo设�m��u�\�!�2��<�h칸�����v��q���D�!�{ ­�K�N�,��$c'���M�9Ma�1��ݝ��/�Ă ~�7)���Ļ!&j�6�N�Tu�9�lMv>&6��Z\@�yZ�eT�c�>c:U���Y�% ��-SZy��[	�f�;��R�R쨝-3���\3�e�°q�u`�-ݦ��������`L�3��]�������OV<V�t	�������+��鋺2~N D�W�֒-�
�Tc�1���}�1ԃ�z��k��Du���������i��Y�����.��N	�`�;t���F����+W�y��A���j|w�>�"�PO�3otW��@�1����E.&����5�j,��s~ ��jad⯖��|������2��8^ăk�@-�^!e�?��:xa��1\��t�T�����&�DFq��m��S..��vå��"A�H�w�q$J�a<�K���+<��|���el�P֗o��ۉ�ԸN��e;��ԇXf{,��/c��:/嚈ҽ&���x�>1A)���,�Ȅȓ(�(����&|/H��^T�ǫ���CJ�Gǋ�h��j��R�jI턓w��A�
�@Y*�[b�����5 �^�u�1�S�%�#㏪����"x��OQ㱾���U#�	�41K,�(I.l��^�~���W��ՋϼAC�M��K� �)������e+Ϣ�r�Ʒx\�¶���F=E���&8�zl�'ᮦ	G�9����Zb��^��?>��I���%F�o^ZN/�B��.�z���Qa`5/kX+�İ�;����K�g TgA��ԉE�C��c1��ΐw�FX���o��qm�����s�'Q2�2�&Ԭ��M�
���
�	0�nl��0^���=���w��$r+���Mp-cE0{T���8����ڢ���%91[VC�7d�Ơ��#�0	�m&�oan�I�B��1��N;S|5�H����Jm��9�WpB������r���V0Jq�L:�dU��ݭ�R��6��r?^�?��3t|B�*���dt�\��oV==) �-l
���T�[kW�R������|g�@!Ь'���P�U�Q��$��b���v����j���@����������洺��'�����2��|�$*5n���e�ƺ��b��s��6�Z{(s�|���{�+z�&d�����0-۶GFޖ���?~�e4��H�l��`��*���iJ&t+�WYI�w�>�J�=�\���
	���,��	KUE0c�D�����s�)Ec�85K��[��o%l3��^y7Ŭ=�������X,ap��>�7Hz!���5���ߤ|F;~k�:�!�����k�۔L���sHik��蚕"��������O��%�@��q�PT�p��CH��b�?g5jEIV��'�>[��8ơ\�^͏�j�0���|}�H����F�7[�g��7*=��yV$EG��*��/PZ��V�:�'n�L�|�^95��w�P/�A�^�1���@�,��!O���6���7�5i�f�0b�jq���s&�}Ֆ_Jߪ/�WU�ML�.QPJ{�]��q�f���ط�����E�M)|/y�4�'7̙��c��i��*�KʫC��?R�yuL�I�3�߰��@���}�p����US�(��
K��*�I������'�	䨗:�c֐9H7��~OIg�z�U!8-K�.u@8��^@5c�-T���w�Fo3�.�f�q�L9���U����&>�o�Kfi2=H����Ϊ^�	9�vg��HQ�u��?c�!ý��u��_=tW^�$�p6�;Õ)�^~[B ���s&秤�K��Vqt�fB�1�M���L��aΐ��ļy�ģ���K��������z�F��Y`-�����H�of�U�>%�u�<ƴ�~���C?�!�����MWh?5b���A���XhGȘ��C�����@��n}�J���U's�`Ӝ��wHC�CV��D�N^l>��_��ɜ�kA�tV����H���H&��.�e`���e�i��uD� 4J�BHxM�k�D�U������rkbhl��� 7�a�8�� mC��>���Λ�v���R�����%锤;�ì�b�"k�#���gW �`62Y�l��Si�arw,Y��]T���2:������.v��H���+Y+	��܉�>A�Kl����j.�,S�^�A?$C?��pR���t�k�Y�iU��70�Tm,���bH�;��!~�.�e4&���U��[1�Z�j[�J&L�r�g�z��u���C���D��:�>�#:1Eˍ�ɽG���8�e.�/j������¼`@7���!���V˪�P���C%<(�M�}�N\<A��7������n� LO!��)�?F�:q<IvDA3��g]�w� v��ᰛ.��sU;��enӤ�|�=�RǇA����/�]�9۽uZ[�	�����ƕ���c$�Z��/3�=�8�
a%�u�L��/)��`���\���J/ɂ4 �������?�L��@��݀���5ݽ�����"@9>ދ	�EE����Qx����[��0�+%�����Ϻh+
�#���`��jK�3�6�þKw �H��$�<�nn�kK&�hJ�A���O�[sZ>�tv8�y�U�x����Q����hM�7��Ķ�6�ڂ5fL�L�, 6�s���)�v���`z�����S�ě�J�wb�3��4�{\^�#h�4������Z;0���d�k�rJbw�-��(d�J��Q}	��=�6�om�}H�'��t�:�g3�0�U
� �w��/��p�C�ӛ�pu�^YOZ��:�A�I1�i@fkcխ�A�r,�!�=�l�F�)���x/g��G9�`�\��zm�ٜ���I��=�-�fsc��b�- �3y�(FpK��ԗ(h;5@^J༨�A��]PS�m�pR���7;}8F��%�����Q ԎOm��}1����B��� H�1{��a=�b�N��VB=nѸR��Z�i�H���_�`� �K��Z���8�����z�L�	�{�Ҽ� X�y�ҿ;cW����w�Z-�fiD�]U�aE=����0J���;!Bm;'��4��D6��/#���}O�����f�Ŏ���H�v�5;�F�S�s���[�"f��͙`�]|��V؟-Mv���]<3�{=C~�>�IY}�T��}�Ks�����ŷ	�@�{�.��xJ�=um�2�ý�axY�?`!�U��Y�~���X�[��[�9�+�ì�w��k�~,�Ӈ����"7�zEq�m{U���y�&���K^��b�����:*�]�u��ɝ>��5�	�y ��39�[�L�,\�h��㫻:��݅_����#!(Y|g��k�13ؐK"3�'���� � b��N�W���Y¡�S��[�M�̩>�`z���W;X?���W|��O�9�R�௼�0�]��"�����V�x�xԹ=��Ѵ��_��I��5�u5�~X�����z��df`�@��3:�.^�*-�'f00s�y����d%e�$XvH�$�g͔��8&G��4�blr��A�R��KS�V֜� z)� �Z�{�r�nt;�E���i�=��R�Rx!�;��s�o�yIO��(�=I �=�L���*�r��? ����"��)`y�e��Ƭ�AL���|� :��1�f�yA׿�N�� �MKNZ՛��h&�$��)�S;@{"��2���9}+fs>�$4�ã:�=��$\��H�����ڍ�]�l����
M�P��A=��Z!7�� ���_D;{@��!��%7�6?��H�⌗LTOH��$�~Ųڧ��_#Jͬ�d���S��H��=
>UI�\�R�8G�\� 
�����ec�}���$�T~���G��Ut:��Pe��n"+Ź.����Q�SS�e[Y=����w ���������'<�?�K>c�b^�>(A<���.���C�S�s��mݛ���%����"��4�klWr�5��G"������&��Q{�W�V+~���^6�j�:y
�Z�-4p�9��Y���:7���,���|GڔΆ��\���Q��?�����<�E���vN�)�`��4Ǭ#r��
^}�����C��`�= Ì��WaK���`Y�W'~��~
v�(I�O��N#����æv����7\.�K����d��8��(\�Z�Ok�����4b�s���ۼ�.�����P׶���8�&X�(�����j�
����\��%b�]�%��i;D��E��V��`P��E���?A�H<�.��͛?- �O$��x��<�37�I�	��=�K���v��#-�fv���X�t��ʱ�=���٥\ʚ�����<�q�."��јVr���ȴ�.�8k4�bl@�pn�cu�bwڦc���%7i�e�$�t�Iے��T}`�^
������G��\~(�5j[�d���h�X����ܺ����x1*R��6=ov ��i���F{�V���/.���a%�=_�v�B�t1<�w'�O ��Y~1��V��E�LL�	B��QR�Lw��e��u/�-�����S�X^�r~����)9�]<b�
�V�zc��1&���+�)m���v�e��'�)�f�Xd�S}��tr��N��0�8{X|NO�Ѱ������7��>p����	�f�����x([���=��k�ߘ�����bt���a�TS��#.���y�08���i�h�2��bX���P)&�8�)����m�����b3���sw ��W;>#"�w�܈�D����Q(%�^s3e���)gB��:���ـ�hl�P,�?�YD�>�L#bERR��{��oba-��!4��WXJ%
g�t�ٌ�Ǝk� [/��
Ǔ��<@1���G��i����a��gl�o�;$�(��n@��D��;��;)�A��2�?a�ά�g�3���؜qY��6
#x�,1ȋ���}�����id��'�����-rW� �!d��R���#����������:��cS��^t4��pU:�o���E�A6�VDq�+A��c�׽�TĒ���[���^��5ϟ�� O!�,'�F�6	��b)�@[������ŧm$�V�>?����vum�V���A��^
�P��G�[�Z;�-B�c�����V+NCw5V}���mT�7�L��da����0s�a�,Q��+��
p;�~k�,���NH(u-yo�7���-� �+%l��D��UH2D;�}.cs�At�W�@ׁ"��J���#���1@F���?�b-�H�3qi�dW��ݸ/�e���ڨ0�nY�T�ڏ01��|Y�� l�ڏ��~�4�c%+�R˵w�	�Y������~aeW%M�a�W��x͠���:C��1.�9أ>�����=Xj
���T��M���ý
0����.»�L���D�E���	s�}�1d@��h��e�V9c7���l������5���P8%ĝ�P�Q'B�8@h���e���W�a�N6��oa��L�$���h�@��sݓ%��,��L]����&���ת�Fo���2����<62w�o ��&�I�L��m�\��{$%�r > �[
�!�����"�i�$�B�^n܃���C��&/Zn9и����`�2yx��ʩ��4��Y���*V��� �]řV��BF-5>���==�����Hx����gԯ���l���mwJq���9��^����܏��'
�r�0��&�h���B����������@{�V_	�^�����5����{�����׊=�����o8?�U>V�
 �g���s��+i����D�QZ(np�Z�O椸!��^�%�F�HQ�5��fn�^�ۯ�Mښ��a!������r��x���B>_�|
wT�բ���M�� _�	�~�C0��XZF�p�����Jy�JC�(��֮��� �Ì�.kdHԜy'aV��<�r�ҁGC�5�2��Ϟ��V�7Jh��\[[O���f|�fƈ2B�'|�h!�Ue�:����굷m�� aM�#OV{9(�)����7�7�^�WI��hPH�����e�
����* 	���!)����5��D8:��26z�-�N8��\Q�/O2��S?.�o��u8�E6
y�?��U
��_$1(r�P��n�"�����I�����W$�M|��D�L���zil�O�(0��D �ֽ�L��>�QqJ�,�]$�R0�Ր��AO��&������x����LN� �u�Az=j=����!Ԝ�x7��֓K`���Q[�}�ڏ͎�f��~�V�N2��x6�u3+�Sw��*sK@�h�f�pNe5S@T��Zu��v��T���4y$��d��RU�e5���?�Pj���p�����ٲu��\Q���;�x��vG���W�{o�����^C�̓� ��������q��M�?yo�h�Ӛ�j�0(j+��I@��>E�&�u%�:�?�6zp;W�Z��;�pQ�k��"t�|Q{Y_�K���$̜�6U�͹���v�������3���q2�i����&�CB��2�&�q���jdyh�N��\R��.Q!*FSkp�c�"ިyQl�w�#��C{$ 	|���1����ʓ�����f"���4M��Ԧe<��� �h���M�D�bj���H2X����GȊ'�!H	e�v���-o��nS�N�J��Ѝ�,��hhQd%�7S�A�o��4�ɩ���QS� ����Ṕ4��X|t�]� �İ��]1��/��x�S'f�)����Myj]M�
���'�y8�g?�s�$9�IlMmwU��`�;�a)눆E��2���Ҝ��Sܺ��nQ
4�y����8�̬+�N�%��VY�?2V����ņ��m,A#����f'm����1Zܧ�&1��t� M���mE��ܷ���{��?Xv�L�L�Г�Gc�A�#�6!���yY��FI�@o}�b"lGr	�a�ߢ�Ԍ��?D�}0�#��5Ʒ,��iey\�t@K�q���N��E���kL^=ݥ���d�����r��
���v�}�U0u+U3$�֣����$/��.]�KEt-��!��������;O���oI��
JO��KV��0^�D� �C���PO3���?*P 8tM��V@���n&BFk��+]N%�C��#��u�����C���_���$Hq�M�}ԩ�-�Т�'		��ټk��C}Ʀ�����z���q�t.��a��	����*�Pd��oO���^�p��H�$"u���h�l�N0�jNǪ�/m������N=�<U���L,�&W_m;{���o�hJf����X�2'
q�RY_i>��|�a��kX�\6����SBFE�NÈ��? ��~��}���}�����?��I�ߍ��i��@͏�B� `��N���XEq.����Jf�܇�9dd����ш} R�L >A �|����dE U_�;6�9Q̉���Ӝ��v}֠�-��%�k��Z��oW��y�]$���\"�f��怒��)�;�:6�5w{f��%=�ؿM����<;�,����a��Mkx�k�O�[a�iU���ُx�����)�L�0�u����<��P�F�'�yʬ�����՞4%]c�f~�]J�&��� ��3��t_���6#��n�y\�����O����'��.�C�h}^�J��L��qTw�
�\�l�"/�끺���l$s �P2r�wR��Li��y¯>C'M۶�f=���9�b�t���n
� ��|���)��o���"���A���P8B��uu����M��VΑ/�n��6�r����l0?�1s�]n�h-�/'�N�ۣ>�5�Q��4��
72�4%�G��$AS�'�/�G�?�D)�Ѕ�d��g���7���,p~���Yv�]�T�1�.�=��N��w�oy��2����yAL��\9
��ڪ(	���/�'�����kP�s��F��9�pQw'��h���T�JɎhE�^^����Ө��of��Pe�dr�{����b	��:�J�J�ھ���������ȍT�hr1�Ax?�6���ú\3/E��S��B��'�&3-5ح���J+=��T��T�,9Ζp���ďىK��Ǵ6q���=��i�+��W��iNl6�
)����DB���	S�R|��+4T�n2nE����>�^(�my�K7�s�~t'�r�dѤ.aQĴ[A1B��l�����_-_���+Y
/����g��l��0� >(�]ƴ�h����g���w���HR���gX�� R�(����E	��B��sXm>"�S��*���Ts�Y/Sm@rf�:�Dͽ둹���0�!�Ǌ��1�F0 ��a�F��>^H�"��3x\�R<4���M�nSXM�x�V'������6����a�09�Ã��yN�R���"����Q�$�a��mO�Z�Q_;�@�DYSn� <Ku�3��H���=qxln��_ģ'�l��;S'Ӽ;#{ɡ�e0�Iq����^�;�ăv</���6_����m��G/�w$��$��R�V�k3��.TA2��m-��HLtM��EEJbBC�1��y�@��=�h��3�[=a_\��j��t�vad{6�?󺩰~���i����=^����a
�����Ms�Z������|�ZA��S֞�0O��͚ �|>I��L�`wϏc���^����@C�%�K�~W�p�&7���p-&�ާ8�@M��P#�#��ׅ0��xPӺ��ҿ�s�䵣}���t�����p��_��ɉ�����R����)h�j
�h�.���O���hd�D�~ �{m�A
PI��&i�RM+d�y��p�5#��]�ݑ:>d��E\:�.cE'Jz���u<겅 �)����.��0˄�(I�4BKj����y�����sGL,�ԔV�7d��d�ѝ���w�yם4�����;Q,Lv&�� ��n%�:<}��X�8m5RZ��^�f%v�9�D�T�<��A[D���K�dj��]���m�T�\ZX��Y�њu/����[���d+Bl�[����+�y�Т=�9J��z�ʩ��^ei��Z-����H���	��q�jz�BK@����{��M�~ߴ�i�8p��L��Զ{~��<~�`�[��X�
�%���x_��	�n���S��\����xpN��r��9�5�~St���~�̌zi���E���yk6��c��B�J��]3Q˶��z�_l��4����߆zM�	�4/j� �>˰��;��j�A,�IxT��N-+�VܝK�����$x�A��$�?�yv �e��1��5�k��i��k�q^�����~V����R�c�6B*obLd��mI�{�<#��"��Gc��M簠ߤӄ0���u�d_�W�o�^���Q�)-�Y�TSk���A�8��p��*hα8��7��t9��Ri+�߽�{��7���!��oD�]�G%���r��gz��J#�e�����t��]�(h�Q�rW��a��M1�u��a�>hs�3񶁛k�.��@ ��8�U���!�6l�1�&8�c�Y11E$�k�Ϻ��7+�x���ns
[�:���Iz� +�-�dl��IL���=XZ����Ѡ#$�:����}K�}������c�buO?\�{�[�v)�c:l�&D��>���m�����N�+�4*Ĺ!��͛�w/�o�[,H%{��,�l����eMM�w�&�c�a�v�|�&���E�U����u �q�+m�f:����E-��]�|�S�V��<z!>@��tBe�����I�|ѯ��*"(+K ���Ax^�e����>�o�w�/�������� �uZ�ʷ+��kp-�O�U�xY���}�
͎emC*��w����䤫t�(���}��FZ�e�ܔo�<�+	�BMXđ����*3�5�u"��]�-�ܺJz�ٗu�6x��S�q��T=1��OeCC[j�
�k�'C���{���5��0�=�68�M��U�{ [���z�(�zbg,҉E��\��Kɬ�h?�����/�n�6���a�#��:鰐
��@�c�Ŏ{ͱܙF�$<H�w��J_�T$�k�1PS4���bmc��M���S��ܩ�s�#��>,�
]�b� !�� ��M"\ZӉc�.|R*dR�H�IF��Ql]���q<5A�ҏ��~(�����hΌ�!2Jl�v�k������������tx��@�(�����Ɏw��6&-t\���5����8#�;8��f���`��M�6i�	���E ��:-�FF��:�Shi�fsޒ+@ �D��������o#�)��;��7�f���]Ca�sq��g�k�%N�h�R6�P���ǀ4��\�\rI�\ =O��s�'eh���S�q���N2�(�~��D����L����m�j·r��z����/!ӑ�*H��<�*B��w��w�#�db�2��?6��1�r�/�B�i��ɮ}3�K�=HP��R�.�1�_�#tN���֎g.Z�
�Q���E�zCN\1O��t�')3�.�@RV�X7�ZP,L�#�A�vM� 2�4bP_�R��f�ِ����vׯ%Y���s�.��zm�<��q���{��dZ��m�RNzD�F�]��	�[��ަbҨ�2�"ͩ�J�B2��֥@��0#��"3��w'8gc9��:�@�<� ���\z�?ցS̝�����e����˓7Q�fW�}W셶�n�G�ZB��?���I�yX�3Lxy���t=c�$����IFBV����(��Kw��rPnY���ڕ���R�ﳕ�'ꛌi>]z�B�>&/ޏ��Ž1����p�Ǵ#���V�Ϋ;�B����Sy��5��k�Z���P�d�&Y�HS8�)R=5m�g��U˔!߹��M�"�پ�P���aZ5S�|h�n�+Xf�=�X�JnJ��(�����k:�3O�:�z�B����A�P;8"�$r���������(��� Z���ީ�g;B����k~���}���:���C0���d��I�K1�i�i؄��_��b	JqPQ᱑8��/�7��-p�Xw
�3F4!����T]y��M��i��̢���6����ze?ü���i�U��+v�1���C�qP'hyB���t)��S�h�n7q_]E�Ȳd�K\U{x?�Ӗ�������y����뇏�`�+�2��*״��U8۵x77��!����fm�x ��T�/���xy�P��L�W�_�0�c�N���Oz���ଚ∈�'"�i��B�a2��;���,TpA�ܲ��v��"'1ޙvβ��( %���P�}���8&?eow'��bv{,�AidCc�&X_�
�LE�����_)Jt�-l�&���"�V"4�Fˢ�|k�jm����
�,}�.ˮ��T��?2�B0���o@�}�!��9��1k�b�,�!��ȎAA���U]U���h�Ly�ȿ�������ԁ[{2zm0�fXlh�\c�I"�K��U� D��B�j��Y��j� �8Bg�럿\���G��!.tG[��E4>���t�qS| �;���:oG!��\8�< �D��Q�,
M��z�Y�R�N��NCo��9k��}�ٓY�t?x�Q�ny��ha�	i�{6 )	�A%��Zvj�^�d��U�ې0���`~F@��~'�
���L��_�[�R��W/��j�4�-���ݝ���@R��	����-b�`}�E
(e�����l+�ٽ�*(��|
�`f������f��� {��i;�^��Շ[�
T!��)>��A1Ҁ��Ќ�^~*�����b���u���r��*�~���]�K������4R,0���E�| �����^���,D8װ��o��*����,��<;��ݏ쯩i���v���szM>�9�����Z�K���-\�ӣ�~�ؑ�^,5m�т�����G
o�}1�b�v	�_bu[j2gʂ�RlײV�ՙ?�������D68����"��/5��'p�2*�������1mZ���ê�̃��(Q�a�!� d��A�r�/�	>�/E7�x��0�|�*W�7��-]Zk��ǐ&�z�?�Dj�����\c/o�T���3��m웁�Z|���n�p$ՒH��%�A��;�5�Y.�./� ��x]ѣ��OS�ݰ�O343>Γ�h`d��{!���ިۍ���֕8ӓ�v5�C~��B:��rC�:�����:̠�r��ûy{-�'c3 dPxF(�������������K'eϫ�� �t��I5�VΕ�B�	����/t88&\� +�̿��_��δO�5]W�$��c'��Bs�},!J<����=2�������t�;�B�&��`�o�jy�+�K��<(�Ɍ���Hx���P�7���<��A��Yo�sqt`R��vG�m�ӟXЖX)�+%�|�i�tB�u����7�'�憲�|��(f6��9���=�e�xK�l��/�� Sb�(��:cPV"\+X�Ŝ��"�R
����j�t�������$��ai�H�D���nba��2Q�f<H�̭cT@3����2)0��@�	��X�\���O�k>�f���.F�M��|������"_��a^E���˔#Çdxp���7IFRrc�Q,�d�J����p	a�4 �`�#��nT��%P<IV!�2��@+���ʛ'�YXr��ZI��a��Y��g� U�
&����}�nN��r��-(�n��
�� �!*�
��l�_f�e�<�440���ӊ>�;�(=�g,5w��9:b���З��͘���ǟ]aH,���	q�U/(1u�[Y9��J<��?�j�7A&~GQ��ջ"��(��"�����K�gI}�c�ظ	����DU�ա����]�g��N|���◞t�h?9�B_�f ��Q$�g�Q�]:Ь(��%�Y6m]�	��� ؀�&�V����
��*CE��h���秢J��=���+0�&9����b�cGV9���e�&���!+�7���5aQ��OqV��I��*��?o�_]�hwi[����[�'=`�9�����.;NI��|
S���v��������B\��?�_O����O�T���� ��Ӆ5F��x'̋C�p{�$�`�p7�+��<���gsn۬lE���+��@��r@�7j�J��b� t+�/ �l�T�oɂ������������ul3��`��G�9=}Yj<��@Mjq��ƿ�n�v\"���M;e�\�n�٣{$�%?W�vP��Rlh�΀�5���w�����VEf��8����
���dzZ�����'D),�dl$��߅&�q`��l�to�0�}Q�x�����B����=��R�]�S�r�w��6^��?�qqb�b��O��'THӸvI�Q��p�%C{�S�r#��{Fq�.�9�������o�"OB��cS@j�՝�2�yh�����V��?�k�z��Ke����ٗS���i�g�􇿣����R��0*t��̻��Ō<�e�i�K�f����)�"$�@�6�&�S�o��������@RUB�Y���k�ʽ���+>��c��*(�\:��Y����3���$�����v�R��~���jU��4j�ٞn�K�
�
)�1Ki��$�5�1Y^$.P+B����q]�4�y<��A�eH��ճ^C�L4ArC�V��I-�y�X?����5�{����Y�o�NY׷���uZ:X�t�`fד���O��5\H�/�q��٧��^�;�P���)5�8�"��w*L�
`��RF6&=Ƕ(��sH0�������aZ�d%Ч��s,��Q���G{����Y��rNէ+9��l��^$�~U�>p�K`�Y�g[p�w�P���$D �^��h��ۚѐ9X�x�\J����ѕV�LF�.�T�O���r{)7
hH��1��1b��Gٯ���x�
� �N�����{Ξi�ȤP,^���0�p�Vk�7���3�|��ɒ�j�2n�B��ߥx���"xvܨ	����Q�s�K�?م���΀�܂�/�G5�vMU�%ܐ�7���jv�'�ǥ
��P���Bᄈg��(��t>�a����V��w[8.l����3� �H���k��⿹�IO��Ù��ʥ0��ky�������9ע��0�7�d]�����8{�_�;�\,[�PUBy����a�a�F4K2ʑk��~O�����[Kb��-�#�)��1�̊@G�3�/�(�׺��6n]�ܳ�N۬�%(B6�R8����>����34���J���j��tYs��{���વ�ޱ�������A�S�Z�`��R��~��7<Q���BM7�:X�)�:֥^��%^!1ާ��[+qN7�|Ä.M��P3�$MA�/�*�/�� Fs�I\;)˕p�H���Qt� h��'}c�ЙΌ�4-��������T:��Q! ��>"+4����3�@!�7���O�6u!��1};l	��	�+7I4�6!	c��Ndx����V���,~��l3�tV^���4[�Ħ|)=b��ɓ��Ϲ�
_��y���_� fC>�f$�hD�%���eMI�`ŕ��mB� /��,k�.�<h��$�leՍ�0�:%���d	_��`2�����$Q
[��!��r�WiW�A�j�?�'l2� �V�����¾���8$�8��H��MR$�S#�p\��y�ê�7#o�G&�Jzd�i��9���Ż�m�Cc17�����k�T<j��(U�mS[*�����ּ�x��a^��r��=T�~JL*����\��䋢��z�&�&k�nM�$r��*���ϐrd�1-�/�5�a��P�(����p��[��^U/Lj�R��Rɐ״�U\ U�zx�W�ߔ���k���Bcd��*�vq�7�[|�Qw��6��� ��Z1�$��U���6����͟@�8���Xx�>q:�H4Q�����'r�Xb+�Pi\��v׏B��*���V��y�㍼.�
B�j �DD�Q�;���,=c\��`��Y�3_�����7�k�bl�s���oJ�q�~��v����°M��n<P���c֒Y�~�y���r�I�_H鋋&�pM=������ҀD��3��gx-Y�s�c
%!���Ee^C�Df�bt�6�JϺٺ!�����H��#g�ATm�;�L��s��nb�^ڳ�i�h��z��K�\!MH��I���O���x��[��P�Δ�D�|Cf���u�'�
��9����(�Nb��� ��'��u�E�<�y�^"[��s��_Q�cď�-�����d�e�jW���\Œ��?3��E �7�1��[�/q\����
?ږhL$ �Bj�z1:�W������� Q!����@�y7�-�})�Ag�l�C���$���o	���I�����Q��
2}��ۨ��y�����e�3��ȇ,TT�顜�E�ad��j��o�������M-��3E�G�MR�X�j�k!r���4���B�ջ㎁o�|=�@n+28OA�q����6�;��Ja�^Q�%�
��|�x{�#���\@فE��u�|�pAS<��5�oU$ؘyEo�9���7�`q7�'Pz�Y2׬��π�!�p�w�a%���:s
xҐ4$ׯO���Whq����Za�v7g�X(�Q~X��1�E���yh�E;�:��2�ߛUv�[��T�=fC6�����$~�!4TR�p�-��|�Z���q��r��c�R���7�l��Ɣ�7>���!B��=[�v���ҕ�<����rs,���g������ĂU%�3�Ew7���)��s2�ZA�bK�IT|%�b�֌̘X<�͌���0����9���'�����9.���)a\�
2��K��d��F%״��#��֜���Oj1�������x���7{\ݺ_k�]WPI9+�6o޴n���,�_P�ma!�҂�jc�Pi*>�\S� ?s�j�z�\�t��_s���l��+r�;��婄3��g��%v�7�U�0n��� `�s��W�-V�Ak�A�ʼ�ʿ���7]�<�~�g���#����5i�������Y	TY���K��A2�␶�>���l�Ȓ��+_�@�}/���"�al�"A����@�(��^y�!�23*�|j��9@����HvDy k!~N�f�~u��u�u4�%N��<]�I�p�`,�J��"��Lӳ;է����5���C�]�v�e%��}�48�
�k>�F�����,�EE�o'���8���^�����0ُ��'M-�ĉC]��Xs�+��q$��%���ߥ�~R�7WFg{0Q�yْ��a7[ �Ce�v�X�zC��e7 ��P5#k:�w=}!�Lq�|�XvO@�?5U���YF�N��T�.�˼�kSa�0��2��2K��sk�⺴v��1�� ~�~2�{AX�3b��ⷊ�����=p�o��74x�t��1���^���奊�����%�/�%��k���LHo�k�m�h���5i1�t^�W������A��7X2ֈL	M���%ǺI�E�Y�1yulE�����6ut{��z�J8{��[�R��v3��Nf̮��[>B�{�p&큒�`>��t��a�H���ԉh��]`�֒Z[��]7��:�e`�
�iv��GSΓvHL�Q����Bb[� )<e�����p�ޝ�+�Eo��&��b��2����<l�.%|Xf�{QH"y�� NeEo��,��{����<}WE�e&A	S�.C��զ�큭�ʌ���Bpn�i���R�z>^kx�	�x����2��v]d��$j��n�G�X��RN>�s�ΛoϏi*��~E��DI�s��-�8`@���y�,��B����f��X�cFp^L��p�%�����MRy�o��13��H�V@Zw�r����3�,26yh�I��;�@<j&~�(S�[��?V�� ? ��8�>���D��D�[2b��Z9ܗ����,,�������y�fR�o���hy`iŖJ 1�z!��c�'ѿ�h�)��R~��#m4�\�O�P�i�/�3�)=d����̪������G/6_u��E�@4�x�&���]�p5h��K�zX�9ڸ>/�
�Ue�ꝝ~X� -������+��8|)>N�����Y��`4{	[��P[���Ɛa��w���&���đ5��Xh��'/�H?���V�+�=��ٻW���7M��L� el��a��%"��=xᶩ��a��K�Nt��AQ���Pc�&��ر�n���$���+cw0��l)�W��c��N&=��,�R�S4��h�?�Zﵒږ� y4.�=q���[��������{.�_3�亅��N�/-�2�\�������!ϩ߸.>�
48�|�d�u�?�jk�ʏ`Y�>��En��$��+X�WP����5������#���};�Bj�I�;����W��4w	�4�Ɋ������������VLg��*�E������rN$\���T������WXTFH�]Qk-Ώ�����%��4İl*��Hm%۲�͚��b�m����wen��I[/[X-���?P1|n��T��r�y��Te b�]�~��_��!�렞`�����>x|IT���i�t�~r[�m�]t6��V��W}b @D� C����7_�?J��қ���U�5�0�6vۆ	��s��N��
�}�7m���ܦGda4w^�������Q�z��׏v�$�rFg�|{��xmYRw}5��zq�\8���4ʆm��`0ܳ��3k�ґ���9���:�U�n㑧;�S��`AiƸ��$52�7���-���ion�F��J��PG�cX\ޓ���x�L�\J_�ź�c �p �HFԎ�RG!�~����|V#���M(
,����o��9�������1fu�4�;p������LVO0줊�MI��(���l���m�J�Ƭ�vm����@s�	 �7}�7]�����z��Q�c�K�z�|0�P%)õ��]HAS�cEO�g(Z�.��'�!�
��G��(ܣ_�ՆZ�"�>��"�Ԗ.��S��Jt��{������FI�u�O��V��k𛫻�$��7��3���ڮeK�66�K��m��u<�i�h�K��)��r�oY���������|[سi�K�+�s"p�%��L����t��	�J�Jw��l%l��@D�!�ߘ�^�z�k����#��"|&]>�5��`鈯��j�,�dEZ$v���u��/]�� ��:y7�	\�4ʿ�n����qݸ
r-��X��!��q$^O4�3j�0Xs��m)�ߛ��O&�� F&&dfj�>����f/^���d�:ͫ��W0�$+m����l)�a������"BM����۽��	\h��޹9'ƭ?(}Ts	Y.��r�₎�E˰m��>�>*���4�%�A�z%?e���3BC�OǤ;�I��:�c�=��F|D���Ŭ���y����(#��x���S*\�*V޽*�S������W�D���d68[�0�w�k�{�Y�N5ά~ğ����=��M�ub�*����_�O�V�x�϶np7T�Blo���/2��+�7��\��g(1�׆H�G��EH��O�U�bl�� 5\����ؒ�ﱪ<��	]WDX��)��6��cV�����Kh����P�#މ�n�Y��(�r�G.��	���9���BHJ�EE��l2�p���l�KmE�L%ˎ��<�.��������&?���I����=f�X��ZX^��ln9ɢό@c�<�`�h�Jg���+A`=~͑��"Q�Mk�t��x�����kR�\f!.�0��)=� �^%U�����PU!9�;MV�DW���PK�����˄k  �ŭW��g��������΂X#AS�r��u�`��Ϋ26L��(��S� m0����9���K�cf��-����u����ə�D̂[��̞���VzXGU��q3��K��Dˊ�����O��$N�eP�Z���q��R����c����Jv�N0�WT����w��w��_�A�>g�R���-���wU�j
73���W)���$,:���{��a�=������2^���)��`^�h�!�de:�6�4F��=���7Ti~}�p%u٫��:�jL"ԕz�)p�����]]ͫ:絷KY,]rWα�p��90
�խ�y��KQ2!#N�~���K$ʪN��!p�3Gy�v-�8$��.]�O6���M�F��b6 ǝ7��Z�8Dڈ�ޏ�}�0��l�+I�;� 'F��8�÷V�F�,���T\����:պ�C����*�I��<���uI[7-X�ن��Rf�:�2I@�U6|U{"�Dv�3�38s/���HzB����3ϙ0q7��gGK�c�S�Q��d�&R��q� 7"�x���#�E�@�uÏ�)��t~�	@&���ȁT�?E��d2�B���>��҂)��c�4�A���zi6EB*�#���?:��Rh;���m���<z,��]�0������\����f��Vzr���{Q��潺�SbA3Y���ܺAb������'���`O!9V'��'<>���S�w��:ČO�-�*�I��,���õ��	T#ZEqQ�-��v�,.�Z���0�a��q1�c��� ��auI�n��WH�.�^�v�Z�*s�"��j,�o��{��z���>;��
c�6��K�n
i�`d�t+��%�y�l��ez����O���6-Ax\�}�G��n�<ۘ,���e��c랐����J|�T`��%� 1̶��"�l�Q�'EBc��!V���Q͒f�}Oz-
�w8	+D�M�_9���J V�`p������9,��܂@�q~��=�r���&��K(�@�ͩ��A#\���&�d C��5��G֐ɽ7S�#���B|�i�tڲm��c�Ӏ�)-~"��<[p��#�Cy����1e�Z�6{/'�3Y���1�酈�L�%���"�<';��^*�ź�)���V�D#Pp	����s�	$z~�B��M�&e�G˞���R���=;�3�6���OV���d����y.��N:�����}��ͷ�g��]L�rGr���ox�a�p�a�K���$�%2 1��`���wZ[�����V�@��b1��SR�"����m0��������]��a�)�9�UH��}z �q&u+I��ζ�v�W�\�T�����I��a/{���f���H��Y�����-�x���9���O���&�z)��l�m&Y�:WkG�k�&��B;�ٛ��Z�Jo�+fP���Wbmة�X�}�F��kK�t=�Jga(_��K�D"!�z"��}a/$��/��e�f�9t�����o���ȆL�i:���r�}+?\��D.�^��ވp0��7�Kzj�4���=��9s	5��DoB�f��M�����1�˔	����]��]��WL�����ǭ��/�X Na�v.�8����K�$�(�Exa:!�J)^�hŻ�뛫Jj�j�=R���"5-���=?���Hd�=�9���P��@�O���?��ye?	c/Ӣ�T�ڥF����~K��-�#���]0�u!�?\<IX="j�j�r�� �喽͊O�S0,r{z�Y&)RE'�}w�S5F���Oω�L��'s�*�q[�f�_�sp��x=��h����[� ���~�9ӫ�;���(C.ʗ����UH���k-$3�F�)Jd�ۉ�T�Ak���ۦ�����p�r���)���/�,��̫�xS��s��ƺ��Kk*0"�.��}��<?��u��ϘWËU�Ũ?�{���&�S#�kRW�V��])kE���B��r̞t��{o��۝NڡX������� ���j�es\k@�Q)H���@!Sן��ǴB<���z�����s��A� 
C)-�<�gcE�������E���E��@��}�r;DG( �����k��4ߐ��c���uX ֞]������0�ܪ�(�,P5���ήۗǼA����9�}�j��),�H��N%-����濻M�h�,����=��S^��``�f�Hv�JD�T�b�.8� ��wn� iv(Dv�m��e{�G�%��.�LF"��|��a�U����߼8秉Hd�l��@�; kX�B�P �E,�)��~����Q�>ʼ�^6�2+��mG;�pq$HI�������B~Zo�7�`� �}�����0Lc�䴸ϯ���O�&a�ҿ���A����f-L����~-���[H'<�.g*������6 i�,>�.��v$?Y�ݗ��vCp�������Ba�:����/���hC��]ӏH2V��"��t�ݻ�N�>��삁@s�rV�K�>��tA��鍜cz,�1nD)�LW~6f_Q�87��l��q�y�J��ś6�XBd�7lZ�A��G6bF�����[��8�:S�\&�賴j�8�B���Q@V�&�#�ǻ�{�w��=vW��0b8�"n�%ZD�g*��"(�U�
Y"hu�d	T���l�K�z�?�2UK(UE�f�;
	SY�lj����s�}���݆fʲ���S��7>Õ�k��Ǵ'�A���ν�	�V+��ⶂ6+������DҾ��ݪy���]���xR����Ci?�[��W��7�F=�(bu�nC%D2��m4#/�t-��h~kc��Y���F5�s��6
����.F)�7�:4_NYhf��F��9�鄪�	����	jB�6:$��A��~s�r�RM�㞄"�#� �� j!c-l�:zȤÈI,su&:[-I�`�pU�9�Q԰7��!���W�G��Nu#t�ĒK��*��&d�c��t�W[;�K��iW��!Bj��&o��L�x��,�֢iL��T)����ۺ����e��g��z�(�CCa��UΈU�Ō�І��㑱'�R�2w
�(���D���+�>��An{�s�5kl���Obw����:ꎖ��[�8�??c�s�!����-Ϯ�BtI�GH}�ǳ��_%��s۠Gd�q�;K�iǵC��#&��/M���K|"�q��%������RC�l�,�j~�7�p��زI�b�]����Js/R�A�G��v&bk&�����xM�Tk$�2K�u/�5��tI��-	e��x��%k�m��PT�ή�������jhњ�m��t����U��tL*g "1i7�g�6�75nw����p>�>�4�;j�_��Ċ�z�R�IPu-Y� ��|�:�������l�/z��<@����䦣]�ahD��pM>��H�A��ȥ�>&������.1�4M{�}x�z�Լ�� U�_!����w�\S/�]Se_�������0�7:�}yF��}���-���q������p����]uV�T�0�o��H�C�oFͥ�Fp�K{}y�=�yP�Z�@��=G�T��FҦ�1ƻ�d�=�2]��R8Qk��'�Cf�z�㍴<HB,��XGq�}�u�7de���

�(� ���,�̈́c!	��Xf��D�bԬ�!>)�0�3�M�fZr��� �����jk����Ɏ�A^�$��,��l�)�~���Q��8��7�m��Ke�ҏDm���dp���ě�ۥ���!�j�(~��p�)E��]����? Y7�$���p��6��J��[��bh:��`�B�#��!F��W��	t����r���ՙ�g���I1�|c,*��n}!�s����*.N���Y�R�T��|�-���'qT"R�(l��D��7A��at�$���ν�7��8����C�b|�6^��
��`�fr��4�A{ѪP^s3ܡ�*̌ȍk�b��x���ɗ>#?ԛ!'̑2��`�4��\��-�ST��7n�(ۣ[���³�Յ���M��Umz�� 5a��(Q�#�?�b�3�{�����YH_�S�
��Ҙ���u�ݗ�1N�̙3�$:�U6^m0��Ț��r���eYI�2uQ�}����j-$
�r@,����-�ֺ���[�@���3/��q���ڏ3G�ۡ������0�݀h����F�DԖe��11sB�W�}XKq�&����,BB�����;��F�Q������Q������"�N���A1i������v��yH�̵�*�{��F@R-�F��.����O��ʛ�|D4wD�Mr�`�rWX$%����p�;���g�o�b�Ҵ����-Q�aK\�j�����Q�M!J%E"����K�>ab��I��t4mۜ_ ��'�Z���5U�8�y��̼���A�u}&-��R>��Lӹ�������+-�a�9u��ϗ��A��6��P�!��k0B&�����p�D�q���X�Mάq7Sf"8i�i��F�|oR}�0J���ho�9��l�[�uD)^��A5�;��	��i<���Q2p���b�Ӓ�q�Cpt��	���O�����z��[W�i�o�M��EO? S�?5� D��z/�e�:����ݵ!��~�#.�i�ޫ��+�{7~��\����V�=i.��=����;n��|����\�� �����d�˵T��0�sG*B=�4�����I�uw�D��fHMHX�/r����H���oG~��a^�����;����kcrt�e�Cya��>��U}��b���Y �K�$�=?cⱳN��*��Ƶ���bc:�#[c&0�:��D�ccֱ��EB�h���A������H�F8�f����숱�	�K����L5K�-�1Ѿ��X+�.�aя�N @.������ҍٲW@��K�'����(���t�Z��W~pcQ��� �.���{�̈��US�&�����>Tn"Ij��,�[�!�R�`.>�r���=� d�Y��g|����{@�9O[6�N.3)�����v�(�;�V6��i0��<٦,'Sc��M��h��_�����j����c�?������������pkVXjŪI	�Bd^qE^�6%�"'�����������ib;�?��Y�"��Jo�(_�S�:U��F��(O�Gp��`x6)�@l�"�@?MR�:i�zF�R8Ș,q��$m�:3��>V@}1�E+^�1.��c@��Q_&�����ٺ��n����w��������,zk��g�`�7	��龒�O���Z��(J�H{Ⱥ2��g;�Z�=�����8{�" �ZL�|j� �!�QI��Xo�j���+�$�Q�!��;P?4�F|�ڿ6�������|�E�FۣFhR^�?�Ã0����jGT�Hǘ���ւ�Q<�Ǩl�O���p>S��
���r�>Ǿs�$o�=���t, ��z<�;c�,�!��&	XH���;���m2�h�`]tx�|����Rm�f���qN @х��l� θY	�VEky�C�/�&e`"D�X�bL���T�+i==�1m���
�1�m� �E�̇'�� �Wե��R��R�S�8�d����P�-��|���7��J�v
()�T�� ��,)8KT�Wӱ{Ν*�����r�0�E��Z�d<��K6i��OF�ҙ�ɐ}�	U*�zE�t i�fh��~�g��/]	���0Xћ+{ͨ"�LRlk��Mq�yp�v�բ�ɜ��L�9��S�J	���z-��|�%��5� W'«X�B9,)>���bj�)0*D� j�L�����L?r��)9</_�l�X�+4�yt�zt\S���7�p����D�;SA
���sw*��yޕ�a�6�W���?�O�%
.�mb�\g�,ՠ:p�B�ܴ㯇L�
�`"R"C9�zu-�o>�>��f��ly��Qt2�<Q�O)3�j[��r>�Mv�����W$TI���g�S�-�r�1B�,�l�VǵSw�V��#��d����S�5,w�8Ԫ���U�^�]Z���\5�g��n�հB�����\lZ�	�=f he���du���aSjM�);nZ.Ohue��y5l6�U��4��v�=�#��6z�g����9�^�����hhd_�UY;k�wҭd�M*�i(i ̿"z��az|f�'��Lx78�_�_H<�O@j�^�&�A�s5�d�8���{>>��^.��z#0�vx8���J��r=�>ڒ�p8�B���RE"7xz
���lP�̗V7R(Ӹt{��B_Z��ּ�34O��/�k/Zd�
�31�y����q
�P-#��Z�O�W��(o�*���C�WwX�N���V ��pߤ<	(�R0��}nt�����e�I��z�4#���w�IAok�q=*�K��t�/�+�*X�"��7��p������&ڎ%�:Ɖoa��i쀌<�������ǚ�W��w����XR=�p��^ �?#� �2Re��+���V��/iBR��es?�[XӖ�TYocFõ�Ƃ�������+�I�/����|�������Դ�T�,;�^�2��^��O���������\4��4f�P���Z������&�Gj�KGJJ"��;d!y������^�7?�������Y��ۜq�&Z<�����J9�i6�b��(�& �2@���. ���u*�p��R�L� X|j��h�͒�i��&��B�a�]B��I��[˒��N$e�_u�k՚�,֜��)塵���k;�Qi]y_�O����<�=�Q���Xւ�ѽ*ҏ��n:���k�I�'�E�d7䚫j���`��cw��3Q���L�@���S84�@\������d8n�i�fuI�,)	x��	[�r�1\�\�urk�hh ƈ]pngS������� �������$�]i�o7!Q�|����@���)�R��������jR�ӽbFX9 �U;��E��~��(���k"��G����j��}�z�
�2��9��^��䶨�~�J�>��#^�1b`2[a�@9��� �P`痝�R�r#Q���� ��z��m�i�3��x�l���j����biI��[*�Pz���%8ǔYmJN)㤎��]�~���x �����eɝtl����:�*d���h�f���	p�;�%�'y�HҸ\�l���%`H���H'�yM���u}몼�\ ؊Q��Ѕ���iُ�J\x�*b\��3L���
�u�t�:1R�W=n�=����[_����5����I� ��F�+�k$1�1�Hu�X�*��v�;��#8H;�����2q�i�\��,�!
�L�{_v���v0�T`T�|�z�Y#r�ZkxS3h:�4� �T�$�)���î��[�l����Z 0�*��!�p���,���|{��lt�<�QI���ɏx ]B|�"�3zՔlev#_EN9]�%�W�\��A�)n�'�|�jqX�q���"%@���A]FpkHa�
a��93
�qv��d�IƇ	P��ˋ�K[�C���RV��x���	��	P��;�_�[»���^M`٪�* Z�mi�.J:�>WW�(�� ����z�j{�<T��J�@�ѥ4n@�� ��a������)V"��p��r-wA5�"r�C�	`�[��=���R�H���� "k2����W	V\:�1De�-�u��(v�F�W���V?s�5I��#�޻hZ�u�AN�spncf x q�A:�������&h��1;��H�U�,_���{����6#f��m����@vX�s���L�c.��Xڡ%������=�����A�<3uf�:�ʀ*�T˯mU�?f$�Q<-hIG����R9�L%*��]A�A��Y�V�\|�ͦ��$3�	Ъ�Mݪ����ǳ���!�^�k��)���Q�;f�!l���~���v�v	2��Kd ��f�o?j17d�O�Z��p.�+��k<�Z<��C��,�Y�����G1q!ܒ�j?'�e��0W� Dr:kSȪ�� �r]4�C��=/��j1v�]����\����6�-R��i��O�H*G=�G�p��`�$N���Dk������TH��_�
����)NR�PS�Ƒ	����S�_�Y0�f��F�0Z���a?��	-��:W�59����ժ'H����ȫ�V�{�|l���S;�}r���7��ί���Ȥ�8D��Z��%��kʟQ�t�ȴm��S(A��L��;��Bx~����2��E�A��m�6F�b
Ta��/�)6(�[SV|�t*oHg%c��ƸuL�+�
~˃�"_�o-�]�T:�L�$ꠜ80��4�c�6|톟�������^���y`�pHI�.�q�8��u+�4jg��ە�r�`�̓YY�/uv	J����jz?����cz=��&���ѳ�!�t\�]Q��5�v+��<Y��v����b.`ց	�y�P_��r�_yLDub�/�}�ۢ�i�~�e��4� ��TN�<��8��x�9�m��j
�(F���B?w�O�Y"�{���g\������G��'J��_��9�k����2]k$<�0�W
�3��ph���9�M�ٽ����#6\�߾!���(���R�>��c��h�i-̹m�R�y��0]3I���KLo���#!�F%H�\Ha���C��8�����5Wk��3�*1�wɋZ�硌������k��%�>M:����{>��Bk�Y�3��B)��P[5���l����P�e%����V�ej�c{s��U����;��m���'"?�hIad��+�9���:�1��.G0���l��H��<�����8<�>���^��;?0���{��g'�=��}?����u�{��0�Gg��ʒqKy����*jm�Q�<�	|��}�$?�{`����\"��ڭ��P�̼�.��y�;8=���'��s�TY�>Jx0{�r���P~n�̮�����y%�!f��r�I]?qk{l���h����'�j���f:Q�A��K�='�4�\���R���'D�s~�����)����e�{>+����G|P�-d8�e�/�vۄ���D�4� �c�5��ooAC����z8�\��	]�~e��cYt[���>�o�Q����
�׹2P�fg�c`f�9g�}\�rI\������;�}��1�Rx5���<w��5�@4�ut�q藤����p�I17\�Di�Ht��<J��_yD봸�G ����FLv��ҏ��`��ڹ���$����5�ʺ�+hf4�p�4��ʘ�0��9�L�ƨ�g���<��*ؓ���MA�\8]�	��n���5���h�THOG���e��H��4���Ha�b�X����b�	2�2�ը�)�T��G8����BZ >�6N��1�)������습�	5�����^��5'u�5U�`~ժB���w�M0W\���'J@���A�G�k�	Î���V�v��dy�Ō( r�aj6Ԓ��WE�A}���rRS�e�YQ��p,�Mht�VL���2����C�\a�T�x�4T�4>h��-5s�Csg���71;">��ߩAgv�Ջ\}�2w<�pefLl:eA�'���[��ws�A���
8��Emn�hnq�Y|�S�w��R����k�i�1_,��~*j%��t�Y��� Mq�R���m��Ѝ���}�bB���{#q�o� ��Bd�_+����g���?�P�TP��WY�O�N��o�4د(�1�u(�K�����*k�i-��t�5��y�ӫ� O}|-�� �ֶ�&K�e�#-��͹3�)�;��L��>�_��������-��{��^G��3�J�O�z��1!�	�q���B��_A3�]��n�[��>+�� �^��X�&#��4%���jN^c�M�!�MN4!G���X���d�&$����X�Xd��=א�ȹݔ�N�۝�oD��*)D�-�jYF�POVw���s��,9_���� ���W��Tܘ@N��R99j&Z�Wͱ���֠s��V<�q�����֦��!�������br[k����?���-�m!�D%�w��6��TA�N�~S�@��k�A��9!���ox���O��uRD��c$.9��Am�AD����C�<#1eG,���j� M���鷶f�6'o� �eK�
Y���J��#��K֓T��5ꋿʣ�+�\����KR�K�s�hFT�ֆ����?��{x��\h�(�M���m���/��CO�D�����Ѩ z.}L�v��s���xH.Uױ<Ƅb���/8P>h��tn�Ӥ]4�ĔbeX]�+��u{H��]��*��U�E�Q!��y(��e"D�%�6��ί���2�`�R�fD����e�"�E��o`R�ZUJe	]�*������=�{�(�;^���[�������8��6,�a�.�	a:C�={5�l$��	v�<Y��+e��wS��՞ؽ����覘f���`�S�/�e?^������M�n3�R������q�nf��m_V&�6Y�=�$���nJ[�|;^r6<���¿r��9��;�%�b�-��o�@�L�:���k�cΰ�Qr�OGC���e���sHP���ӳG���p�L�.2�ڗ([#�/���L��#��7�$�^5<��%�>����΢7��h����ڔ_VbR���X@��jx����f�<_�T�����}xVГ�݌�|����?�[��R�l�(~�M���������i�K'����e�%-d�16D���Z�V��������O"��x�,��{���������k�����ف�ws�WO5s���`ʔ������b5^�����gǉ��Z����Y�|D`��ʔG�}�B���s1{
,.9Q̣���nƶ��ȸ�K��ƶ97�������0~;):��0�1�6�g:n[�.QyH��먂9f��dٕ���IF�M���:�X�N���o	ߴ�"�S�u�o�� XtۂVm�F#|�yǑ
�<դ�u,�+4׎���ń;҇�w�������J��Ϗbp��\�=�a8�!&_�<�m�UP���h�hp���]�*�̄Ƥ4ʘL7+��.͎�S�F)�j�v��'����T�g_waN+4Sw�w� ��q\4��Dg7�ʳ���&u5�Nx���V�ҤC�F�x�[�S$ё>���N2��j ��b����eC��&�j�,��8_�S��*�bD!�s�P�X,�
$"p`��+���XH؀O3� � �#�ݰ�����S$�E�,���{}���dC�&_w���<�r����S��%�6��h�4�v��!b_�(�$�S�J'�j����JLs+j8Ԅ�:�F;4"7�?���O�Ns�7Dx�����)��!�����}zs�?m`'$��b���31����p��J���wv�k��n�
��=,�>'Q-/[� &3\-Yb,��C�_���W�Ե0b�<o�"����P���wYg�8`So����v�	j헁�0�=�N�	�
V8�|fN\�~ɧ�
�bt*L�l��דm�QcB����tz�o.쩏]]$@��w��Ȟ��"�l0i�y� �L{�}��q��d�v�gy�G�Na{��}쀱�y��m��ֱ�P���o�0�N9�t�ڪ�8ʆ�9��C�"�;-%CQ?}"dI$6�ho�):�{�7�ZD(Ew��SA�(Dw̰��\�Y1ؠW7AE˼RZ���F0�;~QQjEC���fז�}
z�B_O8
~�f"ӦR��Q����۠�|\Nc��@Y��/D5��f�a����fԭW%#�M9`�ӌ���{m>�ڳ��'l�İ�L3d��z${�=��/���W���=�8ŋ�D#�$h
���8���Jn�Z�._�,�,��]Emr�mxreV>T#7���5���nP� ��o�%#v�0���ѪM�����pJ_u�"��:�j��f���U�h��:<�ڙV��nF��}�Y�C��� ϑ����@l��%D6p2�Һ������1 fBr���	�N:�'����Z���	M�W�8���t]?E)� ڰsq�(�0a!�H�F�n��n�7�3x��9�e`�poX�SO�9�9Yk�ru����s�8f�