// (C) 2001-2011 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// $Id: //acds/rel/11.0/ip/merlin/altera_merlin_multiplexer/altera_merlin_multiplexer.sv.terp#2 $
// $Revision: #2 $
// $Date: 2011/02/20 $
// $Author: jyeap $

// ------------------------------------------
// Merlin Multiplexer
// ------------------------------------------

`timescale 1 ns / 1 ns


// ------------------------------------------
// Generation parameters:
//   output_name:         application_selector_cmd_xbar_mux_001
//   NUM_INPUTS:          5
//   ARBITRATION_SHARES:  8 8 8 8 8
//   ARBITRATION_SCHEME   "round-robin"
//   PIPELINE_ARB:        0
//   PKT_TRANS_LOCK:      72 (arbitration locking enabled)
//   ST_DATA_W:           89
//   ST_CHANNEL_W:        10
// ------------------------------------------

module application_selector_cmd_xbar_mux_001
(
    // ----------------------
    // Sinks
    // ----------------------
    input                       sink0_valid,
    input [89-1   : 0]  sink0_data,
    input [10-1: 0]  sink0_channel,
    input                       sink0_startofpacket,
    input                       sink0_endofpacket,
    output                      sink0_ready,

    input                       sink1_valid,
    input [89-1   : 0]  sink1_data,
    input [10-1: 0]  sink1_channel,
    input                       sink1_startofpacket,
    input                       sink1_endofpacket,
    output                      sink1_ready,

    input                       sink2_valid,
    input [89-1   : 0]  sink2_data,
    input [10-1: 0]  sink2_channel,
    input                       sink2_startofpacket,
    input                       sink2_endofpacket,
    output                      sink2_ready,

    input                       sink3_valid,
    input [89-1   : 0]  sink3_data,
    input [10-1: 0]  sink3_channel,
    input                       sink3_startofpacket,
    input                       sink3_endofpacket,
    output                      sink3_ready,

    input                       sink4_valid,
    input [89-1   : 0]  sink4_data,
    input [10-1: 0]  sink4_channel,
    input                       sink4_startofpacket,
    input                       sink4_endofpacket,
    output                      sink4_ready,


    // ----------------------
    // Source
    // ----------------------
    output                      src_valid,
    output [89-1    : 0] src_data,
    output [10-1 : 0] src_channel,
    output                      src_startofpacket,
    output                      src_endofpacket,
    input                       src_ready,

    // ----------------------
    // Clock & Reset
    // ----------------------
    input clk,
    input reset
);
    localparam PAYLOAD_W        = 89 + 10 + 2;
    localparam NUM_INPUTS       = 5;
    localparam SHARE_COUNTER_W  = 3;
    localparam PIPELINE_ARB     = 0;
    localparam ST_DATA_W        = 89;
    localparam ST_CHANNEL_W     = 10;
    localparam PKT_TRANS_LOCK   = 72;

    // ------------------------------------------
    // Signals
    // ------------------------------------------
    wire [NUM_INPUTS - 1 : 0] request;
    wire [NUM_INPUTS - 1 : 0] valid;
    wire [NUM_INPUTS - 1 : 0] eop;
    reg  [NUM_INPUTS - 1 : 0] prev_request;
    wire [NUM_INPUTS - 1 : 0] grant;
    wire [NUM_INPUTS - 1 : 0] next_grant;
    reg  [NUM_INPUTS - 1 : 0] saved_grant;
    reg  [PAYLOAD_W - 1 : 0]  src_payload;
    wire                      last_cycle;
    reg                       packet_in_progress;
    wire                      grant_changed;
    reg                       update_grant;

    wire [PAYLOAD_W - 1 : 0]  sink0_payload;
    wire [PAYLOAD_W - 1 : 0]  sink1_payload;
    wire [PAYLOAD_W - 1 : 0]  sink2_payload;
    wire [PAYLOAD_W - 1 : 0]  sink3_payload;
    wire [PAYLOAD_W - 1 : 0]  sink4_payload;

    assign valid[0] = sink0_valid;
    assign eop[0]   = sink0_endofpacket;
    assign valid[1] = sink1_valid;
    assign eop[1]   = sink1_endofpacket;
    assign valid[2] = sink2_valid;
    assign eop[2]   = sink2_endofpacket;
    assign valid[3] = sink3_valid;
    assign eop[3]   = sink3_endofpacket;
    assign valid[4] = sink4_valid;
    assign eop[4]   = sink4_endofpacket;

    // ------------------------------------------
    // ------------------------------------------
    // Grant Logic & Updates
    // ------------------------------------------
    // ------------------------------------------
    reg [NUM_INPUTS - 1 : 0] lock;
    always @* begin
      lock[0] = sink0_data[72];
      lock[1] = sink1_data[72];
      lock[2] = sink2_data[72];
      lock[3] = sink3_data[72];
      lock[4] = sink4_data[72];
    end
    reg [NUM_INPUTS - 1 : 0] locked = '0;
    always @(posedge clk or posedge reset) begin
      if (reset) begin
        locked <= '0;
      end
      else begin
        locked <= grant & lock;
      end
    end

    assign last_cycle = src_valid & src_ready & src_endofpacket & ~(|(lock & grant));

    // ------------------------------------------
    // We're working on a packet at any time valid is high, except
    // when this is the endofpacket.
    // ------------------------------------------
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            packet_in_progress <= 1'b0;
        end
        else begin
            if (src_valid)
                packet_in_progress <= 1'b1;
            if (last_cycle)
                packet_in_progress <= 1'b0;
        end
    end

    assign grant_changed = ~packet_in_progress && !(saved_grant & valid);

    // ------------------------------------------
    // Shares
    //
    // Special case: all-equal shares _should_ be optimized into assigning a
    // constant to next_grant_share.
    // Special case: all-1's shares _should_ result in the share counter
    // being optimized away.
    // ------------------------------------------
    // Input  |  arb shares  |  counter load value
    // 0      |      8       |  6
    // 1      |      8       |  6
    // 2      |      8       |  6
    // 3      |      8       |  6
    // 4      |      8       |  6
    wire [SHARE_COUNTER_W - 1 : 0] share_0 = 3'd6;
    wire [SHARE_COUNTER_W - 1 : 0] share_1 = 3'd6;
    wire [SHARE_COUNTER_W - 1 : 0] share_2 = 3'd6;
    wire [SHARE_COUNTER_W - 1 : 0] share_3 = 3'd6;
    wire [SHARE_COUNTER_W - 1 : 0] share_4 = 3'd6;

    // ------------------------------------------
    // Choose the share value corresponding to the grant.
    // ------------------------------------------
    reg [SHARE_COUNTER_W - 1 : 0] next_grant_share;
    always @* begin
        next_grant_share =
            share_0 & { SHARE_COUNTER_W {next_grant[0]} } |
            share_1 & { SHARE_COUNTER_W {next_grant[1]} } |
            share_2 & { SHARE_COUNTER_W {next_grant[2]} } |
            share_3 & { SHARE_COUNTER_W {next_grant[3]} } |
            share_4 & { SHARE_COUNTER_W {next_grant[4]} };
    end

    // ------------------------------------------
    // Flag to indicate first packet of an arb sequence.
    // ------------------------------------------
    reg first_packet_r;
    wire first_packet = grant_changed | first_packet_r;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            first_packet_r <= 1'b0;
        end
        else begin 
            if (update_grant)
                first_packet_r <= 1'b1;
            else if (last_cycle)
                first_packet_r <= 1'b0;
            else if (grant_changed)
                first_packet_r <= 1'b1;
        end
    end

    // ------------------------------------------
    // Compute the next share-count value.
    // ------------------------------------------
    reg [SHARE_COUNTER_W - 1 : 0] p1_share_count;
    reg [SHARE_COUNTER_W - 1 : 0] share_count;
    reg share_count_zero_flag;

    always @* begin
        if (first_packet) begin
            p1_share_count = next_grant_share;
        end
        else begin
            // Update the counter, but don't decrement below 0.
            p1_share_count = share_count_zero_flag ? '0 : share_count - 1'b1;
        end
    end

    // ------------------------------------------
    // Update the share counter and share-counter=zero flag.
    // ------------------------------------------
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            share_count <= '0;
            share_count_zero_flag <= 1'b1;
        end
        else begin
            if (last_cycle) begin
                share_count <= p1_share_count;
                share_count_zero_flag <= (p1_share_count == '0);
            end
        end
    end

    // ------------------------------------------
    // For each input, maintain a final_packet signal which goes active for the
    // last packet of a full-share packet sequence.  Example: if I have 4
    // shares and I'm continuously requesting, final_packet is active in the
    // 4th packet.
    // ------------------------------------------
    reg final_packet_0;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            final_packet_0 <= 1'b0;
        end
        else begin
            if (!grant[0]) begin
                // Note: if this would have been the final packet of an
                // arbitration sequence, but the master ceases to request,
                // final_packet_i will be active for a single cycle, even
                // though i is not granted.
                final_packet_0 <= 1'b0;
            end
            else if (sink0_valid & sink0_ready & sink0_endofpacket) begin
                if (final_packet_0)
                    // At the end of the _actual_ final packet, reset the value
                    // for the next cycle - this avoids a bug where a master
                    // gains multiple arb sequences sequentially (no-one else
                    // is requesting) but its 2nd or subsequent arb sequence is
                    // cut short when another requester shows up.
                    final_packet_0 <= 1'b0;
                else
                    // The share counter will reach 0 on the next packet; flag
                    // the packet as final.
                    final_packet_0 <= p1_share_count == {SHARE_COUNTER_W {1'b0}};
            end
        end
    end
    reg final_packet_1;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            final_packet_1 <= 1'b0;
        end
        else begin
            if (!grant[1]) begin
                // Note: if this would have been the final packet of an
                // arbitration sequence, but the master ceases to request,
                // final_packet_i will be active for a single cycle, even
                // though i is not granted.
                final_packet_1 <= 1'b0;
            end
            else if (sink1_valid & sink1_ready & sink1_endofpacket) begin
                if (final_packet_1)
                    // At the end of the _actual_ final packet, reset the value
                    // for the next cycle - this avoids a bug where a master
                    // gains multiple arb sequences sequentially (no-one else
                    // is requesting) but its 2nd or subsequent arb sequence is
                    // cut short when another requester shows up.
                    final_packet_1 <= 1'b0;
                else
                    // The share counter will reach 0 on the next packet; flag
                    // the packet as final.
                    final_packet_1 <= p1_share_count == {SHARE_COUNTER_W {1'b0}};
            end
        end
    end
    reg final_packet_2;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            final_packet_2 <= 1'b0;
        end
        else begin
            if (!grant[2]) begin
                // Note: if this would have been the final packet of an
                // arbitration sequence, but the master ceases to request,
                // final_packet_i will be active for a single cycle, even
                // though i is not granted.
                final_packet_2 <= 1'b0;
            end
            else if (sink2_valid & sink2_ready & sink2_endofpacket) begin
                if (final_packet_2)
                    // At the end of the _actual_ final packet, reset the value
                    // for the next cycle - this avoids a bug where a master
                    // gains multiple arb sequences sequentially (no-one else
                    // is requesting) but its 2nd or subsequent arb sequence is
                    // cut short when another requester shows up.
                    final_packet_2 <= 1'b0;
                else
                    // The share counter will reach 0 on the next packet; flag
                    // the packet as final.
                    final_packet_2 <= p1_share_count == {SHARE_COUNTER_W {1'b0}};
            end
        end
    end
    reg final_packet_3;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            final_packet_3 <= 1'b0;
        end
        else begin
            if (!grant[3]) begin
                // Note: if this would have been the final packet of an
                // arbitration sequence, but the master ceases to request,
                // final_packet_i will be active for a single cycle, even
                // though i is not granted.
                final_packet_3 <= 1'b0;
            end
            else if (sink3_valid & sink3_ready & sink3_endofpacket) begin
                if (final_packet_3)
                    // At the end of the _actual_ final packet, reset the value
                    // for the next cycle - this avoids a bug where a master
                    // gains multiple arb sequences sequentially (no-one else
                    // is requesting) but its 2nd or subsequent arb sequence is
                    // cut short when another requester shows up.
                    final_packet_3 <= 1'b0;
                else
                    // The share counter will reach 0 on the next packet; flag
                    // the packet as final.
                    final_packet_3 <= p1_share_count == {SHARE_COUNTER_W {1'b0}};
            end
        end
    end
    reg final_packet_4;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            final_packet_4 <= 1'b0;
        end
        else begin
            if (!grant[4]) begin
                // Note: if this would have been the final packet of an
                // arbitration sequence, but the master ceases to request,
                // final_packet_i will be active for a single cycle, even
                // though i is not granted.
                final_packet_4 <= 1'b0;
            end
            else if (sink4_valid & sink4_ready & sink4_endofpacket) begin
                if (final_packet_4)
                    // At the end of the _actual_ final packet, reset the value
                    // for the next cycle - this avoids a bug where a master
                    // gains multiple arb sequences sequentially (no-one else
                    // is requesting) but its 2nd or subsequent arb sequence is
                    // cut short when another requester shows up.
                    final_packet_4 <= 1'b0;
                else
                    // The share counter will reach 0 on the next packet; flag
                    // the packet as final.
                    final_packet_4 <= p1_share_count == {SHARE_COUNTER_W {1'b0}};
            end
        end
    end

    // ------------------------------------------
    // Concatenate all final_packet signals (wire or reg) into a handy vector.
    // ------------------------------------------
    wire [NUM_INPUTS - 1 : 0] final_packet = {
        final_packet_4,
        final_packet_3,
        final_packet_2,
        final_packet_1,
        final_packet_0
    };

    // ------------------------------------------
    // Compute a "done" bit which goes active on the cycle _after_ the arb
    // winner executes the final packet of a full grant sequence.
    // ------------------------------------------
    wire p1_done = |(final_packet & grant);
    reg done;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            done <= 1'b0;
        end
        else if (last_cycle) begin
            done <= p1_done;
        end
    end

    // ------------------------------------------
    // Flag for the first cycle of packets within an 
    // arb sequence
    // ------------------------------------------
    reg first_cycle;
    always @(posedge clk, posedge reset) begin
        if (reset)
            first_cycle <= 0;
        else
            first_cycle <= last_cycle && ~p1_done;
    end


    always @* begin
        update_grant = 0;

        // ------------------------------------------
        // No arbitration pipeline, update grant whenever
        // the current arb winner has consumed all shares,
        // or all requests are low
        // ------------------------------------------
        update_grant = (last_cycle && p1_done) || (first_cycle && !valid);
    end

    wire save_grant;
    assign save_grant = 1;
    assign grant      = next_grant;

    always @(posedge clk, posedge reset) begin
        if (reset)
            saved_grant <= '0;
        else if (save_grant)
            saved_grant <= next_grant;
    end

    // ------------------------------------------
    // ------------------------------------------
    // Arbitrator
    // ------------------------------------------
    // ------------------------------------------

    // ------------------------------------------
    // Create a request vector that stays high during
    // the packet
    // ------------------------------------------
    assign request = prev_request | valid | locked;

    always @(posedge clk, posedge reset) begin
        if (reset)
            prev_request <= '0;
        else
            prev_request <= request & ~(valid & eop);
    end

    altera_merlin_arbitrator
    #(
        .NUM_REQUESTERS(NUM_INPUTS),
        .SCHEME        ("round-robin"),
        .PIPELINE      (0)
    ) arb (
        .clk                    (clk),
        .reset                  (reset),
        .request                (request),
        .grant                  (next_grant),
        .save_top_priority      (src_valid),
        .increment_top_priority (update_grant)
    );

    // ------------------------------------------
    // ------------------------------------------
    // Mux
    //
    // Implemented as a sum of products.
    // ------------------------------------------
    // ------------------------------------------

    assign sink0_ready = src_ready && grant[0];
    assign sink1_ready = src_ready && grant[1];
    assign sink2_ready = src_ready && grant[2];
    assign sink3_ready = src_ready && grant[3];
    assign sink4_ready = src_ready && grant[4];

    assign src_valid = |(grant & valid);

    always @* begin
        src_payload =
            sink0_payload & {PAYLOAD_W {grant[0]} } |
            sink1_payload & {PAYLOAD_W {grant[1]} } |
            sink2_payload & {PAYLOAD_W {grant[2]} } |
            sink3_payload & {PAYLOAD_W {grant[3]} } |
            sink4_payload & {PAYLOAD_W {grant[4]} };
    end

    // ------------------------------------------
    // Mux Payload Mapping
    // ------------------------------------------

    assign sink0_payload = {sink0_channel,sink0_data,
        sink0_startofpacket,sink0_endofpacket};
    assign sink1_payload = {sink1_channel,sink1_data,
        sink1_startofpacket,sink1_endofpacket};
    assign sink2_payload = {sink2_channel,sink2_data,
        sink2_startofpacket,sink2_endofpacket};
    assign sink3_payload = {sink3_channel,sink3_data,
        sink3_startofpacket,sink3_endofpacket};
    assign sink4_payload = {sink4_channel,sink4_data,
        sink4_startofpacket,sink4_endofpacket};

    assign {src_channel,src_data,src_startofpacket,src_endofpacket} = src_payload;

endmodule



