��/  S����3�c�ub��_NЀP���t�,ï�!U;�P{�g��Oj*�x �*�'|�N�Q]/]X	�b4)�Ob��8�O��ȸ�O_�&��*��2����K�I:[�Q�Ar���C�T&���Ͽ.W�����C�e8�<K��L�J[�(M;���B;"|�!���6?����d�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P���l̓�����y߂:���A�D捻+^N6�'�s�3�XF��[�w-��oџݷYt^����aEgX��Aa�`������u�ETfo�i�.��I$�F0�h��4�8�@+�n������"��RC�;�7P�BU$b���`��*� ���(�6ŧ��ntǧ&5�Z˥ �2��p�w[��@��}�E[��6<$`�+dHH�˙�	��E!`>�u]���\
7�~O�+���K��t�HEK���E����w_B7�Y��}61>u3� �~��.�P�E�����+�T�7�$C�ީʎ)�<cҌ���Q�����
^���gF��q�YY��l�hJ���x��*C��룞8�Ť��e�R��{���n&�RW��v/X��>h��cgot.�-�z�8kH��0�.�\g i��Z$x[�o�ڼ���+��,<�����^�QSb��[�����x��� [@ ~㚢L��W85-��"�A��]�xq����zD���|���ur��ͻ�S�&z��|�m�S9*U��V;z��T��a[f����0z�R-���_�yk�G�B,b�*�ҥ҅���W�:�iX����m��_�����ZT�����v�	(Q����?�Ǝ�lC屖2�9������mf~��^cO�zL+1�����Q�}��4���0�����Ǐ@��l���˯`���ᔪ�$�o�<c��f��	����UG�v%&��{S���~U���}�@K�"���=C�$�
I"��s7�D����@^�ahB�P.u��������0�=��Q���><\��a�-�%���|$��~�p��6�hs�ז��<_`����'c��ס���d5�%Ϟ2H.��)��F*1�3��Z�-Ô"����B��g�N'Px�>n����<�M叺0���;FەQ����S�wK�Y�f�/D�;����,�������G�Pw7{�����åƧ �q�����|�Ov,1t�_tg\�r����xs��ʨ�k�\�k6�l�˶�W�4�Si�gX��{͹h
��'p���G���	�ip`�{�x0Ι�(�z�10�>k�!��2�W�+��7��XV���KJ�ub�<� /��c6�CAd_g��?�2jR��F� K;\Vˌx�����쨸#PNM��x���fx�
T���!Jo+E�h��n"
f6G��7�� ]�R�!o�81��G�aƻ��Ĳ��z��,�^ʱ��^B,H�/l�:7��\��x��1��2���*ӷ��~��aþ�?pIi+��@�q�o�l��k�*>B?��r� ?/l0���;���}��k����_;gB|�Z��K�$�Ϭ7��HP�?=�^��I�#����pZZ����SY�AO9	�Dĳ/���(��0n��-j~��9�DOᙓP���"�.5*X못.<r� ǁ��Ht��/�K��ɕ��Y�v�"�곬,z �N��H���v�x��%���B�B6n��������a���t*S@��Bj��$�/ķ��Z�>��'<y�[�V�&; ��iA]Fa�ٗ9���"ζ��X��M����	@ �"�9�6���m�ҴF���F�y�%��ǬU��ӍÍ�>'@���g+4u�f�A�C��
��Op�n����5icr�q�K��G9�����s����RXe��+�ݏ�=����Ɲᮌ9����G2]���h]�w�*Kf�͵"n��]��qс��E����t+l� MnQJ�!����c����?z��z�|�I����c:��DX%�ѱ-:�TzՃ��#"��Ё����x�V��ߴ\�J�����k�T�u��U��g5~=0ZO���[�T�y�:��UݳPwj�0�=Fvq?6��yG?*�2[Gji�[o1y�!����$�,�I��._'M�B�|������b�.޾?��֬�i�㴮�����~����'�M=�	-_&W\l�Od�/��m������c��(�t1i��/OoC��z�)MǱ󭕡c���7�S|5]͔�����^��h��Ѵ���`�K��Z��B}�>ԅ`M���v%HY�.|�?����c5����=dk��g4M��t�ę`�8�Z*�$
)�Y`S��Ί�kZx �v#-묙�'�,	�X.=P�t^���nfI�/ؤ��Lɷ��$`��-!�k]e/(a�v��,���t bB�t����;���W�~f���E�~[�5�F��#��k~�كXS�ٝv��f��o���\쑾�/2%ܽ�<�6��[8�ɶy炋���T��1�~�&ȧ��ӎÜ��f&���%F> �Z��i{��v<ķȚ]-���B8� �!�ŕ�&����7���v���E�8p��Xg���	����5��`�����]��rļ��@���� ��֙��]!���ϊ�=��`��s2C)��;��M*
�=����
�v-����|Ҷvu�_�	@���bY1(��x�o��"��Px(h��vJ���Y��(}h����^|Z3���` ����L�&}?+b�q2oQ�]�'���L�K���.
�\"�j�#P��D4E���ʾf+�Mwj�#7�#r)��08)�6�s-	Ҫޚ������<t#J��a7 �ı����
0Ip3�^_#��R�֬�]^�k@ה�G��~���5{�C�.�9�gl�@mU��w3�H��e0	����������k�� P��l}�Ḛ��N��H�R��G��!�t;c��Q���i*u���-6���i����v���z(1'�/u�q��i��_�T��&H~T����F��̔Ӝ���!�A��g~�6�^�k�'B�3���8���y��	UC��Wj���u��� �ˌR�GtY���6O�hH�;��7�Q}�[�������y*}�k��`z���J�������K�Eb�h��Ι3�-L鿬_��ZLQ8�Wÿƽ~W�;�xO�KE=܉���SB:���S�!��-s�f���OOk��  B"m_3�[4
�|ls:�aH{��]���Q����[�}N����qҸ��x��*=䉘�hB�8�=�Ơ��Qiԓ����l@�&i�ϯ�s�3<�D�Q�`"�@��2�Ҋ�.<�6Z�זDlW����
[�p(ݼ|���5�uUVi��FW���8�Aq�/�a:��#�G��C4��R�� �'�G]�d�Yq���	Bt ^|������5��E'�T�+R����=�@����"Crf��f+�y.����̘��� �Y�m��n�|�Zt�2Z��*����i��*���b�����׌N�����S��ޠ$]��L��<)��
�0�*޽ry��y�����Ok�O	̏k�Ge�Ҏ��s���ﶞ���c -����l�˧ܞ��ʏH@Y�Z�q�~)q�����L�+k5�J�uP{�W�����q~�-�k�.�6��O�����wT���X��dB�z��y��E'��n�s�q 1���̋Zk �~���Q��ԇq1t��h�� ��������'O��V��)�Z�Kj�#)�À�U���٭�������.@�~��;�{J�^S(RR��N �WRj�EԊu9�:�r�&3q0_�u����S(`�ڑ��F��Tv�� ��`e2����Z�k�^&�|L�ɔw��Z���M�+��]���|��yޔ�cW�j�٢����>��ϰ5MA�Y}��E?�b��xD���p�M&P�Z�r�G���5���`��P��Zڪ?__�Kx���N���vB̫?,b|Q��Eu���/�3�F����kg��~}���0،�)1�v\��������#�ZW�D�AO��T��S��<
Zk0k� =�z�o�7�C�r�>���7{�*�V`�+��#d�I��jJK�yJϕX�VČ�T=��;��moз�0�� Eo��H(�~�\'��7��.f�Y����-<j�ؘ���'�?R!��f���l�D�a�a�5��i6���? �X;���	" �l-Dt$CX�Uܲ��{>�:�h����"Dx5ve�/�����f2�^�!���JU�
G�M������h�Z^Z�
D�J�<T2��9Aƽs��]�|g������]��)jB�C<��E�8ws�֑���>�5� �GWr>j�΁ �h���HWGa�F�k�I%�w!��.��l~hϧ�O��.����ȶdm)]���x��@>��!�v�^~di��3tuf��M���ME�%ɽ�Ko9��m��?��G
��\����w�Ⱗ���Q�UzX��-���ug7�GH�	7G2@�u}����0eW�����?�)jȮ�=�{��4jq��?i���	5���/��	����«�s�w��o2�P�x.Ō=���}a|�*�$*�*n'K8��l�M���8܏p��`�����(�!4B|�sv��S�,�gd@U���zZP�騡[��&�q���l�-��8�&����!6���݁�E<��Du�� ��s4�H�Ӄn�\�^GK}Z��0h���H���='>�O�+�Z��GO-��4�-��[/!y�<���_��P�^�2| Ȇʷ�0G�����z}P��d$A�W��e�bT�d\Z�Uү��S���I?�;=�>�JvPE5oŧ�u'�NGn��L���Q��'����Z_�b�V���I�d9wL��?G�J�I����ٽ��øF�]6H�x=we�h���W�,�Ŋq���B�d���e���XXi�P�v�)� ��k0�'Su���+��P�\A���]9�vv���J�MJ+�#:����j=4wuE��!�� �E�h��dn�o��=kU�T-R"�ϝ��+B1B�A���l���Ji��j_�ݟA`O�;y�n�u=$�T"q���DuA��B�U�`��g��	�.�>?��r�)���<9h�l6(�i���j9`����<�2�8���\�I��%���"\����y��r��lA�d���n��l�o�g�r�N��t�V
uuBq�8�50��[�T��J`�)N�P�Q��N4����`���02���l�^��eօ�1�i�h���N��_my���_y(�ס�w�������b�c�`Ѝx��r6�W2S���_^���]��~�e�L%gd�s.�sU)38=���z�a�V�64,<QMKoK�����	>b_5�Q,=��1�~�ǳ�����^CW^o\���F^R��W�����s��oHs�O� x�7���S�F�vH@��43*��)*�"D^�4��+��& ��Gb�
h0��L�u���S��a��ӊ���9��qc]4о�Am���K�l��#��FI��6���ɭ����7t����/a(�x����݌��_z��ڪ�ח�@�`V�2�}�dw�����[�",;�°뾃�m�fPy���m�ӊE9Z�K��h�V�;�A�5�*��CYC1ȶ5)e�.�ǢX�V)���T���{���`�۲Qe�X����p>H`E�����݃��QD+ۣ�^4_�i�fjw����%�� ѡ�ԋ�$W7~C��}Q� `7�kj�m�nE�bub��Z�g�y�wʢ����*=�����`)F�]���N�Ʒ����'�s�צ,�l��p:�%�yҬ�y��B�Fn[5��d��r���r����6?�&�.����9J�a�X�v��K���˥+�=���LxXs�2[����oy���A��)g}�"��G��D{��L�.��[����|D1ͨfN;�rL�S\�6��N�1T��	JY1L%I�\_gf��(��qI��Sr`N��<,IW~(�;V��?-)��N��M���"c�"S��c�?���d��,
�6hO�Ud�\��xb���(͟p!cy�%v���+M�-q���[��p����6�F�o�.U#A��\x���M_?�ؕ��,m^��v�ٽ_��.��	8���&nh�1ZӄͰ���|�v���&B�Az�@���y-�i0��=}O��E��UE�bͥ�+�7�ʰ�SH����}$�`�H 罹l��0��
b9�����.�ZK�{��~�+:��MMXS�����+NN�����4Kgq!�`���oֆJ�奟aXI���q	/�_�cH�#|PÑ�A��t��	@��Rq����w��=(�S�Κ�
�/4�7}P��Qj�r�HZy������GՔ8�0I�`�d���m�SR��6	�U�YI|a/����VE�T�:��%�_�"j$�� ��/C(_�|�Ysy%j��X��;�#$A�ݛ��h�H�`�l��i����7��h`�ЦT�Ď�Im���8|�%�B�r"(����Z%��p?����7S��"qh1����?9�����}=f.u��X�K<�
24~��>|�2����{;�ai�}8B��C�Y�@�x/��Ob�lB]c(A��0�N�X�cn���q���>����ه$Z�1�7 n�"p�k:%]�տ����D��j[���1V���Y��J拉� ZĠ-��rFjq��[Q���<)Rפ�`:YG����#��U���W♝A>����S�"m�9���Wa^�3�ԙ
T^�'��Gc���/�����UſPUUA vϴЏuy�X�I3��ɺQ�a��l�������T?\mk5��$��3Fc!������h���M��ӳ��[�����%��G,~��?�KV��A�-;Y���j
��'.��*�Q[�+l
�ԭfު��w�q<RA��tGE{�'��(��S�m���a���1;�U����dD����/�{�X:S��-]웏���ov=��"��D��֣\S����������x��9,���8��n\��!�?�f���5[vl�ºID;�J�
��1nS� C����C�n�M���2��N��Np 흛T���጖��S<�H��O�a�S�󺑫ssl?-�2�*��ʁ�\���O>	�)F�ؽ���{y�������r��X���aJ�7~oD�JH��<�P ��4�6:�/f��u�J�PO����{
�B�E_�m)6�@ӇUk�d������ �;�`���=��=�����(���1j�~<�� Ry�����X�r�A��S�pG��>��F��%<;lG�Q.4w�ع~f�> ʼ1���P�X�f�����Wċѫ���}wo���!�Z/���J��KM�������G!�k҇`���Oɧ��|�g��x�ܯ��m�"�u:>�]��$�, �U�>�W<���l�տ��]�u�5�:��_�Ϯ��� ������G����ߗ E�����ץ.�����,��o���}��s&�jQ����y��^�쌣u�N� �����z	�ξǜ�	H�te� R*/�:<䁋E�e��w�d
6F�aN-A�?�l�^h��.^SN˥�U�� Z�T�T��Ļ�z&v�$�{��HZ���5Ws��͙O��M���m�#|pž��o���)�pϐ�7jzJ�K���	
<O��Ê����R�uy��(�#���^��	mK����D����]'K�9��41�me��A��%����#�C���-k�~�>E�9�j�{q��KR�Ҙ?�#si�\��o�S��]���6ͭ�F�,��iE�K���So�У��ik�1�ⓗ�M�Nױ�X�����â��R��f�]�Wr��oAY��#�V���'��f$�A�ծ���ޯ��񳎢����n`0����t����jCk�����z95꣺:�܊��'�[&:�0�S�R��q̯G�H!u�𕐒4j�]�*9o0��BT$K�i��2󢊂��c ��V�N9٦gb~w�[0���{d8�����^=���YX�YӸuE�@6@R*����菆ՠMJ�197���k��(UıVM���	u���8�?�q_8jk���@E��Cp��3��R7�ӽ��<
��|g�EmU.���؄L�s<�����Ń4K�åP�J�x�xX>:6�Ń��S���q��&�b����L�c8�D!��F�2��؉Y5�ki���E���z�G~ʈ��%n�%@#~~��-��XS�f"t�
�� ���i<� �"Ƶ*cZ;�(=7�g�f�'��j�9�5���Z\��D
=V�Nq���ң��;9Co�s�Ѹˁ1��Yd�(��K馞'�O��8��y���H�y+�G��s$�m��0���2fc祰�ltu����~�Cw����y�qQK�V�^�7�V�ÌkKV�T]�8����@9�6~�a�a��z���@�#=^��C�Y���u�e�Y�ȩ��3���?�����m�[��]g�j�jĨrǜ
�Z?k����M�A=}ʿw&�Q���Sn��FWO|Z Q'��	�� 0�QF�� ur;�9��[�p.��/h�#�@��x��k�NU㧯��~��Y;?�IVt��(FR�մ-A����.���a+$��&&����1	/qn�P�����?h���E��ͣ��q<gA�k�s]Y#�wHCH5���)�X�r�t���fb�ĵ~���a���P�$0)
��(�s�,��U��X='K�%G�_o�:ԅ��$F��Jot�g��rg_X|��樉=���Ec�[ /{�W.�����(��i5�"$u���͖{1#�,Q�d�Y�W�]e:�Kh�(~�Y�2,s)O�:3@��	�~Si��%ؔ�i�}�u�2��*�wu����̑�(�T2���5bL��7G�R��A�}I�gЦ$�^�8cK�,_(�4�ܴ��G^�����]QMs>�i�h��w��Cm�쟧+눂t�!ީ��ò���uΘ�WƓ�h"�\�ƭ9~C%���曀;
D�J�L�r����<��9�x���S[٘yԖ�R3�3�&5t.>;NV��,�~���"74�QȀ���IDS4WʼS0'+��튿�����jx"�\����Ř�+�����j����`Z�!�H?@gKt��yC���{%iʗ�å+g&̐H�a|�~F �IT�x�3�M�
�{Ǭxj&��!���Ǜ.�䪆ԝ�QG�l/l��T��3Rq�-��D̅ �+'����9�4�y�ȾD��9c.�)PF	2��Tzr�)__��-�V����M���ѩs��� ��9��-_2�`�lk�\B�jr��S�v�}�l^vЀ�5F��Ղ�[�ϟ(�q��g8ڕ��V,b[t����#�)A������_��N����i�3���H��4;3�����W�8��yK��2	��l����]���ɮa�,����/�a����[|3�&�e�(�M6j��h9�jt��1/8	��z��� }H��7�y�����`>�$�w���B�UT���R�˄^�s褩���gxK�Ĕv�0�Y����IT�� �z�$��Q��I���;%}p�9<s�<������¾�-m|�PHhtC�O9Nᦘ��L�v#'�E����Ļ�_��^/S$Fy)�������9I��]�Jc]Q��C~�m��o�5�N�^mӛq�Qe�X��~f(/�E?HI	������UG�yy?�����@����	�����8��.����`W�@��A!{�f�ѧ���4���\��2o�N��~�oY�o" �kh��|{A�"z�����QI�(��~{��C�(=���}-в���i#�*�N��$8.W82�Ti3��ŭ�����~-+g��_m�s�G���-�r=`��`Zٌ8�����nr��6�j�/�^!�>ͧ4^�I&�� ��c`�MU�7�� �o�Y�*Y�_ѩIc��W��@�L�z�ƿ
Ft��ʤAr�G���.N�f}�4�i��zc��x�D`��Z���ljK���8��r�:'�Ig>a#��6�]Y6��Q��-�޷���Qrڇ��O��m�#	*=�UX�Zj�N	�r�� ��y�ƭ�����d���h�c���Y��َ�no����m$r��;8�&3tGi�srJ��bSc��,�2��v,:8>U�M��($��N����*&�]�=nz�[o��b��7`4x#W�?8M���"�)o��.�gk��o�����EŨ�̘��5�y�B��n�����5C���z3�&�Yҥ/ۻ}��U�P� �}��P�����s��V�#p��z�� @��j�Q�CB�]�^��2mݷP]g�ػ��<!�l�*。mgQW@�)LԎ�ni��XH���@(�ן�����8��O�F� !�(G�S��o�_� х�&mX�c�^=���`r{�K���g{Fh�k�[�/T���~�m��V�n P��Z�(��#���۬eeYv�GR�6�JC�1�Ո�2K��jw���)�۸eo�6��Q�hi:���Q+k�ײ�J�l�HGo���(�l�{>+�A���2үԌ�����7�|�M>�Z�Pm�6�G�	䳕��cG�F � �s��I��
dٱ8�h�{3I�<��fxN���i��-�G\w��:ܕ�X�,�͝��٢qo���]���֑5W�_�R�`��Y�T�����WF����m[��(ԩ�ZU��}�`�,k�Xb,T�&&A	� �2�0ŵ �_��>� x��T����[�̢�([�r�	���)��?��T�	E� a�  �Ħ�Ӿ�E��1՞���HnP�������r)�E��|L9�@��6Q��X��l�k���w��q�
e��ĊY�~x*������eAű���jL<�_S��m,�� N~�HE[���rL�,K*�C��8$:ozs0[�u�e�p��f�Mo8���,�b��J.M�d�Y���Z&t���*�r�*0���*Y3D��<���]�?��>�2ux$�	�,t8�-	x�]�n���M^��|Vڐ�փ��0̂�@�`h��ʐ���,�g*5�W�ݢ�R6�U�?�f�
�e�p�笊ܯc��^�v��M�՝MR���'�/�#tT�1����3j��V�x����e*Y�{0�F��Ҩ3c	��܁v������9�D��`��@Vi�g�8�G\	�l�!j�d,G�n௱�Ĉ�F�ʥ@l��]�oc�&�B��{*��j��!/)7p����d�����,��Kv�P����T��K`_s4�͒���p�h�d�Θ�'�fܥ������|��t�5�tT�)C�p@��ʋbQ�U�)�%�i� x��Fw�Th0dN����׊z��虠����h� �Ӯ^������ЩU:_p����_�Q���4"7��q�8P/%%��wF+�0�?�Hx$��@���0��hQ�r�5D��|�'H9U����`u4���nĔ8�YŇ���1ٺB������c����>@��+�V!��!���
ͤݠx4ǌ����O�?]c�]ڢG�rb�(O|=h���$��X���eOl�x".8������~�,%�>�K�9�<@�`������M'Qh�����2N��� dr��*����?ߧ����Q�=$��Vy�n��V�TCɽ��SG������꥕4`Im_�M�J/��ɨ��7��ũT������������8�s�*PI��O6W�̖x��NE2$mt�03J)5r��x<4��d�^u@.��wJ�%�Q��e|W*�;s	�� �\.�F]bE��Td�/���YCv�f��Ko�k��C�,7D��j�����.�h�sӧҺ!���{s�j✾�N�$���d�64�蚏���I�(��r��6�����= ��A��*,��F�#�=~��g��a�1�U�����3�f���L�v�w�z���0hh���yj�R]p9s(��l�D_%_p�g�y&�&$�쯉Փl��ؑ!�9�$#���"{�:`��:;jQs�-B&��xH�a�b�ޱ�e:q�_x��I�5�f}��V�|2,d�=4�9���\e��)#f�������	4g�齻$���5���]��.���;ZQe>h7�[��L9C�A"��^�M�����c�`	=����)��#Յj��4s.t�>�`S֙阂�g7���ύ� `	֮��s����-{��4��'��Y���?H&���F��b��Z�����v`�T��.���:d!*�w�x� ��w��@"�^�v����M��w&��>m5���6�ph|��k�@�o���מ�5Q�����{E`��9F���M��j���.�/���S���Fw���hQ쯺5)��cr+�)ئһnI��vԹ��J���娄���\N���<����f������ĴL�OX��	=."Tuf2����$�`�e�	b���IU�S�8XUe�S�b�� �z *�l��������Sշ���V�ҨF\��tČCh�q��v��Oo 'mv����֍t�W��j��@x���.%�* O�Ԣ�쬐L�9�W�HP�W�O-�����Ö5����y�z �J��3�o���T��\����^�]j���Z�7䗱�eW�.{i7�u{wn+��@�x�!ڤJ�*��2u0i[�Ad!To�P��?�����-!nMk���HBb'�{��f��Y2V�ʳ^[�%��RW~q�0�+�d��~�}�Q50�<s/@�'�)03��S(Q��� �0)Tl�%���أ�I}0�i���9�����.�z~�m�:ho��X�@������{����"kx]��|U�攄I�`�X�9Sex�C���Q�����!]Ү" ]�dbz�An����6��k�;��>���gi�TG�����~e{-���Ι��<��W�J��D9�q���� :ȵ�����sEF�c�9eFrĐ����s֋� ,��5t��ϧ�J��E�	v!�Д�`%�s��1�k�y�p�؇���!��{ 9���y~�nw�c>���fI���a��:.�^�Dd�¼�y��%x�1�i�<�7�v�h�&2 �7���\��n�G�7����Åg�)�OcG���ͲlD=���(!�mP� �c���Q;�a�L���;>�b�J��T~��CV�q�jJL�Ԛk+�����35A����i��<J�L��4C�>X�,/�k�2c�Ρ=�e!�׬�r��%STH�jb�WJ$��ԩk�<Ub���i3R��t�o��GWὃ�����&4
q�ɐ�m�Tv�&���� |@/p�x����%>���_;z5�H���0g��$B�8OY����p��c�O%V��Jݹ]��{�i~Tit�M�hT�@�Nev���;�Y7d��R����k�9@�>0��9��+1��7@e$?0LЋ�n�����ua�����G)�M:�ꏩ�wF/ON�<Rd	W$>74eB\ɷ�s��h�1�ȃ}o#^̓�;�k�x�	3�T�����n:C��\	 ����t#�R��7$��efz���m+Q8ݑ����Z{��M�]��j��f��$�������}t��@Ӄ�I;�8���4�!�g<|ToS��g��Q�_J����Bv�ZuCN.U��%�����~k�UT��K�Pf�Y�*�'l�9�8R��t��;���v����~�V#/��2#ƛM0����.��^����N����49j�����<˼'���WX�������a��>��)Y�LzPHWn@�pS�ﳞ��4�bf�kC-����B4UJƼ�7�0	kױ	 ��C0>��<�B;q5�gܛ���%Q��\��
��*L��6�������P��X�7�*ͧ��Fu�D���MZX��Ǹ�7��@�g�h}u����#dc<�'���>׮!4Q/,I��X'W��cӋ�$]��S�Tfj~9i���1�����8����觻��F;Bj.��ү�l�
�U�@�\�M�Z?�k����ű�2<y?�T��u�;f��%
26���(�`"΀�D?�Ii�{���:�J�G!{3�c)��6�"�>J���J���Rs+h��ɯ�A�s;N�� -Ѯ�G�	�2��k�U�!M�Z�Ӽ\1�)1]0��/���NS�K���<K�������|��U�EF�ئfddNV!�+3:	0�̨>dE5��z�΄s��.R
�+�Ȝ"_j�HQ��6�,J㭨cևV|�i�?�͟�l��֗�r���!p-ܔi*��T�����.i��nl�p` t�O��r��e{GT�;���D���_��9>�v=�Ľ ��k�t�4��t��q ����'O�.�B��BMzW��_���#���bض�n�v��� W�8�'��-*�r\�N�Zm4��ǂ�7���IQ�|Lxq�0��T������E�đ%E�ONXS\i�4 
���bC#O�ɲ�	B����\2�x&K�NU��g�g����?�͐@��a�'?���KH�?�D�rR������գ cZZ
og�\��f� ��"�8�n��e8�F3�S	�y�h|Aw}8�&#舴������8yQyYP��O��h�}�睜g��'�2Z��ǖki2;���?��m�ab���yvO��/z�v h�[�A?��<�c�}�ɒ)K�AJ�C��xB�b¢a�w�
:���l�<:"-xU�UV��8��E�e�m^�Z�$�ʆ��2�y�s�{��K	" �/3�40S
���7Z?Z������c�Y:Tn���}ը]fl���W��>�X���Bǩ����:����٣'��L>��h2���^}�,:�������^2*5_�&��P�P�4�i,lmʾ;{�'	Q�웯�T�V�`�Ʈ���F�]���4�-�t8g�Ş�b�7����[#�/�Ew�^*�U^�m���v_�uȓ~PbP�Di4Z��ÒFVg�M�]�
��>:��?�E�n8��Gw��h=p�:��2��	�������>�]Q��&/v"��^���F 
-��ob�A^�\��A���ͦʽ�&,��#�X��L2����� �p9�����!i��	%�����R��_vT�<�̿4]�2�C.���[w�`_����F��:�EW�$	��P���5��遃}�ߦ"���L4I�^h�Eq����?�����Ԕy��soX�h�>g���`AyZ�h�	��
X�*��H����S�C�=p����o�����W�>8�h<��`���`;���%&"+��o�iU�^X����
j_�bc?m?��Ѧ�W`����A��/��t�T�2��#X�j0ǔ��E�Q�A�����&d���_Sɪ����$����Q5L�n�ܸrCM4��fF�_}e�*����c�;���r�K{,3U�c�MC;j _<Qӈ���m�F/�%�.dc~CY������'t� bs$f����1��g��n�:M��F�&<DX?ȏwKX�'�Y�8SC� g�-����QZH�6��%�;�r,�+�֋[w_�(�������U���PlO{�X��<���y�+1�n8��7ŁcYD�S�?�}3����{͹!���J�4B�j�o�D;��d��s|����xL��R�ҜJN�"m3z囉�%:4�'���d'�l�����J2$����&cWY�������O21/0^��	]�l�==Xi��\pd9��m�b|�)e�Yf��)��k��8�����E���kvߜj�-J-��Z���V�wG�nr��4>�^W�'+��V�W?�M�;��z3�@}�
�OxR8�eÁŉ�`ƫ�8hA���I�L�"�Q ��XM�åW�k��C6"��j���L�!&����[/1b�����z���Oi�F�˨��p��q�-���<t�~T`�(�df����nD�����T-?�#wa�¼�����-�QV�4s' 0��I�T)u\��.�9Y�� ���B��"��8a�ރv��Rg��<���p0:�����#�|v�Q>��Xk���l��Eo��.KJgm@�f3�\��TT�4SLPړ�$(N�H^|�O��|^�����"���W=f'Mq16�W	U"o>X8��E�W��G�c��T��0W��,���(�Uw���z�b��ď�B�������EÓ��>EN xӻ'�!�Ĭ�[E��%}h*�O�0�W[30a��A0LR�M$�����Ǣ��n�cvN��a-�ӷ&����&�]˶�*DXey{m/�A+ບ�˄��e>��"_-�'x����R���\/*�u���w�g�>�������T8@ɄߦC|}�p����;�[oLS�(c)��5
�=9'��E�ǛG���"�yn2��=��ʍ�j���6��ס���sXs��DK%�{�������~P~Ӡ�Z>Nzծ�q�@�P���В�@��}����_��#�ݸ�1ӈ��/+��V��=�����;=�vC�P*~���G|�p3H�����ɑf�B�W0v4���/���^P��}5��Rܠ�s�k���`��쌡����Z�%�����Q����7�19NPm\8w��ONw����y��ynt��y����(@�u+8Gn�>�lXJ/tZ��(w������ă'z�#mq�ڝ?I~�,*�g�w���w|���/&h�q+��o�#��şbx`�
$p/�}�.�I��n|G�x�$>���_'��OfM�ִ���*���G�%���H(
�wg��c�h�F:��hT�(�����b���[�oq�_�զ�������mN����P��zhJ�6-���1q��Q�+R�NL?ts�=j�z���������#5�4�pn."�]* ���+eF��{=�������O'�.>L����FL�q��ZƱ�WA�d�rx���}��`���[�EW���H��*�E�,��{��8�䖺�u�C} 7i�N;�'O�T��Ȼ�hP��̻��O�Ԡ�U�Cޫ�C�u��}�ŤH��gT�k��,���]�����f.���cMO�#����R�5���<�ǈ��g���zMtWU�nlN����]�ok���x�Yz��m]�+��2���B�*������|J�q��L�P��UnDQr��`Qq�/T �>v�b�_��U���c���(fw���17x-j�Ω���t@(��C��d3�#�M��{�}h�>��0�ؠ?���ꝗ�䓀�cuSh��[Lty)0��"�l��?q`�8�9�Nl� �M?Ѻ������^�
,Ez+4��w���8��5�"�=�����0�f˲]i[���%}Q��ʓe�5JJ�i/b/�|*�n̹�u�CZl���ޯ`�u���zŌY��&�S]^����0�C00���њ�Y%ss��	�&� N�t`�'�����Q&XmZ+��s{����Q�eJXA�0)A��?��)�_����%n��A��������͐l�ܤ{x���?����Z1�J�"�ત�{ ^$Vy�kܾko�^�Gr���t5��i'��^K��T��C���5�&�5�tRɓ@xh;��ZOo�B��68�J�Je����]L�J�v�A
U�v�����)J�R�ȆJN^�=��xd*�s�1�*�C+F�ʚ��?�Qֶ#���f!����샿BqQ�����Ml�)"Z	}?�X��Yjc�鄞:�+/�ЗQ�U:�WB��c���}J:4S�T�̪�a�*���bh!���|h�;)O�Xg}����"3�p]�$��
͜��Mvj"�{��S�+��b�ڧ ��F�����+�Y6(II�GH�ar�T8�jp�B���o�9����S�j*�������|�u]�@ɓi�}������*����Ǖ�!�Q���<�Nu�4�iN�W8�+=FA��a"m�~Qm�
�þ��A߷�A՚fé/h���w��<�2�AW�l�tt);�+K%�+1�JS��%@��	g����+�)!�MkQD�0z�ģ����6�j	n�3L*t͗�,iI�P܆a�3�U����C�)�͋��B��+��N2��WJsީ�.:�����_���aaw�$	�d5k�~z��I߅^�F��u��"��y���ِw�+�y6t(�*�ý���/	%hn�$�$�eM�C>��9l+�ꘓ9L$��O�����j�d�;�`[�8�ۥ�u��t�K��}�=�K�_�oT�1��&����q2G�&��ￛ��|ݭ����|�vů�o�v;a?G��l m���UZN��<K2��fB�׊���GH�%��&$��mvH-���436�Mۮ�m��
})�aͲ�"���@��"D^���֙��)��`���a�K �q\��F%�Bn~�*o��|]s��}���L��<�9!����g. e��^�����1�+[�ʽ	d��7��u�UC3G� 7W���4�M��:�?_�'�x�%����},>�*����Q�D�f���#M�_������X��".C'�����q'N3*֑_����;!)�	/yv�!X��Ԑ+3)t�lR��H��0��zw87��VLm�� T5����z�֔4��>E*e�M�j�Oa��3� ����5n��2n�k�g�O%�7U�(D'�L�G��;!���'�uY& �<1�y0x��C4rTsciM��\NʽC!U0����1x�r����!��C���1 �~� �^�xҬN��ٳ��
���������~�AG��+�"�<�}熒T�����D_[2��m\��Dz�3�ƐB�r��{�?g�p^/y�`�#Q�{Ydɰ2I��}��c�� !��!'��Oh_J�_Ux�Ϫ�N�����ռ���G$[�vpҺ-�K&�+��b)�,����7�k�5���L�"�S��0�[��N�1�V��l� .,R�rޘ�D�Q�!���@�"]XrP�s�ԕ��d��6�c�L�Ν�Ѝ�}0���I܇���X�� Ev�y�ؙOi\I���2���8 ��R�ќ��p#c���S�i���ײ�Gay
R�*U�\�^�Fjn��uו�X�2�5��^FyB�fP�.��+2R�y2��)�_��OQnOk��[�'
��<m�����Ys*�����\���#��,��p]��(V��԰�$:{�Z�u�M�e��D)z�r��S�W��|mg�^0�J7��ͮ���l�=���ZCO+9b?��-�,�б�H4��M=��R�ѬEц}�U��:o��b���DcZ�K7+*1�OL�ܲ�uK�FR2������Fh&����:u��R8�e�	����n��e�X6bN��wal`�ac���M]�^y����xI�H-��
ɜ��bo%�w�O�j�V�!���յ��:c�NR'�I�th�<`�� �_c��V�k*w�#����[����lD��K�TX��ҵ�L�K��y�tɪ^7���]��%�m� ���պ2,�Ƶ�8�k�eE��K���A��!�tػ��0�g�<��!V �H��po�>�6���1�㓐��-Jj�'�R��1��;���ܷXs�(�Xf�b����-'��7��1`⏚�戻�ߥ�«�+��i�&��k�]x�gz�P����7- l౼���3|R)����K��ui���Q�}�PM��љjMR[T�w�ˢ�'��zC��T�~q �)�~=�E��3W,���ґ$)��Ҙ��H��i/��G*X�tL���q��|S�s�C�2#�v�%�2Gh��*��>�(����갎=�mX�6�ӗ��i�5�7�r���Ō=\Y����wpDe�a��g�j�m���7�U����apT���Y�+0��on/IjK�cQl:\���O��E�K$��1އ�$.�Aq?���3��/�
�(����l~�� N�Rٛ{�Kh��D
+pt�`����iu�]E�{^x�]ז��@��`a�l2����q�<�o�X!=��h�b�D����	��v��z?�Uco7�55��2�/�����a��JgtBn+-�IZĩ1jJ`��>� �n7��bXw����W	�o�Ϡݩ�i�3��J/��Q�~���n�=�P��Z��.fKs�s�ׯN񖀋w�ʏ6�w[*�s^>�k�Kw�$�=�D*C/��̴A��+��y�������	��H���>��<���tJ��8* �x�]�N�������Թ�%�� �u*eE�_�
����X�y���?�'���Qn��ZF������.�j�ˉ�m�վu����ik��4
�Y�}�B��l ?B��)�guh�bc���!j_�C$(�<q�{I)�V졺��0��3`�µ�� ��2`�㣌:����]{����e#Nn&�o�
�pf+��m���5��3���\h?�I���k��E���q�[ ]TF�?=���ܦR.�j��F��u�����P�8�bXJ���d�a����F��{�#��o��L��zD6���v�~�T����g	��u�>|"�jY�,�KԜ�ʻ6��=%�v����L�l6�Ɛsbg��=��I����!XcGɏ^�<�%��
�7�z����:�SZ����P�+j���p��ۦJ�]̧�h���w�U=�SY��LX
ńbh
���<�ն��J�L��s�3?t�p �'5.Ԟu��p|F�O��ƪ��U֧�&� D�����}�M�zd�����`��>���h\�)��e����łԬK�ŋ��t�=�#��){W�iF�tv�^Qr=��!�(�f�D�4��&�����nk'�-���"f�gBˤ5IO��ɦŹ�<�J��@���ĳ����[ ���ْ��c�Z�"c����5�-�#w��<�=���;�kJ�R_
�Ԟ7��i�H�Y���u��nd���NF���Eғ������ :�nv�6��/��G��]�$��P��x/`iI�ؤ�(�M�����K���Xr{�(��1L�̢��<xP��%���K�j�,���:}�����Q�N�޶S�-M_^i��ܸ��i@;+]W�'z���_��l	�Opl��I���u�,��Jx��
MJF�3akm� ���8s�Ӑ�X��O2\5c%�C�H��e3��(r<�c[�����~3uZR�t���:��+��D]�k�r��A?�RjB��i��yL��V] ��I�2���u��
��2��2�Hc��%�.�ѣ�A�j�Y���^C\;�4]�v񈚾��r֨�F����@0�,5Q�"�ò)$��~�E�x !��r��-�>�D��C�Q�I��!�9�3qq�wr	����� ųR�sU?�C�邇����$�$�ե] #Y��-T!/5E��w�럧�s����f��` ���AC�H��V9��< p��U�g#�v��j��ӶD���5�����q~�'l�j�o�(��G0�OM�I�C�m�1�A���P:�8�����8Vj�-p�v&\�tn�sRm�����ruL��� ���ÆBP�T �!������.��zsoHj�B>Nl���W�^���z��d�;�2�L�c�l�]�F�k��0
oZh��L���{Xs6��VF9�a��݃G/���҈^�b�]=%��y'`�ۅ(�Zj�hV���ƭE�:ܯ�U`�j";vs�� ��QH<����w��7��W~v���Bl��^�H�٤g!�}�'��G��W��cΝ��I7�����G.��, ��@�m��5�F�
3�
"��c���"7�����x�~(�����wf)_�k�K4Rh��F���8�����M*�|?%m*q�3�
F\�C����7�J�jB���I��3Q��D=��w��<��s����h7y��3&3	&���Ej����a�K�	��vM����>�3'����g5�/��/��jq}`'b� �$����;wҨ6omf/��W+�)�o���8A�f���8�dA(Rx��B^_�R(y��*���Kǻ��⍼��ۛ��&o
s��ML�u����D؎�-;a)�z�wq���;���4� Ew_I.��I�E��p*�	��b����d*���G�k��d0�6g�Y҉Z�R��W˸�h}4ǃ�������'��ՓT�:�E)��ǆb�۴C�[�F���ۅ�p���CFYo-(Tƫ�/G�O���Vo�8E��<|� 2��7��)G��۔���9_��94(�����>�)��M�����q\[uER�����X&@�JA$?i�CT��I��AO�I>�S� �e�r��T��֌��������hp1�f��5I ��b�.��eF�CfV,)ܑʠ�5��,��%��:����,�����v˙��"��wO�I�.�5��xNŅf`���e~z�n�^�:����3�j�$H,1��I�{f��rl��"�/'G��&n_�4ѴS!�ѿ��u����˳�3X���m5�+�� 
�F`�[4��\���?���]C������Jo�����l��L�T�nO�J�SA��J��DM���S R;ޖ2�7ٿ���(�mVe�[㛈'e���������C�m�">py���#L
�8 �",q$w,�l(�-0��F�i���3����E���eX�j�/Z����=��XC{��tO�u�B���Bu*��Y�T2��Y=��u��~�dR��U1�gKAm�D���4`%P 5	/Db`�Q�B3�(�"K3�6��'�GG��������F���0=���2&��x��K�ۖwO���Ͼ�]E�|�S�ȣ��(�f� �����/�S?I$���0E����D�;T��掽4�2�1gʒhd�9��� [r�)e�B�%H�W��Jm���9E��s葕~��I��#�2����Jŕ٧"��*ێp;�X�Tu�ܪ���B(�2���~s詛Yѩ��}�۽�D��T�X�0V ���|��e�;��(pP����\q�n�>%��lq�v�.����1g��W���t>��M�I� �����#��Ţ�ɨ!�KØ�t�/�:M0(R����v��A��`�Y��2In��=(��(I��i�P}�J;�D�|F�w:�NXᕪ#��E�uts`
��?�xx Jx�g1������$��MO��Z[�G=�����1��_)#4���ę���7,^>"�`�C�`,F��o�+qp���?���5���g^�C��m���#�i�$����<{�	&|N}o�4i��h?�b̂�lLn&⺕З����[G�%�b�u�pN9����P0s���ep.%=���?�+\�I��m	�"�U�
�r�1�z�g>�0�C��>��w����|>��n�d�W3t_�e�D��;K�+hl�-�~�l�DЅ���2�`�Q�f���m1R�J��@��T���i�1'hQ:�����]�R��=�rx�Jg)�-W��C%��k[���F���^N��Rj�Q]�K�i�6׉��-�<
�j\쮐��p0��x�dų�$�<��D����� )$e��2Ř��Pt���</t��r;�Z�SH���鱖#����C�d%����HHh��@��+����8B�4�ݹH�l�����C)�{����q��+���<��>����
�$-Ɇ�d,��^�����zM����O	�XR�� $�;d��`-��b�5z`V�ﺾ`�,jɍn�5�!��I2��ad��Bƃ�J��8I�5�z������،(_��&'ø5���EB�\��&w�&3U	I����Y՜�!�>a[.�c�xv��?�Y�sg�2�D�Q���4��,RAXj�N���K
YH�U+�I�f�U�0�p���X3~�&������4�#=�g&&���f�SRK)���A ���]�f��@����߬~�D���0�J���$䮽ӻpe�v;����D�^|�c�|�p�,�S�B�ن��7Ͳ�n"���H%~K��t0=����2����r�p�{0�^����D�딌��r�d��#ϡ����/��U�3ާǍ�˸:f }��k�!�mҳ̲��dk<Yz��6�ޒ�F*����S{wr�u��5^���-� )# ���]~�p%2�w�b�~0%����qz���:�y$3����5<���E��E��cbp+)��Ұ)�t�H7qz��� �	�(-4gX	�c%	j�#2�ø
�}U�\�V9[Mq(�P!x-��G+�1��(�ăY9�U������x��>�Hڠ̶Q��9"QsAf41D��
�"�a�a�v�fD\R�;�ӱc�"mo��%~u�c=�Z��C+���]}?g!2��`��nl^8�
�ћ��ַt�eJS��E,v����6��3A�����o4�U�#�͉r��5���ڽb�r6��r��ax�s�|/d_ ������c�u���W3���j�ti��7��2��R�V�E��$�������Ll�>M��iCj\��W�Cj�����5pǂK�F2����0U@�V(r��&d��KY��ֵv�c��O���`)ʰ�� #?�z���|�Pz���?��C;̟�­R�.��K���S����s������K����9�%��y�õ��[��v�k4v�3ASWFzifͰ��H����]��jN����*w~�%��JX�w�Q֩�`k���R�+���d�w����d��D��������eтV�/_�粒(4�����L�a�D��Q	J� ��)����*�eҗsN�Ѣy�FțE%���x�x�0.� ��0�*m,��H�W{����y]Sz�uǏЄ�|���Jd5q�ڻ����Y
gE�Z����Vܱh-�}���j�����|>Rא�U�F��))�"!d
�W0�"ZJ�>����o挩F���
$@�������*�<��d�����`�=#�D�2���������]�]���*./��cK�3g2G���?�6�P�Z(w��dEN�>,I39�B�\�Ϊ��c�`��?�����n�g�793w�wP�Yg���dY	�\Nɔ7-�1�wi��W4�А��9Bn1�fu�XD��p)moaqrw�����yp7(�w���G�V�I9r$2���֐Tt�@�^2��Myu�S� ��:�7���ɲ����a��X��&��<�e4�����'���E5%n-�j%�q�&�l����Q�k���%� +�:}�?���s��I��B�<��o�ȱ�O����J���?��H8��V��JW�٧��5á�TjI�����%�MZ/��s�A��X��ξ�w\T�S^�$om�SM��c�۰�K�{�S�TI�B\�lJo���˿�FSwd���� x��V����\*����~g�b�S4G�A�L���GQy_rM)�@Mf��#�N���9��-��V��t�k���q�f��"���|���1/m�~>��#}6����EP��<��i�����K��y[�4s��Tb�<ܺfa�(=��G�zܢZ����,,"����y%m+# �N�K����K��n���7�v`7��*�Hlֆ:�9��7�eDC�nH����`�{)��v��fo�T�qek�y�v�4�f�>|�[As(�X�`�h4�ӳ�>�W�x͟pH�V0�T��m`�iH&w��NL��=���4�O� P��o�c��v2��	��N������X�B���-9��ɗW��t�O�G
�B����2��1SB�	u)e�����@7�� ��H����r���IT�M���J��;|���}����vmh@��<Ąd��ц��^�9��c�
��g}�_��X�ZbR��Q(��ٵ*�mw�n�AՎE��9���O���u'�SlJ�'�f'�Q�/���\&�u��]�\X��tG��bzm���[ڳ&��5#u�[�є�E�(FTt��w^�:*��,�"�hkr��W}�io�5���Fi�+}�Ƶ#;���蓧ftU�H�����y����U4'�j�����/+
�irg��t{�k:eD*�U?EP2C�Nv�N�A���8�ŋ�\H�GW�c��~�xXU8����of/�X�q��3�_$�'�Py��s�
a�R*�j�{&>rS%H�4M�}f�n�MJGg��5>0,m�t=z/a�!�a���O�K�-z�{��X���s7_�J��k���>�]��Q^R���_|D������HЃ=����f�j�W|����}�Tu��#=�ɵ	(�'�'g\�5�J�s߼-ȳ��_H��*q$�$�DRS��E)���M�&�Z0:�	1��hV};	�,�����v�h�tA�D��w�����k�MJw{�Pt��g$��r�d��g�ӽ�_HNߎ�	7�˝|�Ɏ�6^�a4�Ɵ�u��fZ.�G���ih.å�R����-���X� =��]���Z�3�}����w�����k��y��(#K��YkW��sYhN=[�rOZ����|�P��`vt����4B�� �6>��ꎔS�*c��?�xAZɫ5$sl�����0���2��V#7�����G��m�̰�2"���U%i>��S���b�l�p��>��՞�+i#T�0!¤b��t
�6(��^n��b5�����Hq�ĥ�u	u���%��\���o�d�M�m�@���ފ��z�o��b�X*����*]K/K��1 =/���7(Oy��Zo'M����ɨ,A���c5���HrS�k+��]l;��HI����v�$T}���:���R\�k��	�^�A���^�nkKs���m��Y'����+�`���^8N��?E�֩&�I�W����TÔ��<ì��)�9d?��s�_��8<�P5&��T���~������c>%9���bQE2	˚��2&���>\����!걱���3;��4ϖ��C�Pݰ���EyH=�/Ƀ��D���SĜsA���dn�v����Ŗ̏%ym��P8f�&����4'�Z@%$��:�����A@8��/1�������_����C�S/�ja`��x�<A$Ґ�'�q��M�"+�6ؼHk�R�a�l�zu�A��߽�z�5z\�Q��ĺG[��vw��An��~xֹ����Qoe�t�8
B��哸�=ʥ�^�酳�ږf�y��$0��LTv�:�S`�W�L�'S�t�YMB�R�� �����犰���*q\��5t�9NB�'�_ҥ�˃��<x�⏥�t��(�#Od��B�>->�Q������@���^�T^�{�]��p�'%PW�w^�B{�M?4��E�K�ޣ�&/��IŗJ�սY[c�Ql�G�i8~m�����V�:~����ա���"b��Ѱ�ҔA'��m�$�U�� Ո:ډ8�F�k�bI�d��nZ^���5���_�,-��^
I&�\5��׽2kQY?���zU�\�**a]y2�_�����nx\t���!b'��� ���W��^�x[�F�i<a>Q;�2�n�S���H��T=p�����12�T�R8Z�W��&l���PT��+��s���#/[;�񶓈�Z���\v��1_?�{�Uv���Q�9B�|���*}�
�/�ۢ�+'�>����ḓ$�性P_M�V���\^$���:��T�
���Q�Du��H��9:�b�Ҕ� ZQ[M眵��h9��+������aO쑟�I6���Ï�:c�q�8�2�{B�촹o��c~�c�e!�%���,Ee�����?z m(��&��S��N�a�P,E�V.�MX\#��g'gd�>�#SQ���8����_�y�m:9��(�Z��(���l�G��
|���v� -1k�#u@�����~�'q����u�$L1��M.�s��est�J�#5Z���6��tA�kI�D�ަŤ9�F��ux���wl!new�)�^ZWx�<A(��Ȩ���HA7�s�e�����.�ܸ/�h%���󩞛��ѳ�l\�3����[�������x�3*��M!���.kO���P$�7)0*�I�nXD/���;8J,c}�J�;���\�>�� T��.ʾ��tz!1�`����D�%�z	m���	�5S��J-P��d�s�S^H��p���u���F��ٯn�3B��*�!P_�#;��Ť���o��Ѧ4�zFgW�������.�x6~(	��Ӯ���HT��烙s���ܿ�?mr�+�H��	Ur1u�XL�F-��{�j�3��x��KYt�~�	9��D���=���;/��s��,-��M�����fH��T]�܁=�עcv[_��j���U�3�pu�8�FO��^�j.wzVI�&W��W��e%mse�Ӭ,s1�� �s]TسK~
�uLПd+T/�J��5��+U��8s,���E�����7Y /�jx�$]١E�5[&4��O�S������V�$�Paa�x��q��V���ϜZOfl�I1U:�᭩9D�`����/3�M�{���21b�����ɍ��ln�-z����l���cVRÆ42�2�@6C��(*�5O���!j�徒��{^h3��L�㮗��v&�l4��-�d���K�-���OT1G��Hp�_��ʐ��F2�ш$x�&LU\r�I#�j���\l�S��^�&�N%1s����'.W� �^M�cUUY:(Y�l��ޯL�1,jŘ�"q��I�C,�M�M�TvWd����B����us�硕N��@��z
�*��|�hlI��� &��1��gpk���p1�4����9�s����Q���֨r{R'�f!��7�w/Mڛ�L(D?��K��=���R��R�:� �&�#��\�2W��p���<D(k��^D�<�9k��c���Hܼ�oh��3H�"^؀0�Ptjs(�i*w/�*�4@���{.l)K,��9�������T@���9\�������x�ģ��ï�f`��[.���@p]U�Ģ���e*b��a�~
p {bP��cXt2x�ًBA�C[YYЂ �1mi���%���8P��ژ�W�Ÿ�NHw�fKM��Q��|��vio�MC��J�\Z'ݖ�ڲ����4���+;������:(���HLp���	m����d��v9�L	�|�%>۽���/ލ���?��Q"t���������ĭJi�w���*���	�oC��C�1��Ɍ!�qp\��k�JE����q#�"U#��Q��#��6kj��l1J�b��\1X�����Ύ֨+������Hv���*��r-~r��ix0k�Sj�b@6:_K�_0�.�t�:)����F�B������^��&#(�`0���xʓw%Y
g�`â2�T�P�r�BBI���&JI��9�9H_�TM��P
�)N;ѓ�W����-%���oќ~8y=V��+�Q�Q��:;�X��l'wҫ)1��jS8����4f+Y�|B2!�����3�jm��mE�vL�1bʧi@� ���L,�kΰ�d��;�R<���`�O�&�&��W�5\MCz�A7�E7�l���W�����F)oE��d�I�fk�O�8�/j �mʲ+&���?'T�hnH6�:���l��ߥ!c�8+�jDk���F��t�۱�E�9�N�<E��L��{�8wr]7#���h,���F7�V
 ����p�Q-U�R��IRpF��8������v}�Rr�r��~!N��2=f'����]�/���-V���a�ѱ*��a�u��-Z��_T��6=#ǘpN�����+�����B
tapḑ ,X<��6[�������N�,Ulxd��ݧ�t������-�3fT%�n@nYz�y��j8B�:ax�ש`(\��0x��9�1J��*D�ߘ�i�h��Q5?�v�H�d�7N��i2�o��4��;2�`�`�1z���C7#q�7}9���X����V�2H���Y�S���0���N��P�5@����p�ӛ���9��U˖�c�X���l���tSi�� �U�ih��[����)-�	��Đ���r4���o�?Qc.�!�&�����E�k��B��=ե~�eٿ�u^?ѽPF�ϫ��t���S��1l�5N��+���<�O������𯴭��)aE�P]��g��x=4L�߮uCH�w��i�e���0����F�pd����j�t݀ўU�x"yQ��(3������&�4�K��TL8���j���C'��$t6�߁ȪJ,�T+��0�ڻE@�irNz��6ٛo
�����D���xFkl�����{;��r�Z�4��'�||Z�'łƒ�X6>����M�����z��'�����@KV���N:!ܾ�s�ӛ���d�+�˃���Xݼm � �������*��� �@YnM�z���9Q1�S�m���b���{1=,���~l��D$�q	g��
4�<�3Ԓ�����/�B}�-��t�656��7�"u�"�S����\�$�^�`�x�J\:o[�s�х:ڷ�0�H ��ۋ��}���yB��\n��?���-ɘ����4Z��=��mxfkۺ��eu��W�-�i��/Z�_A���=�,�����]o�dU,Ԗ�0���/Ք�ij��0!\Xh~3ō7<��a�^�-?�sI H>I�^.�>�8c�	ɬ��ѿ�h���	�����}�k;F@�$�1<)�sse�RS2��R^�;$�Wl�v-U����I� �7[���Ug(�������uoT_K�wS<gd��es��2IE��3	�8��\C3	ۖN�Q�]tz��k��$C�f�>�'�B{��D��ݞ���v�6m�FuY���x�/B�:)𴅞E�tiٿ��g^�o��߳���=���b�哌�o��/_�;1�gk�4j����"�cI*���*�t���s��	�\�X��ዤ�Ok�o�
��������!R�o+lh��85�����M���������V�ҨD�jV��-z��j�8on�D2�����u2Q$��_b�1v ��9$�����k�z^=~��G��8s��tJ �>�����J�X"��Fv���=7z=�t��":�����זt���@�ZKF�t���V1I�Ę@J'�d�t�Ë�sE]��`�r��_�*p��ʇ������S�a��kwIV�r�?F���[d�&�mb*�S��+�Tc Ѓ�G[��~]ȑ�&ɤwn�xS�9�yɞ��W@ѧ��"�eΏF�ڦǾ�t����A�o���ߚ�4�2 �G����3�����c�{�F!a�(-/����jP9kwL��N��р;�^�@r�����d�I�-#ã�ݱ�K@��Yl���u�-6=�a�Ѐtu�c���y��u�[f-�4/Od�M�T&L��D�@�<��H4����XãY675�$Lp�3�����Ό�Ԡ��ּ�X���$RU�5F�-��U���z���y������,��k �s�yG�9�[wJ��`��nl�)��*p�r4��|�׳m-�� �M�Ϸ�h^��c��&dހ����:��ܔ�vc�FOj�o}�pp+�^C�{�#o	QbT��ǭم���c����@���f���� �W��\�ٕ�@����Q%z.�5��o NJ��jӈ�sJ
lAV	TI���C���J��zmd�n���	�b�gnRG�8F}��s��
$��K�}��
��e��qA`�: �b��<�{5�x����x���車ȫؤ�f���J�4?���,�(�j
>6���B��Sӽ���MC�N>"����|j�;����d�tM�@���ʅ^�Jq=N���V�٩�^w)ݍ%�x���r�5�|8�� ���a��1��k{I0!=k��4���/΄,F��x�^~�� A��r/�����D�������ш��0�_f-Z*i{��t���o}���rZG⁾;��<��t��b{	Ϡ�<�e�Xj8�SSsq��1��:�=#'/���ŊD[�KP�M�:6M�|�?���.@�YF�U��"'���t��d���:j�}o�T�+�V]	fG��b����4=o�PC��v�2d�a��{9��TeW�VA�Ņl��8�R~��u��{`����%��yĦ����]����`�v�!lVT��W���Ae�����މ�_V����A�1`������y�h��^H�Z�^G�]ދ�
��ؾ�`�ا���9%�#٤�	�~\��E���Nwb��I^u��t��7�0�l�!r��¤3|}�x��*M�[n�@:_�a�������KM�pI�\2āU��T�A:��g�f�Է6"����y	�BU(&��.�"��s�Q��^]t��n�f����z+�Qі��<�>�oXAm��v��۞�e���M�x�G�`eYu�� 1���n����V9�!�%V��T)��4?G�v��s��zL�B�=R%�=�D�	ZM����hi믷"�֢g�j�ȭ
�a&'��/���	Y}���>q%I�m%| A0�0w�d{�!�U���
���o���r�$p��!<���_�b@b'�`�E�E �Wr��c��8n�#S'j�� ����l����m����Ki�]/9C-I�2�٩Zy=�J_��(���>hn�L�[��Q�ϫ%$D���(��Xq�3�bm�
t�BqC��'�+{䨨.d��]�C�xf�*��˦�v�`m���9���2�P5Rۅ�J�1O`��tU��B�ؙ�rS�#�	Ek�Dd?��8˙ރ����,����P�;}j��}�B���ٹ1ע�2ן��%ӡ;���m2@q�u��*"��Qʃ�Ėbt8�1r�b�ز�A��c&�hPŖ�RV��1\����t��S1`��c�T������s��)Z
�6�0�T�5��}M&Ph�.��_oj���]��f�p��	��ba?���3&*f���q�ƁUG��*��j�;��-+5uf�{vɢ/��{q������!*F�3g�_�/+I�h��y��<-����V�������B���^M�'[܃�Sufd�`! *`xq|�4�*�]�cB(x�&vOW� Y�����-�Ή3q)j ��d4�l*����P������.Џ��#So�E\��ߩ���!I����J�<gЃ�"^{#�;�G~�(�_��䬭5��KBe����d�jt�#��{�/9�����W=Vt�} ���j�oq�ى[!J}�}Q��eP]���&H���om@������麾�F�E������2�'	�JJQ��bN�$Î� א4�]��:��H�����'��㡧_~� ;~�'.�v��R%��Д��m��gIm~�*Y`v����Z�ezNҝ82M���<��c����Y��l�i�9�!�z���Wפy|��}��`�5�n�)��y��&��ZU�>�g�(�Js�r2��^�-jS��gyBW���38�@��H��7;���Gvu���"�A킪�Qꔴq#���.:p��e�P#f��v�nCײ�\�@4��e�.����r�Z?��=j�O��l�LY���M�Y�����I�X�40�%Ix;k����~*�0JՎv�M����ä%t
��-���έՓ�#���@��we�-Omwdt�B��Qͮ{z�+�374�1���L��HLŚ���l�xH ?ׁc�GA���� '1��U"���R�=�%E�N�E��	r��S�����~Q6K����)H�I��"�T� �:�43��B�j����H�bQ�ErTT�`$��F4�4$g6�0P�T*=�+����>�c���#P����ڜ��%��qݬ�R�d��YQ��?r�:W�D�"F
���\Z����D5En�����?�^F�h�9Љ��������RV~��oU��?�n+�����Rc�Ԙ�O&��!+= x@��%��/Wz�ٰ�L��9���ZȆ���܆1k�F4ҟ�
c:XU>YFF��If���¼��3@��̎�'�`/�gL��.�ٶ-^����!�e1��7�/\M����^>l������n��W��ߩxM�a�s��ć2	�ΰ���i��P���0=�a�Iă�sĶNiDk^(f��Ϋ�'ڔ��
��Fb�i�B�=OF�{~���pU:�����:(St�����b��a塂;l��S��� ������=+σ3Z
�16�_��Ih�0{�_�Iу��M+T�k~AR񂭎��"�`c޾�� N�W��;�܇wt>�k9 �3���M���z~ie]����g[$��
0�����^�MO겨T�֛�́;�,z��:�e�Vn�P;?X��/��Q�J�@��i*� Rl\P�%Ѐ�p�̗@2:�⧳�w�`N����q��l�1�׫W�y29tFy�7�Ž.�ӂ���B�a�d�+.��J�OH]�����U�NJ�L�)sp�
Za�)_��ޅcK�&����l����;����3�B@�"k3u���Ae:��?3>�q�}�I����A	%��y�&޶�!�Do�r��(8p?��e�����S��}�q͊q��鸓n��� i�L��2�f�Y�%z�g��Z@O��=Zi��EN1e�V+z\�
vCw[ֈ�	���ҡ����a��cSI��o'W�z��W����~�����+��$�C�㶋��0T����ܽSDA���~��?�+�>�q�g���M^�D��0�}�+1 ���>2ђ�Uu����4�41���5��ܶ�wĈ~+��KA(v�ԉq�	�ע�i�@�g[�Y����ޖ*��ő9&��,����ؽ��D��z���&p��M��B	ʉ����cux���=8?~?��Uۈ���cڮ�v[��h7�Թ) ��h�Xw`�y� �أ�����l���z����8|%.V�g�ػQ)�(͡�+;ɒ!67�W��F1F+���-��r\�Z�a�0���G��)�Ӡy|\=�_Lp�- ��yz�� ?.؈dp�0z7Ր�+k��x5�!�y�\A���3J�q위�N�[^u���s�"�+�u�E����VP��H�kk�4�������i����ӥ�KPg������0_^
pq��?�M:����W�*��K'���>�C!E��E��Eڭ4��2�A~L���ȉY4;����G5ᒦ�_*'��=ႉ�ހ%�yi���'�N�G�v� n/|~�C���o����:��G�����]�]���
��j���t�7�z����|�n�-Br����U�#� z��c��Y���QoP=�П�6r��#�͐�+�l�WEy��֌u���5ό��\(RP�����&9د(8�'�B$�)�B�`�:dSp[�*o�����i�;�QV�9�'a0�������R���q��������e ,��<�JQ��I;M�64���X��uA#��P� ���v����A���g��3R��QF�������OJ\r�kN�PE[�v�b�e��bK���(-0�I�KwZc9��E7��g��-�D4���t#�V*�L�_�����4nj�u�4�h�{�	�ߏ��kq��;���m�~ʐ����Lx/9����"�-O�C�H��,uJ\��>�e� �凬P�)`.b��n����L���E�jj�縉N zh�[`�ku�&CetL��s�:�k���4�M���J��2>՞W��
�Q��2g�:gʜZMQ��8���<�%"�r�z���G+,��LD%g�skU�i;y�32�BMw;�W>��}�6�����-j]ɸ?��V�{[uY�ѣ��b�PQ�s�����ZS�ή>��Wu�s^���ӰP>��V���]z
:0��n
��*�/��I���i��WGD¾=J��M�(Q�Um�P��؟�(��b��<�&U�$`��Y'��V��f�-E�"�4=Qf]�\X���Y��y���P�M��h�Q�ʻ���ɑO� >�*�:l^��W�|��z�=
Ν�:*�a�8����1aB��ں��|�q�k3r��{�ہr���uw������Ȯ�{�(.��.T�6�&,|C�૸yC���-�L\jV�\��17a�6-��sl<4(�R*B �0���hd�ͤA��\ȣ� ^����υ�<�Vr!��:U	�uD�����L��� .͘��.��n�ݳ?6�Sn��&��j�מb4G&���]M�؃k��q�{���*
͒7�US��q�Se�3�'�*�
��G,��[>�C4)�����|�}��"ë8��4I��hS�"R ��w�.�8�����?�L���%���A�F:F�1��zHފ�
?{hc|T7b�"�~�Z��d46Б؎�lb���-)��#�YD ����GO]�wW�\�+���B;��?sR� 8Ev�fHA|q@�t|�%����`��p���7���8L�%Ab�b��Ycl@3C9�PD���`f�j��˶���&�8��.���c4�Yj��*i���+�g6 e�旍{�A	m\��;@pWw��-�1 �'� d�IZ~���j���Ç�o���%�����<���KCN�����dQş�n��5�
r��R���-�u"�x��6���/y��L�ᾟúG�.5r��f�۰ٻf*������¥���AcL�{�*rx�%�̬��_'��C��P J�ں\ƫ}��M���Q"�tt��
C�����LL��aַ��X����i	u+k3z슼_:oJ+�}�a흮@�2�U��;C6�JV	������2�L۠�h{����M�3� �lL��	��F<P��L����^$��\F�������gb�K��J1'{��h����@�P����O� t,����18�� q!�Vg����A�3USÕ}��z��?Rp���n���[�:��
��9����(7�F�Գµ�;��<�P�v,<������}����H\T�
|^�dZ#��;��2��@��v�}a�`�hh���UI6�.��lS��$+G�3�|i��a���� {�#�b�����+�&[���rxMt��%� X5���Y�,|v}ާۅ	Y�B�E����LVW5�c�l�3�C�$AOGxP)b��T�.}�����jG�#�60y��v����K<c��$�5��Pa�у�cNmVs��4�p���4/#�Di��Ozs#H̏H�ͫ��J硉�5�zn�)S���9j`��@�T���1�)&�G�/ď�a�&?y�,���3�Ha�Y� �L���eY��䙇����?"�^ 4�\�o��v�Cby�0��s�B](�u�,A���@�ы�'"�t�����O��|��}n�=�����fa�-�Q7=\���^O�aq �&Xv�
)	��ǵ��r�p�CB0XߟUB(�*>�ӝS6n��^�g���[�Y��4Y�'Zb�TM?��q�aL�[�~#z����臚$��b���VwM٠*D\�ȊB-�OO M����w.�(�!��Y��,��Olfv�F.�,)<�k2�F�Z���I�,�Q4@��G9�=�Ɛ`�w��->�K����O�EIO�Hm[��Y+vq�P�i�-d��䭤����F:��!ؕ4<
�W'�J[�t�:{�7H#z���S%^+R�/o�@{  9:P'��}�b��ڳ�{�l9�p�[�
fe���9�(g��]<��e�T�$Y�M��ǂ�=��N�8�Ӣ��Cu�\�}N'R���Ld��!���@n�cZ���:���0��UܒUA�jI����2��()Zj�3���\7��<M{�d�*¹� ���,���|N�=��-�%�N/�G���/5h����θc�~�t�UYX�����&�-���D����2ĝ]3��q6��lF��J��Ħ=�j�z��T��B�@��j��$�i����On(�c��r3l����f$�����
�l���_nA��oW����H�M�^������E�}�� �D.~sM�gw�ڧ5	.^z�~[�ǒ`��zS�� X�uJ��R�fz�q�A[�}��#uQ�W�LYJO�l#�c!(u]T#&na��AE��Tr�7��u`���l�m�H�;��:��caJ�<:|RW؉��/�?���R�!k'L,S�UU)��pd~˨�R����m� ��C|��.S�v��$�G�(��DV�?�Ap�/tԦ:��׏���}*_���G6M�Q�I4|n�x3��'EV2H�$P*��������O���sF��Jx��7ȵ��%(F����,[�q���A��u��'���r�����q(�#;�ܹ�������A���s[b�A-g����i�W��O j����û�@쬽:�$����|���G�u�u�l���������w�d,J6`��Y��j�Q�9�-�K��M[�� �Q\∭@�x�_Z��@��ԓ�Vr����3�?�q��ش��?���H���PE��Q�]�ק+��}kbT�t(rF����E��ŵ�p�k��]�ݰ;~ų�&�8���I�7b���pXER���o2f).�d�	�D�gF�v4B���Gޫ��8 �a�0I���J��D�{��z�;W^m��_(�z��6���N���-?� T �ݻ�c�QR�#�B/��ќ��^���0����r�C┚�\~�+D���|)r6�Kȅ����Ǎ71Q)��߭��f-�H���i% Łk�ʭ�OZ�t��ٝ9������M�t�	�^흄^Q������F��� �����!��_�B���wA�¿Ң�q�'��Sj���п�yV�k���r}���j"^%��S�и�`�����?�-���7a|G4�Ԓ�@�1��~�W�}xc:�)7e�j�N�XkPj�.M���I��($�z������}�fw��^����B��S4B8��T��*B�V�l����N,�Y� ���}3���1�Bfz����\��h˪�Y3�1Nr1�'7FH*�a౰���V��n���m�X ��qI���n�a����;&n�s����/���J����??�qd@��K�� ���c�.�.�6w[`�:y�Od�Gg��[A��d�˯;�vK�����.����[\�4��I�&L?`����)S��^:y�m�4�z�sXN�"��jF������vo�7��{9��Y5��b�Rg���Z��J�{{+5����Z��?�"���oV�m�u��d(J��l�8�Ւl�[��f�6�^遶^s����z�Lm�#p�&��Fܝ��ݒ�m�Z�Q�&aS�x��M�y:�I�ʃ �o^��l�]��3C��A�dP}��W�������t��Aj8�<f�+�E����x��%v#���ǭw!�ۿր}�Q���@4����%�gwr�%=-��A,07VO k�~��L�#nkć����@�mq�I�y_������;�T �>Q��I��9�b���m<�;�̶��85`-0��Zk�=�����n��<���|�=�W9��� zŹNJC�����q�H�!{�L�
m�Bvb�_k�b�Q�>�N	���r(z\P\����ʇ�d"�oɂMf�,�ma֩2'@OS58&ÞѼ3iAѭ#�
{V�W��rj�_�g�y_!��������cqv�l��!����!OB��rz���澟�Y 6{¢�H��`;ꍬ��j��u僿��̓�z�	��X0�p��1���O�������Ov�'�m�[�V#/�ˠ���x����0YJ(F;��x��l<\w�rx�uL+�5S�q�CZ�҉��������*s*�x=M�
+y}ŀ�)����p3�0��.�pb��%X�Pl�E��Q�X�v�tɉ�e��|J!1��D��L�����	��'x��!Qf]���j�%b�"����R;<�
�.��P%zV�T[�����:Tˣ�`]7���P�kI�T��s�;F�U{6VIe@D!�'��?>��r��y`�S1̈́]R�etun��?��3�C�c�ic��;����yʗ�ӴV�^��h7j���8L��\�P����ǲ)�V�X�,�<�!��������੻k�#8`�֤������WbQ�4�F�^<�N&��G�x��v��Lc��j���1i&�Fo�w� A	�UJ~�2-�G�X]O�JB4{�(���DL��kN�.%����;�5�ׄ��f"���"�Xvz��x��oWm�GS,~dz5q�K/)OmSM�����x�[��xЗ�� 3[�I�\CKJ���z���S:i�;�گ�(+�����������C��[�qW�YNCM��H��=�?�<@�����YZc\&;mn�2t��SAp:P��������@�Ց-��R��Ovi�R�q'�"d��x_�x�����D.;�LK1|,��f�B��Y޾�Y�O�+����]oFLK[�0��|�p��������¦˗i�I.�n=�a�//���jL��v���A�S��V�]9ڤ���.;�S���(0a��4A�x{L��]9Ƃ+���>�L��2���GЎ�����Y2�x��*�Z�3-�7L�9CM�T%�4�ˍ/�G�M,��έX����"o�:g��o�9?w�8��X��������Fh9�c��BK͸7���#�Ü2~nh���9`��0����t���p��#�tɽ�a5�W���ȉMñJ<>�P`D���ğ�o�ǈ6W8���Jp�����1�[>�w�ƺJS���� ��%~�]�Lő6����)5�����,�#c]�N+��P�=�4�<�w���.7e5��n�3�g�Tu�l�xw�6M�%�H:�@�ݛ��Xم��&gqRx{�U��MѨ��;5��4`�~?���9�7~A��I���'��$�(B��R���6�<u��V"k�cC��;��_Yz>83�Ks�2�f<֑W�m��Ƴ�Gk��[=X��!��U��Ӌ�����\�_v�PT�����K|��2iN*����]�����-ɬ�b��8���nꢍ�9�B�7�vz�^5�,Q=�>��4g�(�0m331��nE�5����9�;�c��Y��
��o,P�9"+?B��~��p��Ux[%u�����L�t�g.�c�=��}h�u����e�9���*y:|�� 2(�Թ�n���P�o����Nc�s@����P�~�I����VF̒�khE]�)�'�\쪡/U���"?�"��e��Ш����:�0|bm�A&����r�"@`��:���y^9��;�� �	�I�P���'�Yʯ:��o�0#��M�'me	}A�4�B�!���	�6_1K��qr��BoV�K�jȉV�<n������Q�Ulj��ڢE)��]<'g�7�hn��J�{=
r���$�B���BAY��M�Ǉ	nP%H@;�LTq[j��ľ���8&���*��'pn؃���B���Z�ǜ4��Qk�jAi;N~�!-�rk�b[����M4=��j~k�����ȣd��f�͕h��ރ��&1ǿy )�h��?y��Em�g�����a��d�?>��T=<���5��]�(��'�0�	\}�q���:��!b -�7���=�a(��b�߇��i�/���aI����gҍ��h��]���cBÇ�;��QC��K���������I�:z_R��G��^��?9V_�;C P����<�$��'=|�IY[�s�`��_����W��y��_�܊�D^�Ԋ�p�i�ř��y	D�;�%Lu�OHl�⹊g������IX�����n&?7ȧS�=x��V43� �7I�[�!XsL��~��0֭f�`甠nl͑'��9�KL���yo��G�,�{|�'(�Y\#�<H�A�=b�Oi<�1sj�x~���8��Ė�C�3`H»�����ܡ�B�̶Q�)���e23�oVΒ;Gz�1�/:�
���d�Gv�|M5B��޵���E,���/�:�C������\L�:L�԰넧��L�����
r�?g�E�6t���ԓ\׾G8������n������t�(��-o�qQ�&Z�}��2
$�Ո�@H�;+3����h�� ������-��6�}�d��$���xbws�c,hK�=��<P���(-��K�V�N��̻��Qˀm/��� A+1�~�&Oy�tw��-���v|	`�/25��f�wڜ���=�l*�������`���rۡ�n��ͦ����xLW�xv}����Ȉ�֦��1ة`�D��2#nu��@f�����K�L��Q�o_MǍ��X~ټ��T	���+�gƼ��1E>@sU�"��f�r�#��۞,��];7Hĭ���{��_Q>�=�[�2�\�j��4�M�?$�%�7Y�0����:��=8C]�~T����Si���@�0�C�I��˅��-N��]�Ȫ�w�}��)�U[ޛb���]�C�gn��~�k�R��/�y]���^aH'-������19!~
*/����w�h�NnPV���KLֳ��y!ʇ7��B�a��L�������-�3��$Q�&r˻�@�BЗ�9���
�r��6gG��T�J��Eˑ���Ƨ&y�)�K����[#���k]F�1*� 3��ƃ�����.̂%P�N�sŧ��OB�x��!���vY�ߒ��ww��c2�q�Kg��0qЕ*�T�z���WQ���P��8�	���V���v��˔����"��Ӂ�ژ˅��f6���b��Y�󌦲� ����5/i�Ϋ7�'�j�n<�#�bj�'m,0/�&���6�H��H3���52�����ǵ��@����O���>�4
MY}��=�M~���e?��Y
�7��z�#%m�eC���};P�"�\�����/�PdyW�&Wp�U�ϰz�(�- CLBR��j�Zk�����h`�A�m���?BzX�8޴���4Z���a4�{��y4�i�p$b�W��-x���w�V���J��⅖Lx�������K��[��]�k�BF�cSz�Y+e(��.��#���W>��GQBӫ�Mh:O���y?ز0�P	�#3�pp�P�f@C�2���V�q�C��T#x�P�BJ��%T�Xyc�ت`7�@��	��r�
B>�8�=�*m�A�"v� l[��n�ߢ�+��u�}B�4�n��D�Bj��"yůĺ!��G�kÐQ�+�<�,r�zS����f�$�{wsr�}��c�r���ETME?�d��7��:����J��ҐHzX��|�z��0�u���	�Y�$y�����Գ�ͩ=���Ȫ�\=੸6]�!��v"}�_�4b�i5Ǯ:�~<��-��EN�[���u͌�������Y����ɇ<�_3���5���A��)g���a����b��9�ME�B������"������c8�Νf�f �i( �Y'
��A~Ck��n�ֹ�L�:L����ʲ�D��iJ7ۋ�`Ys�Ҍ^�R|�M�)����]�e�O}�2m�ّ���/k�6���|��إ�_�v�d��'o����9E�_�;2{���^~�D�[�2=�wL��e��M� ���$�6�V~�$q���wc!�s;{O�;�1�4es�(����M��gA�Vo����Us����H�1���
}��q5�����L��O͂�:��֜��=�Q��ֺޕ��Q�����ťN�v����"G���Rh�ه�^�V��)D����D/}��nt��i���.Q<H��8���~�-��L|w��Q��5g�Sa�a�qv@��X��_�T]K����O(W���Ժ�evT������<�Z!���KH��{:�V���)�}��Ό�B�A������@�3iH�C"�ϵ���@�C�G�]�m#�Y�
��im����i��e��poW�\�N���A�9� �=�p�?��O]s�m6z\lC�G�ʅ�@�B���[C��i8�]�<he(���J{*��zQ�3��>�P*�H���rT[�%�7e�S����-����j�GLY��u��P�KՄ*�j�V��PN�ȸ�A?���.a��葏��(����<�7��	d���7q��a�
���د�oŬ�ey�� &	�(��5W�p��sC�*����l��m\�w#�Ts}��.�C�������N�S�!���j
���a�8�T�ɞ��<��3�X�4��C������eu���UT����oc���Wv�,R�������;.=�
z�	��腒l��Ժ�����7al�׸0��\��	���x�Bg��H�y�C���~4�d
%լҞ��.�єJ���\j[M�ѯ.� ������tv�YJ�
�)i)��)��0��r>U������Tm�S>��Ocp'T��L@�vc|�no�H-nu�2s5jĿ��jb� ���!�yk���,ix�h�K �0�`K���!"����gU�bdF<яk����#�������aڭ�(˘'Z-\HV�C}��t1�42��}XJu\&���L��� �WQL�l%f�n��%�S4ǛH��=f���M��|�nP�.��}�����C���fA���i�c�a�A����?DLmQ����u�@���w���W��v��O�R�z�����ㅬ
ޟ�xP�:%�{ӥ�=��j(�;���H�<O5u$8�xś�'PJIT4�b�:�'�`������7�¡����N�1��P�Dm?BOT�f�B�V��A���
��~�9L�j55���6'60e���	=���lC��ߣ�ϟ/��u�v��c�L�����:	d���5�"�O  �6mH�8��Œ��W͍F�1����:�ڴBfD��BY�����Һ�#3��T����!�*�~�u�Hi��-�#���
�lB�*A��H�$��V�6ʇ�֫Vv�<,׍������)�p�oA�M#'�H��*i��p��>$�WC9�!�-������z|�R�]-Jw������������w��o���S�\[�HBEo��U.K�N�}!�̠�v�#�/uɩ>�^:�L�*��x��2`��ʩ�ؒ�pUkl3))ӶHP���QF���b���;3u�jp#��|-`Y�����|�_RHw͚[��x*�چ�e�J������y0mD��1��<=��u��ƍ���h�]���+(�
�p�:�b��0�n'gY����jK9�o����P�(�{��F��q��yR9f�؄;��o�hp~X�L�����y!���	%��a��\m���F��|�#Y���E��!+�>�CYx%<��+����ͻWGH"[:P�+���F���RA����oEJg��W2�ouZ�1 �c-�tsņ�s��d�����V�x�I��ؙN�K�0��)�6|�>�_E2s�1����2A����6o>��!�gݛ0�5��s4O�/ Kǡ4���8v�K����1E~Y�DGV+	�,t(ߋ,�l��SX�����s�ի�G���Ԛ�_���_f�cÐ��;��4��w���A���=8�c��q�iĄc#�I�{��إ��f�@ 뀂��$���N��(*�gv��c��&i{`�٢ԜP�t���4����F*�T�����������ξp��o{�����r�dا/��y\\��.eGN	"�s��3JA):
s ��G�qO�=�������"{��������p�N���ׁ9�.-�w.�\<v`�KTv�������;��e�s�GP%qm�Zv����G'h��%�R�>��y�h���h�^_��jC0,�T'G��Xg:�Il�g��a�t�|ps�5l�P�_?Pg�����h�7�&:��`Wy�����$�E������7�o���Ψ0���6ԏ��#I�c췒�7
w�̿�+a1�
ϑ�r��cs�~��X{��g�n������S�[I�_�f�0�F�:g�o��}[^���Z��//'�3�!I�h"$�x�j̆
���x�73gHe��B���C�۠�ND���#�c��͉K��tiD�x~��ëhX꺲�Ć�~}9�}��s��tYo�_B�YP�[kǼ'��j�~�L:�-zL�i�;I�! �S��{�YʢO/E�=�]xK\�$_�P��0��n��/1��K]��(�:�d0�e6l�2zZ�b�w��
?�<"��Y�iϥ������X/�!� ڦ�d��T��W�ok��XR�'<&~���6�f3��#�{/�'1�;W� ���}(d_2���=�)�����d�:�|<Zy:�qA��G;�?�u����2JI����̨���1�9�(���8\L�d�`�S��t�%���醰�	,�N2�N����fe���O\_�l���&B���^���R�:8�g�s䈼�E=��	�[qhO+H����ݵ�,h�E��5�:�pՐcf�J#~`�fL>k��`^x�c��ɜP�r��� �/9�pA}u�I3����٦0������?z`�Ռ���J!�����%��+���X"�������_h%���\n3�D�V�:� �L�W�,\�
��\�P{ER�_������I�8uX!�R`��"��/�,�"�Nd��h�'VrgO�w�j�]Zf���=��$_X�J�BӿBa��~�]�F�T9y :�.�8Aoi&������퇫���!Pl�+V�Z'�V��.T�+�K�mG��Oa,�LZ� vض0��|�,�N5$f���ఴ�Bli�jvkq�\�T�ː������ž� b� `w�3���5	�>"�	  ��Ѥ���>�F<����ώ[���ݝ��a����<w�T��9e��)�W}[1�^<E-������Ol	�'�Vt�J��4�C�9�y���[���d73�#g�.zLi=`S�
R����`���8�}P���i�y�L���F�#��M���d��ҭ��!��9�晧~��� ��?�i�vH��Mx����ʶe=��Y$��0�X�ׄ���kgL�aѯ"�1O��L1��m��	� D���Lv�H�rݗr5�ubIp�fO�C�pYs6Ҷ:�Lྣ�jl_9�b!8��?!�u!�N�f�!�����-&Z�(��X^�ziʴ�����!���8��B���������ϧy��
ӊ��gh)�6Y�ZBڍ��ԬP��N�4������5/z���*�yf���C�t�N�׽`1�:ط�B�)GZ�VH�����HN�X�����k����M1>;D
�Y,���"����e��jj�����ց
�*hzoHA���r����'��zӟ���
K���<�Ti���暣�pF��$��o�S��+����[�����N�V�:u(DGw
U��N�	`�����a=���&���+������zZ�b����x�c�9��������~z��[B��ZD+A[f�W��8� �1�Q��Uy��"�D��2�~�<�y;5�)`P�Y!�����%7��MGr�?T7��d��0�1d�!8^M�Î��B�����I��n}��=��4�<  �6�sc�2�S�������&���Zv�\^�@�!vL�·},W���!��!�_w!�13D��a��H�KX���#͜u�%�3L�P�a=����=-�Oi&�����+�:vMH�;kEK�S�*�Tn�Z�'i��x=�8W�N��#nQuh�WoΗsI�8�P��jb�*�Q^~#���Qzm-Z�R���k�#���Ҷ�掝�u>����Ό�c�wΩ�O8p��IïqXN����j�5P��:������M�
��0�"�����;^����?iX�% z��� [u*Avc��V��X���~Ƭ�5R��v\��H� � �k��I���a8j�`V�iQ�� K>N�'J����y�e�-�\��\�R�0�Yl;�S�)��c��m��"�퇊Ϙ����Ǒ\�+��M2����cr3[��k�2L�Ԟ�̺�i�����u�lf8պN�� m��ƒHJZ����H�W�~���'i$W�)�	̮v����S&*���ݭ��V1۱!Z,��Bl�ߦ��t̽��eyfv�E�i�jγ��K� �a٨��ם2���<��q�q=,;��[~��ކH���"0վ�4|�Ly�pX��j*b�mmP�i�ó����{��9��B�)-F�2�O�;�5�m�|�Ӌ��~�ê'�R�E��<��7D/z	w�VJ-_�Gn~�P�ɋ���FA��`�8p�80�hX4��j� �3p��0���+O��jDg��L�$�z�x�,���a=Q=���/����0��g���e��[
�� ��(.o�7	6����K��)B�$�	ne����^$u6���3�'\�[�8hVQs@_�υбA�H���a����[�Xc&��/!8o��Z���u��>�'W�9���-K-R�m1�ӥP3�a�R�i����!�f&(��id��i7����ޅ��R�����_M�p`;��O���qSZ�X7/��/�����PAUy-�yN T��i9\���VRJ�ڿ.[�(�53�����Ը�Y�";��F~��p�`zH�=m���(t����#��'� Mh�����`�F����!z/.h�(���T��c�5�� ~�ׯ�yĜsI�!1��'=�mN���1���ݻ�k��5��B��e�,��7Jx� ��Y�8:�T�(u駇����<iyq�5�1!�"] �؝��:��rb��w���p�Y.��$9d���l-�ƹ$�c�����nb_��Ղ�AJc3n�c"�,�Ń~�ٳ7�����t���{9s��/:k�pξLa�G�L�Ӫ�C��ɑ�y%O0�Gb��TI�t:�+Q;jكy�?gn��ơ���h�֋���W@�Pl3�cWw�2��+��AJ�S*�/;`�z�o�6��^������-�a���L��&s��+P�|�v~���,�V%뺎�2.(r��DxR�x1[���̊P��YJ&xGk5�!�6�ayxK	��@���`�c��t���$��Ҭ���h�D4��ܒQ
�t��*5QU��PF�f��ީ"+$��
��G��Q���$е/q�?OBS
wJ�
��+M����ԤP~��V�b~L;qs�*�vab�C�0��i?���fq��7�w��tZ��:�D��5K�.(��C���h����d�N�j0�v�����ֲ~)�c�'J���|`����A���s����k^���v՟���� pX�6��dmL����U�8��N��ו���Q{w�r���0��	�Q��31�^�o]{��!���6С0����x�p����tإ�
V�YXJǜ4�b�>珡�K$��Ɠ~gI�R��Lz'D~��<'Hh��I��ofx��=��`0`V���_�t�
"&�o�2C�߄y�S��	i��%	��r��gÞ�B$���O��I��*",��u����&�~D�H��`�<fo9����Q!�OI�s�vB�M��� ��r�۾`���T��_�ʈ�H�N*�V�0H`m!Ɲv�����!t+�4��/�e���k�R�sj��%�E4�����:�t^�d,
��7�o��K��u���ʧd\E�o!t� ��r����4
�A�w �S�6�mń��kM�2��
/=��[1��|�]��/(1�Ps-/�|rS]���%����ճ�)M}Ћ2K`����$�CHh�oEn�AXL\��� ���e��
�I���6kC��߆ ����ժ�* A�/��rT-_sVw+�O+n����:�t���99���S��i�'Q8���>��T������c���h���������`K��"Z\q�C���#I++��Զɘ\x�P�t\�;��]p�L�~:�Z�âB�D�ARڴ֝�)H�q�J{�g��(>q|q�я��g]Iދ�	d)Z
�޸�����n8�u���>��@;J��Cw���`�#�P`�@�5�@�_�0~Z���1(�O��2w�R��AU��,,��%L/��()�T�&o�.�"j
�K��bӠ��K��%��X�H�u�ѷQ�`��KB�L�3R���D��ϗ����`7�ZϺ���4�<���M0����}�7��Xx$��w� �����ǌ�" �~����t�M���Գ��,��ώ���Kv�p͌;0����ư'0{�r�C��A��JВNm�B~	҈�b��$6#�w�^ l� n�V���U�BD����i�a�5m��%8�օQ�L<B���#��;��X�w���1�u�r�"���"N�<ܻd¬�m18�j�������n)K�.%�l��ô�;��b�!Q��>N:�����-�_>,���A�����h��)O$�p �@`�� �#˚��{�i2�q̳��l����>�K>�^���"��c���(N��������9�:ݕ�nw?4Say~���!�����?�<Qԅ�ߧ8"�%>�N'�i�\�M^(�n]��yH���~	�����UB���א\��2����'Qj�ӡ��K�D�T�mrf�}���.�u�a,|�Qa�0��3m�� Q�Lƀ'�~�9E,�3�l�0;�β0�^C���x�S&�>[�C��Vɏ��ΕwI�=��.�w�c^��e�i`#�K���+s��0�=��(pr��%���%��ѓ/�d>:M�ߴ�"�d(�|0�t�u��K{����u?��:F�bdẎx�U��|\�c�7��iL3)F��k[i������ڱ���`��3nF����
M:�~KjL.�����ER������z5>aPG�ײM���[���2tI�b����U�a;�3\;�=�ֵ�:������%~\�ݷ���>�3��:�`��	g����$Xϸ�����H���?�J�W#u�m�^~JRyx�A�{j7�Fq�t���w$kfƄ|{пД	��x���β��l_M㳤��:�+�>[�b���*uż��!J�m�VYt!u]��+�U7��)�}b �dNW��Lrz[f+��n�ܕ9�;q�����a?ō���Rg�S�����\�ӆ���)M����4���B�.���]h�J\Uψ,:�����|���Z���Qv-����gP��G�)���h1�n3���y��F˺P��ae:��������	�	`���i���+.x,�b.�5�G��'Kh	�_�b�a��e�t0�.�nq2j>�C >׈f_�`*k��T������z?Nciϐ���/P=L�^X7�����V/N�Ȕ)������5�5�#���A���Pɹ�;���O틚�|�l"J1��dpq�z���v~w�v��tƟ����W��UA�Jg���~�h�u���"�g~SW���2@��ʭX���x�;���''�:Μ���mΏ7*WB��x[��ҿ*�@d��3��gW���O3�佪$�	����.n�g��ݟS��kOh`��r�ߛ&E+��"K�����cP��Ix��乎2�[̍���{�$����p�HS�#ڈJ�!n Go/W��$�-�\�keU��G���1?(c�8�'�����c1��b�7�0�r��ߊM��Rb3ٷ�(K!�J��b���-^�}}��.Z���D!A�Z-K��Q��qk�	T��U�P�+�J��u:R���Θ��j����ch�	hy� ��7Ɋ�bC�_�J�򷔷q[�h��Rrr3���	�_MT�2��\�@�;6^���ir�����y�ؽ�C/a&(��D�a�E��>J���6P�"@��'I�
�%A�����?��w-*w�L���gSoQ� �+�1�z���ذ2��zMu��u[9;���]�jS 豖�~���i�� I�3�f|4��V��g��=2�����2���V:���+����H �q���Ǵ�J��`5�xn��Gq�I��:�Ǡ���9����9u�!7�ګ��64�M.��N�)m!B�P��b!ւ�1��4T5��EZ�K�&F'���/0�;�H�Q*EB܍�*9�#, !-���fV��CI��m�T��`V@c�?��Y�;h�EL *e}K��;�2���
���4hjz#�.�y��Xe�|�[�(Љ�3��Y��@<h�`�X���:��oR�e���֡�q�iS����Tj
Ё����d-'��nĞ"G�滨�3�%?v|w������7J�G~�ґ3��EU���O��S	s<�V;D�M�Y�[|.<5�J��M�R��4�̚�;ٝ� �/&���l3����m��Ĕ�d�,E�33��~h�����m����m r��� ���Z��G�A�[��@��|u-?PD����"[�hs�˖v�XT�)���E�g,��:�]�\b�>�}�V�������-޲��`z�w�ϒ����}]� ؼ��YCz�|�b�2!a�R��md����a��`����b��������5� �0�2�Ѱ���ڼ���tBS�?�+Y)乁%���gd3:!�ᷟצ?Q�2����I|�Xw��[��S�Lw�b���8�Tg�S*E����5ϛ6�1���xn�w$��o�0����ʜlީ�V��ꔺ#2{�2Ȋi߃4���W=���_z�?��S`�
zU�p��-��#�Ί�x J1���e�\�^�E:���G��� QJ)�5��TD�CMN~R/�@��\(.J�L��	d�r�0+����C>�P*�5$w������۵Y�@�FT��v�KopZY>m�ىS�͎&���>�P]m��o]ל�a y��el�6n=E�����SZ�r��)��G�~p��Ih-,Ev�Xf|�n�ͺ�Y�}�sh�-w̔j����w�F*,�2��G|	!/=,��(+D�|�^��4P�}F��i!\MG�B��(r� )6�v@�)�$<��7ܮ2�3��?C��_�ס,C^{�)��T}erֵ	�b��P�+������!�P�+��8�Y��c�K��NV*���4�x��Vyᙱl�䅢4�ųu���Êp��k���jsBeD�O	0����Q��	�Ƣ?�.pj����U7>�� ��o%�X�IO���O�l�	P����ί����O#�L�t^��+�j]1�}����u󹴦�)�ߴ�ұ>|����r��{����pd �_����ӃCF���nG�P'��0�@iL�al�d�� �Ժ��8�l�9u��B�H|W ��7; d�Q���B���DY\��׾��L��$DyOvwT�8L#�g�L���^oA��F�y��9+KHc���/N_룃�;�Wl��[A=�,�;?{�e���O�9/�fI�
��i}��!&���08O��*˪�Ny�H��
��%i-E��E���� �2����믻|�ܰ\[ԛ����g��5�7#����ȫj����PRkW����L��,�"�9��)�T	��؎��E��Q�h@{�Ax��8UأC�@;�<';Ґ��O�A��믁�����u�� A+v�oPф'z�W�P�����T���� e�ĥ�����d�9W�S�EN�����I�~"'�y@u��c�VJX�[xa�Fyb���e������W`�P��(;�P�φ5h�^2 pCzr��0���ɬ�NoHi��.����E�+���\���-ņ�ˋO߳4PE��ʾ�� �)P@K�t�2�%7����`%Ǒ-z��y�cי��\�Q�T�9ǯ�Qz^g�w��z�l�"��_q(O�m�9֝�/�a���Y��NA|��DR�
0J���p���\��R���0��|�� �����Hx�~	�@F/�����!tw����9�	�q7a?%��qЊ��g��b�K��$�=�R3���|W�f��l�5������̰ C4}��nt��d�*������#&��y]@���07^
�2��4��Ɏ�e�#l�>o0��m�̞�E=�tN�c�9��]����ӌ��#*���k��)z�[ˇ�LP� �!]��0J���FŽ*c��x��
��@�h^1���J�v2{����ʭӴ�7�ZΤ�c8���7��c�O��gc�V����n���ˌ@$к�("�ppQ�'�����I%�{��yF��dؠ�h�ן|xp[@�����sPWq	<��8=畜x�?4�5d�.u+D�q=�m~��V�[[=��8�����X���Q��"��� �g�Q�=G��X!#�rRhǍ�=�(�e���;;�߬��D{�g*i�*���7�������g����`�؝Z���+G�>���Tg��)=.D�	*�M��9�O&�)IX�Sk�!���y�mB�N�Ó$(���Y��2�?
|(<'��s�r:�y���F9�6tk�ا,�"0^�07��iD+���!�x��8r��J�čIt
)�{�!m�@a��2��)��(���p���"�މ�a�����6�9��c��'1{7�؃%�����!�@f+�f�h �cvy�w�~9S|ױ+׎B>@��0��4�I��,���5))s���nV��F��`�uVt�ma�w�;� ���v�s������lh���y�&���--�����/��Aߴ�j����{dl�5C��C�JG!�RU9\	����ʕ��,�u@4Kc�،��*s�f)�}�Fހ(�{%�����4�y7��$��(���}@�-g4>eɄ(�p�%��/*����	:�*oU[VG�_@�h�T���-�=��!�n��)O�왦�^�g���̈́���lt5�&V�[�綤t�U2�oI�1r��ωN"����^����'˞�5c��곝*(�A\�j2�����
��s�����|���`2�݀��L"����
d�{��VG5Ut���/�y�#�c��{	�X��0% ��;7�t�;���
�8��|�i��o��K��/���;y��
���2,j/D�k��Ɔ�\���r�S�"�Z�u�H�3氅�fM�i�?"�-��K[1�~�t��R��r���+���:�Q�yv�a��>���Fvy�'q��GLp��+��f�Q���ߑ��L�L^���E19a���4~�d{9�4:�uzU�d��,kQٸ[ �wu��^	��*<���-_�j���K���Ē�N3�ev���4Ø*����Q��R� �A�B�*����A�ƕ$g��凯e�Բn��X��)iE�w��r���%Ť~~c�ܤ�p��]�G�˙sK�����7�N���@��u�Zߦ�*礜o�z��L #�'�bllY���x�ַkXj�}��v4��v��H�U�@�1 ��޳9�����.�oɿS tи,���i+�;F�ǽ�����̢���!�c����+��X�[H�I}6%I��%�l^uzl>8��{�hk+�R�O�{ld��Ȏ��$g�N�9;h�.�uB�ԥ��rK�f�����"���@�%	��l�#�K2����R������}���AK�`��P��v�%=��&�eb��{���ѩ�j�v�]WP�! Qq�ev�s�P�����ŧcF�'JX9�Ac�����ʚub6	Fw�L�d���H�0�=wӮ������-�8��HA��8(WD/q��ׂ=�荙bt��Up�|�w�af��"�0^O.\~w�V�������{<��v!��Mf�UDq���L�8>�+�D�±o�]�_Es�i9���坮_	��{۩�Ax�����z*[k��Dү�Gf{D���v��%?I�����i��F�0�!�v�"��#[�G/�0���:���d��`ns=��Ujw>t-U���F��5{8uu<��!�K=�G6�z-�Ѕ�"����sr���\���]�,Lˉe�ȫ��:,z�eXI��)���j�p� ������W�k���6��P�P���x)��}>�Q!i �x�M����)csP�<�h� ���t����Ɵ����0��oj|t������Je���y���l;�A������jo )����Q���/ǯ�9R�I������':��T" �3����Q���-�����D�MqW�a%�]���s��'XT+��ƅ@���`=>�ˁܛ�oFu���{�fI��p��b�����%M���8�(E�rT�~n�����(���>1^�5�Ũ�};�u�xl�+Gu�ӥ�!��w(�k& J9>�y���.���kM�T��f��$��e����U�ɝB��{��
�kR��v�G
K���Q��&{r�R�|n���k�2b��Z�p?N�Ig]����x+z:�ǥ���)�������vN�d���x���H��5bL�j̀-<f�Yt���q��g�O}��(?-EA���Y?1���zJp����?�����F��gj�}ס76��;N�2��^!d3Un���T'��+��6�qژ̔6�؎���W���2�6�[3�&���J^��I1u)MH�A��pG�3ˀ�lB[�e��J�"H  R�$��(I$�J�h�����<A��N�4,��� �C�����L<M�Pb�KXR.O�Iy6���$�4��%~ۼ�G3$R|���`���^p2��:�Q�iF:��^�Q?���|!��a _$L~�WU��T	d'vƊ�@T�}��u�	����&ٷ��'Dh����͸ɀ*�����k�0��MrFn!G��kj��9Hqq��7b�����>m��D�Z'}GV�������^^�tϹPΥY�����>�5�{��@�o|�XU��v�XYN'�fj����H�q���Q�-�?��U�����^dn��S*�zz�\L�M�M;�!-3Ap�����sN�I�P��C��)�y N��E����u�{��� �{���i�ѫ�s�QxE�r,�!�ο�+��^:,�'#a�ƀ���H5�J�.�P��{Rs�WEz��ϒ�{ذf���G��V���N�����w��3��rb�40��oKO����9�S��z�r��ā��ɮ��䂩f��.�o[��\<�$t�˶�����&��>f Ε':*�6���&TS�����^PJ��P"zm'�V0�������*a��T&�i�y
��͕�٠����^sY)`�2������m`!��	Ýԥ�	�����K�I�ߜRZ�����ך��WѲG,�:���|�*����VXc��f��6}���1�o�YCă]8�����*�/#�|��
H?ф�Ư�m�� \��Fp*K9��w����$G(���cOfhZ�;g؞5-R�x}F-N�[~��>�v_=qk4�Մ|~>n��?>���RCQ���}@�r$�N<����e�'Ty��఑Ld�G�vw}�K�^A��Lb�%$��8l�
҇(ɯ3m*�\�����"�
ތd�.��&.�4�����"s�>�#��Vd��cS�E%a�˥�bD��`��#k1ʡN(y+4��������Y�Dk z���u}�UM�J$�:���R�poQ�ׄ��G���3l���~�J�<o��: Qͳ�}�F�@����%����ZN�Üd�C�ʿڒg�H$ݐ`�,��}z&ޕ$H�-a�m�����♉))��\�P�u�x�.��+�w���}k��Ӛ���n���xB�>�W��F��&�ޢ����@"�܎&q5_�-؇��z�~���=�7��+t�^����R��׶>�y���H{��h�I�TE��n�0�VO4����.�L�#�%,ot��#_��b��̶�{-W���e�Z��<h:,��������ܧV�n����$reg��F�T�?!}�������(�$@�L��Kw�Dc��u�|�����?~��3gX\u����u��� p*���N������[r=��E,���M�d{�J��|Ǥ^�����Xsc0\���i�d�G�'K�hI~����O���(��K�ǣ�'�[�-`��k2r���7�;�R!0'����s�'$-U���#�u@�T��2���ZU�ۃ����-7VS��M�v�Ca��ѷ�+����
��_�~I,��K���B��@�\���'��G�o��?���g��x��)1:�|����$p��K������+���A���*e�
1Xe���t��:t�\z�W��+u�9�v�7x��#�="�5���tA�"�)l��j�9y�Ae."�����71F��^�J��a-��W:�f�a��'p��'���w��z��:3�%Pž?�s��,�i�6T�P��9���O��L�>����?�`nf��5ӛ��jy��O�wZ�\Co����IQ;ο�g�ƚ?p������(B�j�o�]��|�|�~v�5��<�q��^�7i?��ߌ�'��������VH+��G�����Ĭ �*xm,5��r���$�������{#�ʲi��yP�Ga���m�"Ǡ�������8����PF�f;M�rےT�v7�.ӄ��>-J/iRB�ϛ#b���Z���h�7�{��±v)�'��E��$$��ڐW��@�6w�4U&J����m���DEr�aFIÐS�i$��	�E#N��}N-B���}B�L���3FӒ��2^����1v5 �M"7X���hC���")I$�C ����&X�rN
g���bZh�i\���E(6�n5�`���f��;����Y���G36�f�9;�Y�k�{�jO�`��K�?�f&�T�[=���Q��l��f.����2+�����KOp�����LH�� �ۦ����%��>RS�|��0�LZ����E5���4*~����/�m�0�.��L��(�^l;�L}z�q��/Oyђˊ�^�/J�8�ზt]G(����L��#��w��6�C�"j��*�q�"�VI<��ט ��ƻ	��U.@O6$�Y��t���3�:�SS	u�uQ� HL�U�v��%*�+a��>}P[?�9H�Lq�t�~É��w,/�P�<�v�[�QD	j�R��?���?ORIA��5��<�S�FUn���w[T2N�|`��Aw�=i�A	{��� �Ͽz-)�)n�k���<C���A��H�A�6��Z�׶g�c7�א2����F�G�TjB��=�d���M�l�~˺ە�q�p炄��
i�ׇ�a~i�s)����;p"a��|}f��y!�6F��^m5X�9���\K��������풪G�=�v�S?��Ar��t�S,��(�3RҰD���Ǌ	R��k:&��M�ḋDcv�	R�U]�82��ES�X��3H��ϱ�m����TI��5�ɐ�*E���+.mS��t�Et�8�-#�G��l0�Z�<G�n��>3	��ـ��2`�FeS�<b��~A_�7?}���7W>�޾[[ܹ]������Y��W�k]�~�	��b���ZW���h�q-x'���7�M���9�Xс���
a���1�	� �I
8���҅3�.2��7+�{��e�M��ȜHPw~B��s�ؓ++�^*�gu
�ԸN�R�U�WIkC���F��+�����3z�a�ݙ��uzA,���ѱ׮^�\
\�4*���T��&��4!��Z�e5ߚy%���o�[��o3y��_�}Z�(��Cv��:|�N|b�q
챴��b���܍l �Ή��y��:��'�+�1X�I�b��'��C��>.��av]�(�E�u����=�I�MK	��-J����NȄ��F�t�ź�;�m?F>%6sU�"�G������Żv/�{�|��%��y�]����2wbD�����#4������1�rM�(���� -�c%V]Ԕ���<5�:SuM����k�.��\k��O�Iډ�I��2��h֏��*2��7v�%y{���@(���b�@�[c��?(b*_�k��x�T,�|�-6W�S�W=��@��Y/��y�l!2d$`�v������en�����#��;J�^7�{s0�3V���HK�����5�j��+�}Y���A��A��F�=i ����:Fۥ�yjFF�B��RQ!� /�.��]�U�il=�G�V��	q;,l2[��� si�c�H�<��q�:�6Ȍl��e��g,R����O�4bd�P�4��-�����s(4êx,�H�5��0$-J�dE;hl�n������~^t3S�KQ\�ǰq}Eq2, �c��7�;���ytϨs&eM��(���^^�H�We�\�J$��k ��@�d��n1_M��ou.O�sͣ8�V��3�[��F]o��_��fBe����0����ی�Z.�"a��n��}>:�����!^���>(^.�:D��s��&;�砬�Rdp.����5�`@1e�%O��62^zn�r��U��崇�����I�'�FS����`���ͯ�cy�$=�a"l�ee�U� �[�H�����!kG�0�:A�e\n'� �E�G��J�r<?�Un�gd�x��k����1��e0,�drYkh[[
&����p� f͝5����	lx~���z5���QǟQmĂ�c�e9����u�9qJ8#<������`��F��d`WK��;	�Tȵ�E7�T�`� %Q��EͿ�g'CO�L�α�����Ħ�$�\__bq����{|��i܆`�F�<	���U���>L��Z:��n_Xa��3�f����Q�@�8��V�ٌ�7� jV؎
ӄ�L�2�I���9&��JE0�pi8	2)��N�2���<t'��Nh�6���>쁽�a�k�N#�� kmVs�$XE��}�
�^���8{Lc��w�\�E�b�6WB��m�=��'��Z胸7�I��ܦ�\ͳ�D��ǩ�ƛ�ǌTg��Կ _���ӣ����%~ɟj���u����t�1ꔖ���8!�W�|r�	x���7��hu'��A�{R�)��(ot ���^ƻ/pn���-5�=����qD��딗�a��J�d�/� e)x1F=��;�R�J]�>+��dRV"��z�gU����1��T�S1�r���x�&�����n�.Q��zOo���ȀP��@t� 9�'���f`�7!�A��-'��r"�P=���=C�~�~3��2�L;�7�u�-s�^�!��+���2+���2���0w5�7��b] �e��@A��6�J  rZ��+�0Qd5��) .����%�C��m��5s<=�H���X	7�}O��vG�^A5H�����<����yǃ.��w��ת� �#R0S�q\�)o u�/(s:��~Y���k�T�kq�5l�L�V�-��cK!�|e����NdELi�y��V�CB�:v�u��{��� �s�4�g�X�P�:v�ۭ.r�7�6�(�<������/|��&�j��E�G��G��2��]دud�_!MK�Q��#��[���)ܑs���I㓴� �߅�t� P�=/�C" �H�+��4'�uMQ�Ю���|ha���q���r�P�ZOf�ZF�.Er' [|"�8�i:���O�1:�U�4RG�R��
�z?�}�Vͪ��
�&��@�˜F��,�k��C{!;$tS�8v�G����|V	�>��w_kmt�'t&u�C�\�(��T�7�^�b�wAَ����g[}rB����޲wu�����ʕy-�����{��I
�d��G�2I�:�ss���RA�E�w��k3�d/�1�Bc%~&����Ր�>��6�sK���e��r��8��-Κ����8r��rA�v�HI�]�N�
 ���)j���>��ә�xQ� J߬��oY���}�po�Q,J�&OԬYNk�W�Up�H�>�f����Z��%��q��~���v�d�B����0H��?8Լ�ZH>�h�8��,����q�>��:Ģ,���#U}����U��_�uF��ڟ��,�?��N�"2Y:���'z�ɡ���Y�JN;l� ���f4�'~e�b��<7N8�վ̍��Z�-"qPѐ� Q�������KX��K����4�OI�9 wE����Z��Uk�,P�oF$�P 4Ƈ�����ޠ6��%�)���p���[h|��(ՄJG��Ձ��O���+��`�|��&��4�P�Gֺ}������>�ü%������o1%�@(�6~p�V(��S.�U��x�fR��--c��r�l�z��U�w�.y� ��(��UM���@�އlq�jK�nGއ�|��Y�p���x�W�ئ� �:(;\����b�7��y�A��^g�/+��*��p�[�h������J��]���j�)ʿ}�/����[-y���A��'Ҭ�֩~�P(�
yz�}flF��k������s������>�"T�Dp�圲t+D��Gh��׸{�}r�4��m�H�t�pg�]oG��vL&�~��Z��IF������~���juTE@#����&|5�6�M^;@`��~��S��v��	�y0��%W��yޒ�Y?����	��1 ͈S<8�d�?�W��Ёr,/�-�Z���������tM���C�fґ+�����J6YB�X�w�sXQ =д.���GSƇ���Eϗ���Z���Rg��uُ�"ڭ��p�F���$�Ay��� ��u���Ae-�.M��1V�a���&��j�hQ�����EM����1L(�2ܬN찭�k�	�U�����bq���0)֋g�(��yd+j�E�ᗰp���N{��gV���)�N��A�B�{=���Q�*�&���̈́��d\r`<ɷ�s	�����c�X���[���\�"d��|��g&�3�_i�k�4�%Y���P��]��³YaY)n=nx����ױƭl�j2o���9:�Ep2w��<��m��� ^��FQ������$DЋ�hpp٣�4� *{�����A�J�$��
������i_�$�z}4����ּ��a@���$��}p頇y�?9<����]A 861������*�|Cy��@?��-,E�r�@D7ۗoP����fO(��q���I����@ 흠"l^���܈�N�x���6�6��r���=ʟ��_6u���q�:�H9���tFb���cB.�O茐�2`�8�Oؖ%�"��W ��cl��x��"1�l��N?�����_����mC?��K�$���~����%����/o@'�y2o���?G���z��r�򲴳J���*����f�P�����A+���uK��@�B0����kiA�82�?˨v���=	���
LJ�Ԅ��ĸ:�}�n���k+�86p8�J|��˿�Up�_ 
l��ꚩ�J�������g~�bFN,��l>1�Ԧ0�x���hk��1��*k�Ǟ�z̛�`N4��)[�Z#L�+���x)����$?��<jn��2�`ʸ�/�b��^R2�qg�A�p!���_�h,Ў����֫������0t�ǅ��{��E2����t*�c֮�?��,��	��U9�8:z?�R�q�O<g~�����+:�� ���ǯ��r#�q��&���вBV�[i4K-��~�hg�Y��_c�R�qd �'��` ܗ�m�:R��VF�ڭ��pDx]���8��m(
�'��� �SS�}c�.�|6�م�f���C4�H�_w�pWz��M/V蕤K+���A{E�Z�t���4��.��>h����/L���r8[��(uj
 6C,�U���qM��^�"в��Y!#��"u^��;9T$�ִj�*������J�|���ȁ��f%[��l	���CE2H;c���_�zV=���ԃ�w�;��}��a�/$�3a���	�ú��n�Z~B!f�0p����=���$' �9���@�ul�+�NC}]����5�4�HR�ǁ��E"֎��~M�6�B�V�So�������\����DQjHI���:�FO�՝c�~�>�؇���j�œث2�e�	�"�#��T��c3350�U�|I2����*�6���� ?^������*���;c�24�"QV��G����������<z�I D�<vD��6�^۽�D�y�c�i_'55C{pP�U�9ȗ����<�����/A�3�z���$8[-Q��a�3-=��oI�I�g��4AP����Ѽ� �%G���'���PncJ}n�����%��4��TJkXnb�Ӷ�)���.�+�������	���A`�N�d�e�ئ�W�m�p�6%�M����(� ��DX�m5��5�(E7��>�����%��e�_�Ѻ�3���,aj3���O�$�{��L>A,��!ЎJ�b����S��CE�?A("�E�P�Ƌ�<�2	[�����L�������WϞ�[c�a����qӬ��-W� l.�/��G�Jh�����a��o��ϣf���i���V��n<�	L;Y�Qu����/�m��5=t�)�j��
��D��"E$9B:8^Q���\M4Ν	[�7D�O�le����K�N���5�?�����l7�2�}̯ʽ��꺫 i�,Yw��r
ݽ�Ԕ?�� �N���7�z<�o��d@jȴ��hR��"E �Cm6B�O��5�J,��0ܼUw%K6��Zu��R���]�ʴ��1�c�7�洹��I�+A�Gs�*Ǥ�s.G��*����n+�C�Y'���m!,�?��y��IWL�U8|x���*r��
�Z�[��p��$̇+�>Y��-����i��9~��Z�O&[bO��?S;;6��ehg��`�<=Z��2���D$cF�� �&��H�G7s~ј����"����c{�jV���p�؅Q��dX�����}N�s��Rŵo7��n�؝S��9�[�S�+hy��:��T���g+��p3't^���u5�&n��`e��?M2���Xq�f6�Ο��pT�Y1�S��8'�.�{`,ˣt�ڸ8��]�q*�op�(M�\*�����p���ہ�l���v����h�Ԥ��첢�xl�����`ݘ��$N��yu?E�n��A��p�G�XZm�wZ�8��Z۶�W�ꛯ`����/��;ȫ�Ĝӥ	[<0�������W${6!$��j�-�E�U�[D͘	�/B")ݸ��Obѽ�̲^��{IH�s���$$�ʌ�&KG�H��7����Y��pW\��	e�/MC�R�Ͳ�r����`5m��H�"�P*?dm���쬣Sb؁XT��q��-� �L:��������<���<�_��w?9�{{�lC �D�6y��!�4���q��"�^�4�;4r�P����ZS�w�����JN�9�Z���V*�Spc?.U;��N��`�h��Z��{����B/��ƒ3w$M�N��~���k�G���;��m���m椄��1���dB�Y�ak��ܬ�>�8S��F����0}�ں7��|�k��ɀh�����E+�(o����Yެ�R�Po����#ܷ�T	셣Oy������:� �M�D�4��k��i]�$�.{}�:84P��~� s�Xn/&�Q;J�_�mon�����K��$�j<�ޫ�*|k_���]�4��
����a���w�ul8t� *B�ρw�I�O+�v�3;������(��3� T�"�;�C
�[j�/�����۸�6�ë\����K#������9:��\��E���8�׾��m5lI�E[sL�
�/# ����d�izp�����K��M���N$E��i�y,�ϗP5,hba����F2�U��M�i?S���xB،��#��m� sD�&VV>�N���eh��Z羈Nj��]wK�ء���Բډ5X�4�e��7���DE�y���?����x���x��X-޴!���g���u�cx��t��*V��s�����b�qSXse���兇�`���u4��5��k]S�c�����a�z*���K/x1�ɡ5Q��v�I5$�#%�3Cn���8'{d��\������2_�ݗq
�JP�����q"3t���m�SA!`^	��}-�w"��(�+-�w��'���O�#<0�ዛ3}ގ�y�'lB�-��k�>�-n�� s���SZ�h�t����d��&!܉&.G?��6��&����������@���W*Q�-�qU���P�S�	&(�����v-b%�+�$�3c�k ��$�@$;��O���`�hi6y@|z��&QaK� #@Qa����O�]���t�jud�cw��Y'�qU�A�������xB}�F��F ��f�%�<��D_��w�#H����p��h1Eڗ�)�{��^���-��H��!L�����K�Gj���a�M�4�
!ίv[�i���U���S��\������|
w���L��'��)���Ծ �CM���e�[��](H�ֈZe�j_ kq������Zٍa7�׼`��m?�M��_X@X�n>qV�C]��P୿j�X~�dB�{���?�|�$�@��a�3+@@��i`�Yg��o��+v�|U�x+�q��-���8K�b�'UW�G��)��
�'�t܁=��aB���DB����S���-K�" �]HS�m8wN�"������Y"	�:;��e�j�4���8��~ջLcs\*H�Ԏ�L��5����	�(~MA�qA�|Tg���#�p����nb�?*���|����tP���F|��gV8�W�7zrը+'$�ۈ4�<���%s�	IU{�ŋ�f���/�J���XX�d�g8�T�Um��n�mg��0����OH���b�W�w6{�4�p���F�^`���I7?��˥���y}9�>Q���KS�*{�:)*�Z���(7��:�}���;��b.�c@��ޑ��k�@#i�q7W`������G�Ti�������~���1wR�̙��w�A	h�uu�/bM�
l/�ŋ=�LHx�[��ݯ��U|��'Ù�z�^��e��;��V���X��rGif8Mh����p��ə��P��Y�MNo�\���RIKi��(wx*+�;�T����*5��X�Y�O�o��"�����C�Yh���D+L��Es�e.WF��Pi?�+�;r4�P�of�S�I���^��&뚀���~�^Ώ3��+�����Oa���'C������m�&���R�8
pc@��L�2Y.m[B
�e�x��"��V�m��i��s�d�sf�4���VX��u_TO���g�Z�uh�����\��A���()D$Db5�ҕgԸ\�D��Ul����W~'�`�V���H�n #���G�� ��*5���ΊH`/O��>����<�i# �>R2�?ҍ�k>��u��g/�'���3Ȑ��-KQƖ� �W�==>�F�{�L��A8�ʊ����=)���$�D5#57k�X@@�I���"Ek���K�U���q��-玺��>6�Ki5���w~>��\�����ZA���N, $(�o����[�1�T��}�,_�׬���<�+�~�sZM��$a���f�_�9q�
�>��L��F�/�%����17���Ͼ��㆑�����h�!�џ) �lL����Ej1�Z�e�u7aF��,�&Yh�v�ss��9�@	;���	�%�[�Lb�~3��8Q���^�Jq�o�Zd`�� <�Ę��6+�m�ITe�v؟�-��=���Qв��Iл��mt��-��B3�-"��9n���	ry�PI�=��P:�/7�6;)�I���I��"��� ��W�,+a�x�$�	�{5����#g�*�g�TVd9��m&����G���_Q>R�lU,��P�NN�+�D����i�Tktz��}Ogw?��h5���Jŝ� 7���-��Xo�D��ǯ��	77��/t44|��V,}�L?P����� �=Kd|��&�-ȹH��&�3���x�s?4� w?�� ��+y%�ru)W�� �"�j �2D�y��@H����fn >-��LO+zA>��T���q6�z3�FQҕ�Ņœ�������]���SȜ�p��"��G-����l=H�������\c����Z�jX8���-����0���-�t��LR\��SK����z�k���2�f'����|�	f��`^�E��z���_|3��{G=���ہ�`߮���m�z�O��s�ղ�W��c��r���f�%:/	�L�����iyC�bـ�y���t�۱�ʸ�)���*	X��IM!�huA�?�C>M0�U&PL��0��a&��}����2��;v�Vu�J��5�.p�-0�)�u�g��u�i�!v�C�x�+�CHC�H���DC���SU7 ���o�#G���|]����!�5P}� PC��K���t^�����{��K\]���oXmq��Ϊr�-v �YT2�_ �<e������P,8��'o<�W8�����6��'~��Z�[������2u��w�$.����M��?]���o��r�"��oel�i����Z2����D���.�t����3<��>��V�AR��;�Q2�����V��ĭqW�!iO��58n?��WÐ��:ڡ�n�
���X�H?�rR���[3p Z$�Y���OT�{��/w�^�f�,<���ޙ�G_��ej+�e`I������"�/���V� &9�N|>E�o٥lGA7L�m�<�c�����~S�`�9=g[��K��u���k|8��:�F�)DM_���P���V�C^�r\:C��`Zd��R�i��}� >ZJ�X�^3�$�ec/�)u�$�����((��F#^�&A3�gִ�*�?���Hd��A��
AD�=4�n������T6�ًM���#�d%��:c���� ���Gk4.�}�\�!va�ֽ��V���$�뚝\��kbe4�)�Y.%���� u�E�FqV�`�%2��w�Cq�~.Ȫ���np�IWWS��e�%��Q8cb��+k�Y��}��*���s�.���<<.�6e���w����G�a� L�ðl2�[K����0��/IJFf<�������>d"T3�׼��6�,��y\땇kf��Y�|�X3��a��c��]�6�{C~�n�x6$l���B�WL��W���me ��^Ζ�Nq3�o������s٭y��ҸT�B���R�������"�7�����$�,G(q��|�Ĩ0�d���뗤Ol��E�X��V7h�yfX�<��[���w�4
)��+���	g��6���x�;���8_~��'v�N<_�E�G�w'vМ��B%D��@jhe�c� T+Cާy��Ȇ`vQ-�#iR�.�$�V]-�m�ƶ�����ѥQ�Of�m�U��p�]#�yjK`�3��w����.�	Ό%���&t�X���J���Y�r}l�����U�����<ȥu�~�+Ħi��ȹ��?:�O��@��N��A,�mLcv@�]����t�'}��S���E���RӍ�� � �0�)�'fL��L��-[�D���t���J�J?إO�2tR�G�������9�������-�>O#�=}�P��F|�p����EgP�N`]`H���mW���o��\��,c3��p:΃��>�rq{;r��������p��gG+G��M��D�N��CY+��DA>�c���A�,i qg�3��s�x7Uϖj2���( (����?��~T#�W��r�jFj��ڈbeX�g�Fa���)U1?Ms�̓f������G���+N�?`vLC ���8�P4~y�O�^���ۉ���.�I81~��:����_�{�(��;a;�r��U0o.���2!�c�ʅ�s9S1�퐯Q\U����@W��&2y ?�?&��5���ް��#��Z�p��^Ҟv�7�Q�����9>�jh�a�qo���PҤ��ua!�4z\-����t�>�fk��DH��Ə���х����;����z�d�H�,�	�B�ZS�	�~���4��
M�V�[^:,JS%&���	/��C��2�U�����n��v�$��� @���|T���|2�~o �xDu��ř��#:��\��Xߚ~���*`-�'N�'I2'�7Y�m�;�m(�����}��������Zu5��bNr����v�z�B���q��+ ���w�R��t<�+c�����#a����)o��$�k~�(`������(uq����yk�h����"�V����Z#(��*�̀<gCS���Ǖ[�� ��U"˄ɥЊh�ԮR�3��r0��Y�ځ�O��🣘�{��Sd�ֲ`��Pzv�Ae2	�H�,�h}?�X�<��f�������EH�&06_I�R��V��6�r �������(�\F���V9�ru[;�.�[�0��Qs�!� �����
��i��{��F�m�k�������8Ű־&`.@��Pwy��$ҏ����o%ł�s��A�S�ipb0H�D�~��0�.A��TBM��j�V�__��:�y+�l�n��>`c�`c�r��Z��>QI^��m��cEn����L�B<�o�݂�����a�a�%�����!��$S3�<;�AUā�j�@pJє&�9 ʭ���>��\�5� ���i`S��L?��.&���a�ܳ�m��ٹ���w��ؚmeM !6k�^��.�e|���j�%�a�zܞ�ZЕ�J�m�mx�Y�u����0	�����"q|�4Q��]0ƞ�`�R�FzY����a�A�zzP���4�q����E�?4��jm�3TEn�y�)Q��,"�� ��~Z�̒����ꗈ�O����{uŘ�|��I���p�ܙ&A��y�"=�R��"$9��q}㔳��2���v�Vh��O�MK����V�_~36�~�$��W[�M��)��z0��q����:Oh��-r<�֔d�]~���c�0�Ro)x2�WĞ�ac{䍸o����:�0'��!��?[��f�C�W[PwW�w�r�F�~�h� �;-�B���{�a�>8H���7�Jg;Mc���-�¯����#1�[y\4.,5�{��C��F2�S4u5�Bs�d}�b��Uq�:�Z����n�/|�H W��56S}�.��NB��l�U(�/m5IG��/�AJ����9�bZ���W���~�(q*TsB�������Te�'}q"l����͈sY��Pf�fW_�T�z(Fy	�mz�8�,��B2<Ԃ�+��+}����O�-k�(��p�"���{��=�m�C���ə8�3���s�A�{kU�W׾m�b*�������In$@$����;^�%sR�ޑ���u˸R�`���25���RS���L�g|M&�.x��t>!�ؠ������M�Gw��q��̤^8��FJ�cD�)\[-�$��|�U��Y��m��ۺ�$B8Lҗ�P�"Q	 �!�n[���U]zN��Q�~�wkA���F� ܌"��Y��nI��.���=�GJ��%m����A*���@h#i�`*>�O��К�-�tYm������&�dWT�?�?d�d���6$�#����c�c(��<�zpq��u�r�y���}6z�;��ǈR����1	jǱ�-ڊ�edV_��r��l��2�J߭�T���F�>~���6g����6k�fcjjCC�>�Gplk���AB�]�fe�S����3�[ud�/ϙ�u�û�GrЄ��|<�
1��2����LSy���8d�Qt؍���[����؛Ϩw�A�E���9�`g�|�}1�p��(APIQl����ǭdAZ�k�@"N_F�=m�I�����N~�#@������.�0�a��N�޵_���z|I !��hO�w[�wXb��O'[:���+Q��>a�Ni)N]|��.�ա�_(�h3�����~`d��`m���iחBv��f'+h�q���i7 ���?w���d���C�[<�\�F�t=ڟI�����ﺠ/�E���CLC�#E�2�ҭ��caNT�@�0�Ŵ$ޒz�wۉ��c����.��r�;s�E���s_-�x�2�d��R��� � ����Zw�M!`v���U��R�t%���i=m�ҨKg�p��u���TyZ��@���T<��\�e�i�1Ѝ_��lpM�b�Ƅ��8gs�F�f�^�I>��������gXt5Z 8�^7�$���|�N_���
T�<�cP��9:���è�7f�!���d�8���/�/ĖN�*^�sګd�a>mK����&����J�L���;��ޤQ�^�`�ZPP��_��C���(��
��H�b�T��նs��M����CV[�ȗ�;�t��<y˰%��EJ�HС����I����i0�Ր���o�����[�_�$ձQ���`��� ��������PQ�	��~�,;���O\�2P�4�G��ߎV&f�i���ey�{��*k3dG����L�+	�%zՍ`^����e����m��j�R�L��Q$�(�Q�e�:>�O�� ���G�K��k�����#��ZP�2�f��J��5���p~9�<�WaU�F`�������9���  1��#}M��au���.�6�u�	�@PqX�����8���b���E��m��ŨK�l�!���Ai�e�٬EE�`8�rA�}:�;�lq���_���fpW�觇v�Y	�m����f����.BHd�P��Y���e)̉"Z<~Ϗ,��&��H�1	e�u@�ȟ��*n^`��o��`�!2Γ�O�]g��p��_����$퍡�pW��4����m,jo�o�R�MM�.]ȃ8sox���V��C``���"�3�a��j0��l�y|�#�>�U����C�h"��ha�'N����?U�ΈMw�w܊M5<1E]�;�	�5��S�w-r���6�]��u����k�3�$iW�i~�vuFԼ�;-y�[��*T�{d[~&سL��x��S�ἣ�p�,�����9Bk����:��U�t��T���y�U��YeH�ka��?(j;�q�d�%����R��ڗ�>�D�����ע����K8(��U��%b���wp��3�އ^�W�{���e��d2'��=���YPp�G��R���N�F޺�^/�GWj1�󝵘�VDәc[$#����ǲfzg1V߲���Hn�\�؅�VMp�a���an*�q[-[^j�X��2���X�$!�Y�M�1��}�[�F[!^�R�g��E���q<7��������w:�3�Cd���_n��4�p=D,��-
[��;n.�^�?C�d�������$�2D�[�ߖ�
�
`��"�헦�����*��0��1�hX��7�����ݑ��[�!��c�0�G����M�2r��@3A����*�����́�Im�y�-�@]�EN����ai�Z�&�k"�1�R4`�O���|�]K�ds��D��������,(O�W[y������J���Z5p��8.���'I��q�'#��#�}^����Io��~C�\c"�,��yr�*�}�fI+�%4Z��u��	_���E=M��B�6c���-p��|�����Fu~��v�� :	�U��S�E�|����R��ik��:�+;Z�ɍ[3s"��J,�1o� ��`-t�/k[q�Á��B}g��}��ʤA��~���o�J�s��u_�L�� {Xw��R��ԢV�b�H��m��h����l��|�iS$��];)ꄴm��0`ґlfAA��o�4?Td��+oG��K�;��4�	`�?�Q�p/p���MuXr̆��]�����|[��⒂B�y����H*i�vB	�y=i�>���p?��Ϛۊ���j�c��%{^_u��2�w��B:�/^R?�ת^c�����b�	�"w�gMiCFCk=�*4oUhcQ��4?TV�K���p�~xR�)��WA�Ur"����g� sQxD�A/ҟ{K�o{�Fہa�(�.�����m݉1 �5�Z�<˷9���+�W����F9�^���H ��!������+q��54�����Ǿ$qGkҐG58�h�kn�^OZ��#��D���U�ޭ#���Z���N�F;�sh �1���,D��,0V�e����0M��W�+uzуi_����4�,����	���*v���(�׀e��6����������g�1��!�^�#���n��yBX��(��J�P�o �Y1Q���@�Y���P�(<���s.�	ta�D�3��޲h �X)
ɔ�Ї�8@��qb�]�a���aJ򻧒X�G}�I&9�U�/c���pbs��vX�^8�?�d�M�Ut)O��D^�ù4z5׳w�={�%�i����ş�p���ɒ=����Ql.L�[8O;k��a�jj��G2Ӱ��o<i�;���N%%�f��da�C����u�IL��h��N�L�7?�0Q�l�~h߳|�ف�?��A� y��.P)Έ�/uNGS%T"���S��LY�eÊY��r��D�b��M��:���`U�뗍�UT��l��5+����N'.����5��[���^
��$�s�q���G�a��X8�����4Yؙ�T���-��g`WE�3�$�k>f��l5p�3��_j���5���a�ѣ��՚���8�`�A�y���'�UBX�Q-g!��b���+��-u��N�\h�� 7,��Oe�~�/p'�&�;q�zX�}�-̸4�PQS�v6h��{A�0���v��B3%���~h�IlE|�bN��l�8F�1x��Zn�:%���/����ӎ*��*�gh��n-��3��)e3��Q�z��D躦�0�`:�Yv�8㚏q�nY+dVs��V�Cs���8�
z��HR��O��4O�H���'�,�J���5t�=U#�!��\�5�G0<�ȩc���{[1خN���R�\t-K��E.^n��ӂGN;@�s7�t�D~aMic�3����e5M��!�i_�%Em,��L���(��W��%/�(��M7�d���O�������??Pn�Ĺ��^��gXV�4�W�a���W�93�^K~����-�[��z`ж9b@#@G�)'�ο��)�\�N�1�B��x�
Br�C%�q	0ڎ�|S�DĈެGa��"�����h�������G8N�A5�jTh��U-IS$��89�Al�0E��Z����]>;,�s,YE2��)8"^׌.Q>�6�k�'�/�,vje�B���R��h ���Ց����O�s���bj� �4#P�V��@[��k�ً�=c���/q�� (����M2R��MS��/�Օ,�g$�+�_w���$�K�o�I�<��]��J{����c��A�zM�w��f[���v�m��|�@�����:�~����dv�Y76,A��\���H=����aq��>�����B|�&���̴\����/3^9�Ѕv+v�>ݔ�4��Y��Q�����w�{�ԛ�I#ER�Ԃ�5z�u�]+�ַc��J��	����q�[��N����:��s>��(՝@�-�#�V�v y��?�%[�7^-?�7�qŗ�sg��0M��hM��rE�d��"p����غ�uv��j{!�XQIO���b�&��ʕ�	��(����{X�������0L*���B(��bĽ�reŃ����9n�"_:*π�u�l�-Ν�+��	�QE�AZ�b���$��`�,���3X����Y��֜S4mo���?y �ܹ�HX^<��?��.+��3z��2Y@�1*p�xB��5���o��-��&Ƚ���.�� ���C��DHY[�p��'��#VTV��;�T�7��y��e�1�=��q<1���f��F*�H��)T9�e��"��DOw�C`�.7z�Y��>;#���s�#$5���Δ�j����0��ax�%g��a��2d�U�l�<��GrkF�S`'��E${
���!x���%��M`G�1� ��	V��S���:t�ck��dw�,���bS�C�f���%���de��XB������4RS'e���䉀�zF{��K#o��L=�-�~�6���L	�v-A�� ��;k��#�u6oH>�I7i"������4��V d��,(2gOS2�+f�; {y���H��ݼ������~?�UQ�������PIg#	A2(��w��Xإտz��`���IaT�\��Yko�U��x��Q�h���HQ�SKӍ�!L�{�T�}���<U	rS��=��(rf��%M���U㨼UV�4\N�<���@�nXO�/������ɤ�q����$��	��7(i���#����߀�q�����Hy����Sѓ�r����彖e+ղR�"��	HI�ࢦ�md��Շ`�V�P��vF�C�$���H���T�.�G�i�Nm�����	l 0C{3z�V����h�E���N²��d�Eo���+�Z����\c!NP�3Q��Ȟ�|9=����L����p�ZQ�fƅ�Q#�!W�&0�U1�f��E�!Z-�q��i0�����h]�cQ���pF�V��c���Ş�"j����C��b�X4Ld� �W0�
O�Dt*��;y��mŝ(�&����M�F2$���\���d�#&�*ĎK�Z
n�e~C�Z�%�\�\ث�ѭ�$d�<PI$�+ߧ�9Ĵ�DC�ǢR��0��;�#�Ο�q�Kd$���/=P�X<`*�R���������BĐ�4T@�z���LJ0�Mk�ֵiW
����5x'W�U���<�q'?��,r̒#�~��Jb�p�� w����P!�#h[��-�h�,9>���Zu���u�0�֪�Q눸������ME���P,"6]X���0@�fR/���{:mk�/���X�JdޥMc_R�go��r���
�"��3�*5|6C�o�c{�;�Z�1/���*(SAg�Y�5>0n�����
p̌�9����lt!���C�"�Ag���,7�l���o�Jh��ko\�=zb�(���'b'�(j�~��=�Y���l�>�(3I����G%��o�9/�fEtfzW&�e[��q��}0�\�~5ݘ�Y�d{�β�ķ=�U�ew�/a�{�����s�������|c>�|�����Ԏԛ^�~�� ����^�i-�L;�4
W|#��$�Y�U�H����22>�	��a�-R8��/������݄k���oF��jf3��ZP��~i]�6��-��$�9�zq��b��u�o˷߹� Fk��)���N'C��ԩP�-�ɢnx`� �<e�Mw��M\Kf�8��&������(-#��G���c"�j�7��R�P�G3��E��cl
O��v���\^�75O�^*�Gn, V?s��� �%`����U����q�iz�}l��7�/�����v�a�/��#NL"�� 7W��Su�e�R����}�{���Bo�Ob�KL��,&��?��d ��?��83����-k���3!�����5D�C_5I����b�u#+74V_�u��웚�I(�q��3�"��n�D/h���O���Nd*B:'��֞wF��7�.
-֖ӆ�8n6Y,�o���qs��OR �a�ɴd�م����z��&��cx��9C/���8|��6�_�K�m��Q�T�G��I��Lx=�Qw���l�(q0�S��=�C��m�X���F;-D'�-�9˪W�`D�R�H�|����\��ʴK�²�=��!�`pM��D8"^�:��<��iH�Fm~�
�8y�%��$�g�
�<~+�\!�|졾Cf�!_qm�7S��!��b��Qg�(���
[�|!�8l!	�¡���E�R�'����x'Y>����cR���e��0�ĕϭ0s��j$�����g8P�R"�C(5F}F�f��q�N<D��a"eiC�N��/G�IQk���y�Ƽ��9�H�݃�g��V���2�W�8Ѐj牵}�dU5���m��N��6	��&��ض� ��Oϕ{dm�S���%�^����hr��t�|.䄫�K�T��{����љ�R�:`�[��Ԉ�����j>�`�S��]�K�t�~٣���d�Z'�s=� !����aunE`"�pg󎬪y�����u�"����q�܄�TME��}��W|���v1gt��No v���3Vz�"�4ś�0���T�q�ʧ���If^A�>���3|����I,�_��éZ��(���Ӥn�ć�����f1^�o�),>+�	������X���`�u������kP��?k�R�On�
M�e)��a %�ehcE�� }|ő6-�3a��%���Υ�[g#E@;$�ޅS|��N���&\��e�\�6	�JB��z���#� z�ѳ1���C+���{w��#��@�����-�ǘڹ�U���j�gI���0�~�r)(鞣cXP��,p!�&0D�QO-N�M�X8rt"@�5�)�(�}��iגR����+U=U�����J(E��D��I$���c�i.��u4hf���/�,e��t��%}� 84Sn�TM��!��kn���âC6R�x��إf:R�{���߀����3� ���c\��ϫ*��I3뾎�j���;�
c�L�R��ݤo��a��e��6��=6H�xqH�7���*�
5�p<�w�-^ �IFy�4���#����Y�Co�%UOv�?I��g�O/q�`�%`o��lK���l�\���8+M�$��ҏ;�'��N~�y������4~��M����&��^��g~�����S�o�u`\8���Tr�j��j��!�d(�dw��w�:p�զ���1E����F�f�>�=��h�,:�xlr�?�l��6.bV$L�Yl��V�ɡhO�Eb����Y��^"G}�0���Z�}�5d�e�<qeZ�ʎ� 
��֗��R�N�ȉ.E�gô��� D ��C�E�T}ߞ.��=w!0�b�ӈ��5^ik�^}��\UCkv�1��H�գ?%w�焰!�.�����(wGn�V�?6���c�LyEr�]��A���,~w ��/L���0V�W����8s�7#\ɳ��j�?BG�hTR�LZk��TТwV���-M��V�k-K�L�+|^]�YT2ʎ"O�q��ڎ���xg�u>��`R�e [��CٸE��� H�b��.Ti518���>�a@;t�:��(�|�V��ә\�DuP#3�{9gv�	��A�^H�C���R�3��`T~�M�[Nc�]
��*a�����-��B��gt+uA���F�����R�(^o� � 7�rY�4��>J�a�:7�}i�w+A�c�~�>���%�ԁ �c������؃[����ɶC�.0x�}7(�]��͵�&�Z*T�7�c��W�뗀j����֧�#78��X��	2v�������*�z�p�oU\�V~q�5���DG������q�I��,F}��,�N�t�r�����S�M��֓� y���,�zCʽ*��	��� N�$<��X�=Ƨ�O�3E�16q��h�nŵm��[S)xm�-X"i^��1ۄ����G����sS��������`=+J�n��DC�V;o��L��r���L��24�>5����Vq|�	�t�0���ZM�ĦՋ�kz�b�\0}T\������B�UomWYc��P'�2�Iy�^8�����v�����ew�G�;�b�����:���P+�K�h�Vr��`-��r��3""}��s�S�SY{��M`��g��^9��b]��2N<���b��8�@����@%�$���p�$�G�{������u���|Q�Xf7O^�P�h�0gZ~
w�=6��"�7|��TVW�2G�ʌ�.���>S��v�3!�3=�D^�~��K��L��L�w�L�gTҊO�N�J��p_~k,e~�Wg �>������m�ʂ�ab	��|!6!C���k3Tm��5�(4�SZb�����E/ʗ'RS�� ��2��+�$0�-�TsK��� 4�`r�WJ�����9P/�+���x�R!G5e�e��\|�k��x>���Y~+#�"wՉ6Lql��f8V}�eԣ.���V[y0��d:��a��ט����>�Of�XO�����4�qL"����N��n.`�=������Ry˪ �a��O!/�]}�@WyյI&Ȣ.
���A=y�yT>��m�v6��[���w��],�G�໒ǺYٔ}9���~�,�e&��qA��o(��JƋ�J��؉i�c2iǬv�6}�����g��܌���JL��*V��0z~{���w4$�p��>#˶�j��~:��� ��'��L��B�_�l�M\m�\�eՙ�{ԅ�r��*��6ρ���6���}^ɜ��b��ʠ0��ȕ%m�|�a|�!�D�1i� X�Q��zD�vzZ
5��8��j0����A��S&����*h�
�:��YW{w˥¬�^l���h8�WMu�%���ʹ�I�{��e���S���J@ �^�ͬ=U �6�rb�I�q3zI�w(����Oes�O�ۜI�FcE�<��6?�_MY�-h���,%�5�)��>�;��B⼽�a� k�!��N�u�ڱ5��ÖJ�͋�!@��<�� ��:M�Z��sށ"K��������nT0��h�T�kk[U��$���<�
��f���s�h�Z~~X��b�"0&�����2"��?Hkh�tP�˅v5��.�$�wcC�����W��9b�F'd��~O+O^) �����YU�)̊�tLC�Xt8��&n���ن&�h%Y<:v��K ���^�ڊ p��:�F�#'1��b��#:tÍz]�U{LO-�)WcH������� �f���߯Y����i`�p-����cF�Q���e�t+ff�l��믆*� �p�Dp�Dwa��,�Z7�tN;sH�(LwƘ�@�D!0j܁G�?E��r�.�kB�[�sh43��8�9Έ�]{B���C1���n�<�%R��ǧ�OՐPqFG�(d}QU��51����c4*�X�cBq�W2x��Fh�=��74�rS��<��]��Ʌ��:T���<�t
�����N���"�D2�I�z`4r��j�g�e0�G�g�
�J��U=��֟��W��9������h�3�^���%��(����dLx|� C"ӂJ��P����$O�\�����$;kc����H>��#�
����iha16H��\gpAEkwn��/�?^Qky������>��2^��7?&�#��=� �S�v���>0Yܟ�)���(c���u�	�b���ӑ$ !�^�Bh|qȷ�B�=��8�͵^Ƹ�0=[Ug��,B��
D��'Ud���5��w�~j���W$��U�
����7k�M�o	��jc��H�2���+/ƈ0c���N?sI��2����I_�"��dY���r3�qN[%��B��E��<�݋g�����dܘ}�s�to/���;q���گ�5�O�q�0;���hupn�Yi9)��&FQ.ۦYO�2V�"T� a��"J�����Fq7j��B݂E�L����m+X���ap��E�1N��Z�3��p��?�z� ��P ��v�[b��ҏe�d4�:6gV�5=c,=��4/��8 �֑�7�#�p"l��|h͗ER�%z���v��@��8�FNm>���#ԚGx�3���(��@D\����0��$m:���3RA�8mFQ�h��{��/�ډ��U]����-�OG��.$�,�!�D׹�b!UKI�&��ʟ.*X	��<\*��i����L�ͧ����1�W$x.�V8���'����}�"ZyHj���,o�˴��P�#E%fA�|�q�wײc�Ƽfa�(V�d���K"�w���rQ�L��g�	�è:6"2�߄$x�&�_�V)�Va��';�����-+4=��MU�!�_���*�J��ݍ��i+����f ��#j��F�	 �2F��m0/+ar��2x��M���h�΢�:�h����/�6?u��o��������3E��Q;0k0��twbIT�ty&�1�*H�͚�=p#���7�C�u����~/��X�\�C������X˴c�}	�D5�G3�տ�%��m<J��b��n2�gIȇR u�X�qŠ3�2����0#{�W�� C	f��(����4o�eϧH�����+�n̈$�	�S˻�j��	��)��^���2�휱;.N�J���}X��\��̞�ߵ 8�������څ۵����ź��¸!ħA���.*�����f�^Z����y�	�sar�/|]T�L��]�.xe�^�T���DDUE�V�p�����ou�������ńmV�lU�]�t�̙��'ۺ~[{�zr��4�����PF1��I�/Ѡ����,y��f�f���ɷV Z�s&�l�6hE�!� ������#U.�J#��m��^K�� ��eN~L�tm�Z[T�"��>�� y��j��Ñ͙�20��67��Y��Qi&�N��,����(����m��e��n��+��4�6r;��8b0�����itƞ��F8��b����+M�5�Ӡ+����=��\;۴�.��l�[��E6c�'��p�W^'-��r-$���1[[M�4I�%(^Fk_�I���,�w]��*ۨ��q���C��1lS��� ��2�{��� 8 ��n���~��s��'}_����+��n�縥� jا�N�92ȕ���'���H�tK�k?o�[�k�B}��VX�?ī9�:�1�Ӂ�c2���dtE8�A��:<���A#�N�*�	9N���bꦹWRW�A�g�!K�h7w�>�`���t�Q_@k��t�"�iǀ����g�]�pQ���[��C���ַӆn���")-��9����&��*�O��'>.�Tk!��}���Xj����O��=v�C�RUN��)ڔ��̪g����oN��	���WK+=�����&��>jΆU�r-�<N�2
�='�H�r�f�#�E��À�m��D8O��ױ�z��#´?�fBܝa�3솫~D��.	�e��pE�;x�r-/�(��;�u���r���O;�*��-��;����G�;��%��[�?�&�S���^�MѤ|�%�E."Q�<���BW���-��s��n]�i>Zk�	�oƋO��Ĥ^+�����lҚ�h�ͮ�o�����%����(�Yo�gm�/o�Lk�b��׬�P�������������y��O�%~���+����<*���phio�d�9$�~X�H�G!�2v��PLx�>w����,�d�*��ُ��@$ykj1ﵺo@����7%Ri�K�Z-�[�_���Ź�Zo61w�wӥ��<�,t��V�r`���`�W�I���\Br#�1d��-*���_��P+S t��J�b4Dq�� DR�ކ��GX�y|]Z�Awrw�s�t����\����C��w��p���4㟠�É�^�l����li�oM��L�&�N�TGCK�R��!ŷ�RU��~�CW����B��P��zC��{e�yY笤���\@56)�ڐ��M�9�w-��o��^�C�6r>W1(����7�"��*��f" ����d�B�[��d, ����r�5��eE �]�֎#��0���*���,o=c�M�;��r���	:{f=���\��O�do�~+��MX}ik~B�(�:k�*tٮ�SPP3�BPZ�O_���P�.վ/ť��lݮ`Q�ӰJRA&#�����^��pw&1Q� ��ab�(�{����l�VyfR�D�{	Q-eۼp����.��&ߢ�D�>s�*�u�B%~ œ2eq6��擜� %�'��E��ȡ���.����3��]���j�x���$�϶&%�̉�)6��X��{=�� ������nk��]�15�sG�^�o�Pm��wtCiQ%^"Z���籝�8��C�WA.۵ .W��d�7K�Zr%�V�Y:���Ό���u�cN��7A�[`I�2��j���"�LNp�/1aȼ�5�4�dO #4��$:�|��c�?�mf��h�;_�t�c�\XDSDp����-��g���ٻq�B����yJx6,�#%s����t	�,\[P͕Tc'#+���A)�*�&�?�r���|5�M,��ߊ���}`*�m����y�1�� ��BL�7MqB�#��%��_#^�r�<M�:��|�`F83/`� ��h=���&0Ѫ4>hШc���Wn���F��X�����Z�io6����P��� ��87=���|�,��*�
�N�>���J[$�&��k�j4,ڋ��݆N���e�?�ؾ�Ϥ��p}��nJȣ���`�ik��%u4́E��ኊ�E�+��,�\V�`|K��^u���ς=6�ST$ۯɮ��[���WVE�[����ϟ/0�5�h/E���Q��m�!
�}��Z���#6���V�!)��2oFUa����o�t�ˡ/b����ܣ�G����[5�	������<�eP��x�ǳ쬟�*T���VO�G��z���UN��z�|ӹ��S�ŌK�@�Bʨ��=��t�H�[��iq��0�>M�r�L���g�*sN��,���j��Q��0p��!\�l�S��
������0Kp2ø��ǘ�ϪC�h���&�2����3��*����@uAD��ٺ]x������oc������h)g�*/_b�
��&` �--�M���&�0��3;���������U�.��A��u�wEW�k�͹�;¿��W�ױ�������b;���Xk��#�!M�]�n�r.��l�Qa���4՝#�M�x��^�/K^2qov��2�$�2=eX�"|	<�!c�Ȳ�0Z�y�ѩ����iQ'�d�Cov*�=n�[)`�QK�L𴤂��|P�1I�_�laF��L�����4����p��\r�e�uM&*{�];��ئK~�3�A�_̲�)�� ���D�!�Efl�oy~I�D�-ypDdl��:`�'3�����iXt��(AV������|O��R�����q�ɓx�BRNW�q��H����Zep�`���б��	�{�+��ob�r	&p���(s����z[�µ�w2�l�)o�.�������i0�����ȸZ��1�)�U)�_����l73BY-ʴ.9�M��g�S3�,��R�4��A����{���
Vk�I:�®WQ���6�x�L��CE���Y v�&��@������&[ѓс�ԡ:�6ھ���u �����(|cblo���5�+�2�i~���\꿙m���9d5��ԛW鰙��^XH2%�n���C���~��dzr��֖��;����~� ��	E�If-H���8 �/�h��(^��2��SB
�1����̅+RGy��4�z
���+�uq���zN�����OD{���u->����YU�Ǉ�ӾJ���-�H]3�k������S��Q,�n�����U;<��uW6B�'b5�͔t�R���gL&u`",spTn��~eI.�4�^۞�l��4i�T�%��\��	��ߗ��n��µ;%������Q��*�G���,uz�o��^{5P~>�4�O�Q�;�	�	E8bᅒ����m�r�����H�?j�H�ت\�^o�l��2�̟�@��vE�������@�b]u��Wu��s���(cq�B���Ѩ��l,?�%bk���3Լ�&�/ћE�S��ە��u3�ƫ�Z5�����T��W�'�>��`����Vگx!�9+�\�9��8
��1x{]5�XV�'?��I���<Ն��Jy��������k�Ue��:R��t~,���p	/(�>��8�i؎��U1XV�-ZkSE�S��V�{�����[�*e�1��x��K�/�G�m�9bĔQ�Vq&���_�(QSd��*������Q�-~R�q�Տ��C�'6�����
��Ѽ��c�>�� ���cM���c�AN���M��9�? ԏ<Ǐ�*�[F9��k~��֜�d��¯H�ûP��
�)�"s)a4��. 鉚�bk��ݤHmq�&9��%I���|�#�@&�qh�d^nܧF��V�B\�κ�00.f3����\�8Oy�fϣa*�z x������ �ӥ����` |�O��/a�i=	_�'�`��%#�C8&!�T�}@�6�ǉ_���z4U�B�dfYM��}y�~�q]���7�b�-{6��\v*UP˹���>�XU�i؀B����^�����t�Z!����턒��'�Oyu�e���¸�m����)�5Q�����#������j�bAF�aR��G�y��1h���O�W��]�Ϡ���r5�ԃ���E��n�����֤�ȼ�fv��O�Ԋ���o>k		<R �"��g&^;X2�|1����Mdha�Q�ҝ�E���pӻ��pv��{ep�&N�hz����[u���7�~�g)v�^�J�
q/&S�$��Ԁ�2#ޞ���bLEj��hŊ;wi�m�
xo3w' �9��jf�-�� ��.�'���RV�� ��yrvW���fܧM����(�N�:�]I�	0P�v�`�N�*,��Ҷ
r�7:d����{|n���꫺�ޗ�`~d�A��Q}E!����͐:��9�~	���Qӄ��SU~#���|��yh�	@�2������N����	W�qM�U��i��8�ϘW�l�{����FF���;�l�ҿ������h�&�G���z�M�r��z�=ۉ�_�����v�(}�����.�@7E�J��\O�������]\)N󁬷!ң��Z1y��4��%� ۳N�~�5��6������C�[��>���;��0&Hu��.���r��$��x������5���w .�N�#�&=��B�<���X&z-+_�{��b|�a�J�泈:��O%�,�C�V����	Rߺ�?AӴ�x�Do�����\a%�A�;�;�LS��4�_Y�4#�-`ZZ)�s: ��W�iӳ�Q簭G*N��?&��o�Y��meF�3�_�6t�UǦډ�ә��~��+����|�����h*ހ��ӂ�A�`>NJ��/�NHc���"�l������w9����u}�p�\�E_�)~�P��LQ5ۇ���!��(n�/�&���������v�FK���6��]�N~�L���E�'��#�<a�s� ��y��22i�э��ӹ����x,��y!VgC�䟚���I2Ly)����혚4_�-/�'ŵ3�NZ�ς�W�5�6���Y8�I������6�\�U?���<�R����Kj�od� ������>��4��O�p�T�s�	6~�
��t݋��8tX;�Y����|��܇��"m��G����i�^^
�� (�p�d´Dw��
;��b3{Ky�!pL�����{�J��H�i����B7@Hm�n�&/�<B���R�U������m������T.��g�as�B�u�.�-d� ��aF.��HD�U�|~�FE�u$�|������wCϓ�h-|�r���'�Ʋ����+àm,\e;cP��lȶ��,�1+��n �u:�֟z���[��,mxG�$؉����A�z��ŔdF3C!~��].?m<kP+�`�*d3���T4n ���XJ5
;VȪb��8�Ϩ���ƍ�&,������v$_���8�rS���w������P����EMN�\��P�0������|L��|5��O+������tYj���tHAR��+�76�>��-�z91���_��!��('��0�f�S��)� !��q�N�%p�%���{ ���yo���]�bs�F�lF�j ��8����v�(g�Qv�)�&!�⫲X���[��S韇�'������+6̔r��2��,��Iס��Ag�'��Ϋ�X�NG��/ほ�pȗ��w�f�'��ж�Q�'�+�І}ǻ�B_x��tB'�`e@�a4�r%z���˅h��p/^^���C�m�/�G�o\ހ ./��S �tֳ]M��;ї���}4j�(ml�#L��ï����Z��߆dk\s���hQ�4��X�|��x<^��
�Q�'�Q-�B��MQ��g(���Y�Z�R����p�2*|,���:#�U����$(��q6m�!]���z���.��	Z�#V�1{4;�"����> K�]�M��H>�RV����C"$���>_%��)��
2����9�3�3aXq�NңӁ/����W�N3��˷䵧�^o�췰t�go`e}�_Z�+7�X� 89	,�W%��(@��ƇsF�W���~�'��'�~6�9��M8¶ ��l�.p�^O@�G���׉[Zl�B�Cp�a�)v*����y|�BL��bzȪ�~��}U�sN�k6͑�2�x�uљO>i_����LdN����ᙇӒ�ؗw�/��hg�7��u��s�%��py�\YN�y1(�ٰ�YH�=-�WV�"�	������acN�U���6cc0j���vX#��$�����ɍ1�Յf������cH3��\n�0�g��*��ҫ��[�%���5��-U#b���h�Yc��B��;����N+Y�=�*O'�2I�	u-���Ձ���� �� ^�N����=.Ҩ�s@�+�o_u��Y���G:C,#"8��T�[t	,���cO��tK���o�-q�������@���n|~��ж(K�����@�g�ۅ�ТmHE9Z 'O���.�ylƷ��\B�X��3�T��!�$������oއm]a��t�8B8c�^�b�e���L`�!��u��=^qX&&I�6b7���F��Cm�BeXCk��8��~ 7�����ݮ.�rH,x���r�<t�A� sЍ;�!*�����m�u�Ŏ�{MJ��:�~�h�x��l�0|�ҳ �r�I����涨��=_����7�!���c�W�4CI��_�:-"�Q;Zc�,;��,3Y8�\�A}k�#93��0�p����Q�f�FV����b�9���7�T�Wr���ڎ�+�DG����bL�&��ݩ�	��&h[�NbPa�'���v�Bu��?�7yF$��	�I]����v%�Y\��6�:79� �C�V�q����',��.DY��ٝ�0ZQ"/U6��Pp��ϥ^�|�X��u���2_��H�
�:@j�5��p@��YySc1�'k��ر�ݱ(-`+
{��D;���=��1B��rl���}��{k!���l���:�T�/��+Zc�j�\���`q���̡��	fx�V��$�6�����8��ZgN�8ep>���L���h$c@�D`���}���$8�h�(��@o�2�(�_7�ܙ)t�	8>��
3�p�����c��<(�Z�$���gD]b���3�D@�Q 5��f��A�@2�����x,z#��Y0:۞�I�}�V��u�{�IqCb�~P`��8���0�K�4K^�c�!�>��Zw�l	���Z�7Ǩf�s:��t�B����Fw� |�w��)�W����N�"�UD�+u�< ���j]�֒�u��bM(����|L'�Ԗ�k�k�����и9.lq���I.�0�H�c��z�����:\��-4�HC�иsl���\�qL�|"��*<|�tR��dv:߈��lr`�o� ��CG�o�f��@fQ&1��q]��w_Q�s�c�L-���w���s�iO�x���p��C�J��;3Wܪ/ۨ����id��9L��}s4�Ϧ�͙�k�1�I68��`p�L{,�
�e���O����9>�����vR.��lo�w�=t� }����cFZ�@���%�T|�����x�.{�]H�J�d��Y`,cn��Dϰ;0׭(��-D^�HDO�0�7[���Y�1�H50��(�};-&��U��0����Ҽ�]>!�v�c�0T�*zj�m����ll�P��M�VN��6��4��䲒@1d�$�I�*7��|l���	�Վ����_`��yZn�xj���lB�m��n�^,{ �oQT~z��w>C�g�s
�w�r��ɡ��w/�?W,��<]K�s�7���a�R`�is;~ .�2B>�!�����,�{Vd��)И��P����X&dѽ���!��I�_�i��:���X�^��ɜB���F�J�gוp;5=q��7O�Z�pq��{\�~v�)�9�"ZKe���^��O�A	�1ӂ.w�`KLO3��1 �E�f܍��w>vW�D�L/N����]����E�Y��:_�CK^ !r�<������kł�����D[/P@�Y8�WN�D��*�̟����������i�$�iN��b,�`c�A�����{���K��������@����dG5�o�e�%zf0�1�#Ak� ?wG��
Jg�4�XE��q�)�[�%2Bu�����&Ț.0�ɑ`����M�[s�`�G*7�>?iF���,'go:U"�	��劐>�Z%?�R�9��Q)v~�?�K&�ҖJ���\	�b>Hm@���ߣ��#�$:��F6�-��צ�kj�>a�a�)t(�M�ʧv�pxul���XP��u�oPe0�/��Q>�E�$O*�R��3>9>�֜���f2�!����s%�a���7�$�'���hLR�; �F��HM�޹7��R��9v~v%�,o���J"��4���j�,������_w�I_�O��p���51�-���:&�L)�޶�=�+���H����#������%��7ρ��0�\f?�z3qT���ѳcf���DO�`�F_�iPQ��G�O�mv��?� �i���u[G�ؕ�
�w_
�����f"´����w��ON�P#1����x0P�Kټ�������U�2���2��˯����])y��;9R��y���b쵿��U�_]M]�D�c����ntn�z�,�������8ψ�S���c���O���bhZx�5��Z���+xc}j�Wሶ��X0M�.]�[s
]̚���iDk�Ћh��D����W�����f�j����"�:<��~ߢ���j�,Ȇ'A�Q@T��w�\�6��2ܖ�R"��c�t�b���3��S��ְso+�*�B����
y��Ζ�O�X�S��U�AO�'1@ULb9K)��]ՇUN��Nj
�'O��t�LJ��ǈ����Z(S�bi����{ux�yBD���tEˠJDE�▕-p����=ﳑC۔i휏c� ��P�כ`tx(�f8��l	EZ�f�wu��?��nׯ�0��m���}�۟u����N�B c0�\�\�X���ӵ���[abq�P �ƣ�Vo��!̔��sFw��.��-fOP�85�?'V��.�ff�^�����wK��<����#�]>Q�$僇�Ra��G�^��(Z��㤽��c��j����c�5ﻧ@YiG���$m�%���ƹc���`���%�b�KSui�i�/��	�Ƕs�6Vx�E�(��r���a�tŎO�竄,G�cG��Չʞ�P����T].�!FQ�Z�?��۟�v;�E��v)��NsN-R1�҅<P�x�Tt���:r�븃=J��1����6�a�f�x��Ұ���FÑe��Zq���`4���>�c��B�)Bm�Z�U�]մ�K��#)�78A$��eG�07p.�C�:#NQ�RZx�����<��֦�^�q��/�m[�)�>`��-�Dq�����h�>�b.*���l�X뾋=�����'St6r�"�RoSrpP)o'1ѯQ-��A�䞙�+*`nУӈ���O+�����dms�J��-�$��2����y�QE�t/B�&C��'�k4i���Bǘ9�4��AN���2���nH�ʕ���W������W�L�
~�
���-��`��$�C��ţ��ʮ�������Op��ŕة"0ɭS?�p���\u!�	.��ͻ�;����[!�/f����&ͦ	.ָK��6���wbEU��L�\���g@��C/��Oi��f24LF�,��L~�ޠ����������ouF�DO��4%;�傉Y�=�����L�/DM	�E��Z�'�"�_�g
DC�Ż���!���	����.���n�D3�+4Ps[5f���,�2�d��`�HȉӵQ�5�s� ������"�4�݆h���F��A?C�/���n��ʂΓYڪ���:�;�\�ۉ��<�,:tv����1K����4.����9m���<��K|2F��� ���ҕ�W>��߅�'7-fb��:���Q�ZV�&�����C3*Ζ�᝛���w��{�,A
�[�<�0�Q�}Pk������7�Y��H#]�6(lU�7p�Ll�s���"�ePόL9�g�����\l]�דrC��Q��L_�'dRLM�!$�2�O��E��*�8�L��As�8��q�u[�f�2$�kG�s%�BȗG���L\�ۊ�iLHS��ѡ]^�[��^t��B�ᆡ}�U+߲��O\���Qɹhf`����o�F��3jM�~���'i��~?A��/60a�Mn�){L��Ʀ��<�4�$�G�(.�}҃9Ѓf�%`�GR���{��C洡P�����63O�r��g�ȸ�5~Jq��4��^�lh������b����x�ֳ����Z82g0:�8�3'��y�c��x5��d5�Q�ț#�Z"��c� �Mfu||2�"�����oO%�i�V���4�I�� ��忼�Y�F�8_��'�3��D��y۷'�3���q�KD��4\F(� ���=�v�O�/*�Gf�VhpY�����c*v�kGNsd��{3�g"hO]D�pn����%}�9�5��z�|�ڷ�<cVX|r�������� |;]�eexߪ� ��@�[�e���O�;��}P�ӹt�\��ɻ�u�|y�L�MTʧ����h��7q>����XB�*Q) �)��\�O]^#�S[���}�d3�(��~�EWܼ�ID4�� �-J���H�s��yj�s�����K���{7R�b_�|�(�'���8��I1��	q���P�|F�E}���%]K��,�g�\�����W�H�b��7<����F���8n�vl��"Oj�V"[�P&����S��t�IJ��Q�X`�����VbK>����[T�����P��?�&���l3�:]MG�9�I���R&ҹ<��O�~�S��,!����d��C�6ê��e�^�d�]�Y���>���T���n�`E@`��X��������%>A}u�#�V��G�s��٘lc���	����pO��+����*�M��B,Tn$�G�we>�ާb��a��]�y�Ձ˰=w���Q]��FA"��һ�#�$��-*�����ҙ.74���k���**��qN�E�0�#O�9�VN3�Ní}�-��y~ !,�Q�������l��K�Wjp)����0�Omȏ���ߋ���L�l�IQ��a�bv�-��:�R2C�DS�C7BZ�F5%3I=�z�d�W,!�T$;�T�!!��ꘖi9!B��ƶbJ�GT�+:��ח����5̺l%���<�P4
�o�Lg
��ba[Û{����lK2vM	>�w8�'�t#���30��R�bE�@�Z�����e�ކ�"x�@��]��j@��Bz�9����*1��˨Ȓ��9�졀<B��"к^x�&�S�C�f��Ch)0�RKT�c�G|슧�/�3�.F��1�Ĭ����& x����2Y|%~^4i�t���Y*�/c�쨻2[GS>�ϣ6�4w%�@,��v��Ǭ�5����z�
D���YJпj���|L`[;s۩0,ŭ��)��Q*��'�C�3pL��ɬ��#�_+������K_:gݗ�j�U?XpgN.�����i;،\�pu�ӊ�,�՜�x�P�	ڟ$1�X�7��S��T,�3n�/aҩڭd��
aJ6�yj� B-£Yi��/�&�S:�$�p%	�@UG��*��7Dϑ2���7�J��B���w7���պ�-�"�=��#�/X-\[u(<�-\o�]���,;{O�@���FWP��0]�� Si���ȆT;�0�.�� ��>ʱeC'G-�tV$<r¿--^��@���B��1dR.Q��0����7�����L�-�x�: ��EMu`��c��Y��礍Y\r�6$�Z�S�$�Jbŉ�����Վʹr�q�'OBX��X���,���)e{Pq��z�<9Kz�Z�Q �9����R<�R�Un��[� >{O@%��S���**)�c�!����]B����X��l�|�O�	L������������'7�� "M��R7�x"?� A�]tx�>ozҚ_��!k	�C':e��x��f-KVrk�Ƞ��u:el��c#�!����&(��0�������y��ـ<�3�! ����h}e��W���:�B\��	xn���ӫ�C?�d�Oι�i��9��)��Ғ}��a-�
�"E�L���Y��(�����*&�ֈ~�+yQ$#\$z7qb�=���š�P�~z��Y�JPK���؈	-hw��Y��"2�vG1NsT
G/�a3@�uJ�6��.N��xvA�r�,?u�J�},r��'+УT��E@<�_Z��oѪ]�Vr����B�>~���~S �cJ?�uݢ��8�����Z�9/qOn�O5� �T�!�����XU9H[Pf3l6�o8���k�V�*��������:82�!/��fR��2Mf�����1-���k9�ݎ���`��&C����ʽ�p"^{�g�+n��{��$�$���[������(�LB�^��aʏ�n^Î�qEc�ϩ��	������xP��%��%�x�5L��jm\��h�R7h�S�4��]U�t!� �$;��O��r�{����)�����Qʇd~��ږ���s���ß"\��!#G���$�w��]1���o��q��⭰ѷ����8�u�˼�%�˰-٦0TX��M$�7��N�������kB4���9���:�G�������_,�)M�lI��7���=X��;��Y��
u��<'�k�R=���[ ���v�L��*�,�5d(rt���'v$(���&x�"57 �����[�72��]e�if�Z.:��X�t�e�S����&�v�z�(h��\��c�<N[�T�S�0w[C̆�����~(1��{E�|���!�$�d;D�Z���\����M %�rW�CwS����dʥ�t"P6���T�%�-R�~�� ��@�����=�$��s�fj�,���V�+�X������Q��mq�����!H3�|��#��e���?64���	")�s�K�B�j;��Y/eC_O��x��A��3v�Z�Z �+��"�^��$�iƮr�_}p9�j�L D��h�uZ4.�� ��#�k�����mj������z05r�*�����jǭ��dXe�*"ę�����G�]��9�I�_o��_yx���E�k,���MS�g�����(�N��7�?ȇ��0��.6\�E�ÞZu�jTS�JB/���UoP�G��Knp�t0�g��a,.���ZR"l1�Y�	��
�aZ�x�ؓ�~�e ��%U�����,�T�$���b�E<�b��U��'�1!�Č��?����^H�Z:Z��O5^��
v��9�v��ȭ�9�S�m��R���k#�o��æ���x��b��5漷����"0�
��w5�3.*�XN��%��I�|l`^�j�8�m�$r���(-�<��j��3s/3����^�83�L%���|LϷP9&R��Ȋ����a�Y
	������\� ^�.3	����������*��D�ňfu#tO࠽��!�LH~H���ܐX>P�Y�표���U$.���� hR��l������\����1��%|;���:0�wI�(_��f-Z�.����;��g��6c?�gMPv��E�ąP����@��5�Km#V��$Յ��Hc�����uȘ��� Ʊ����gE ‫ôyUo|G�ֆ�z%N%�^��С�|�@=cj�lH1M��� x�h���|(�7��!�/QN�L�I&?�duF���������Py�!#.�K0���?���9{66��n�	xe�;��̪��L��M��69:m���
|u�f.��H��������h5���J��ЭX��I$vs|���L��fN���͍���@��(ܣRw�σ����|�J}�I@)�a�h�G��x��~E�9bӛ�ފ>���S�h�@=�iUo���|�� ��')�VYOk*�h)Z?�v�f��K."�)U�}冈34��l|�Dӥ��#Q�u�/��C4�Zu�k8��v�VEw1m����~��5[ꡃн���u̫�^cbB7O5:n��e���Q�^P_�����"��;SpKh�{D���R5uZV]���SFW �`7�|����~�c-ӟM�% 1 B�ɮ~���T�kA��0��x�s3�Fj���y�W_�!���5��2{����`�.z�S� -��)⻤�OT��
��K.�Yu؂�;79��^�܆��DLw��T��ړ���0-��{�Zu�������Ͼ ���N�mJ�G6t�c�?�W�;b�9�1{����C��~�ww)+�[�x#�%�n��1���3%�D@o�f ܬң��3��{Gy=�F����Ɨf��έ��n��h�¨�����3�vڎT��8{��4iҦ�t#��
�z�)xp?�>�Y��]���t�s|p2�#F����͸'O9Š�{u/�V-����{�s�Cʏ� L���V\�)+E�ƈb�^�Ia���@B��>Z���QW��_���~ �邑I!�.��=�?���Xo�d�}� ���+�� 
�J�|�,�7⚒����>Ilg�m*Aj��ar��Ȿ�Rd<�N��*h���[�N�y����ۣ�մuà�Z'�]���q�{Z&S6��-��e�C���.[do*;���(7��?�}#��Q�τJ�!7X�q�w�/O���lK��]�����悢q�s�G�
��>B��{ah�e��?��+�gL����S���K�6��ZYb�����;�L�;�f�٭y0�Ɍ^aw�[T�~��,Ö��	����R^M����X��'|4O�����K�t�b���Fz�����#�@S�'����P6��1R��Xi�F�wϒ��ce`��(T+nj��B�'U�H7r��������R~!�~~�AӍC��P�E^�L���G�jR�����H����y�T��]z�9;�(t�s~���;�e�K�h��S ���1`°#ʤ=�]��d8Kw\؋���.���p����<B�n�5j����8�]gl��&�������$����u.�:��I���Z9ټ%��ڂ:�1�j�`Mc�9p1���tf���a��n��|�Z�E����O�NS��Ƈ�G<��p��4��g!�۱���ݙ�Z�e��>;$�)��� Ӎ�LK�c��ٓ�v�e�8h9�5��o;~���gX���LQ��9���n~�u��p/�E�o�l�>[^�"Yy|�Ʀd�i��
�}e�8@]<��L�#�j)���U��gBE�6y
��xQ�uF��,�����)�7���x����|�n�ǆ�������r#Й<�U2to��@��k_.�	S^;B�GE��A�8��H�M��W�)�F�ύ�ߗ�4�f�
�$�`.���#�f�(�$Q�����x�x�+��x��L8���G�f�vwcaaU��H�:�����	٢���u��7=��Pɛ�?�No¢����x�1;�"��e���a|�Q�S�'�o$?
*|5�y��1��	Ļ����_�"��l�J�4��
m��eN����cJ�	����H>Q!t��;��,o�b`�y�!�ࠅG�����g��9� ��q������p��3u�A�L6hd���Y�@��:U	a˨qqC�V�wƌ�c%[��#�����)Fo�MB���&X�& u�Z��~[9�/})ti��Y�r΍*��p�r��86�a�1���H܆�ev�y����S�4��ZVn����y'����jU����o�8rǉĲ�x�]��q�j%������I\�禐��ἀ ��:Ҵb�n��\>�\����s�������	�oe�2����Ssr�d�� &�1u*�u���/��/,��#�B���n�7�"g�+�^� 3�����$ꠜ|��i�;&�\X?�Y�G�Eژ����ЯbN+s��\��tX�&�$��4���sv�� V�T;���h\^���=#��x��N5�X�4J̏�q�
�����u�A�/r�ߺѵ��ܽ��azdq\(��_�|�b��M��-Xo�0ܫ�̆X�V�5��?V��"��haG��F7�H�L�\�|�U��ݟ�Z䎮WYk6]��� �?��'Zl̃,E�?��f\-V`Q��m1F�ȫ6,��㱗�d�s�>y1R��>.��]]Iw͆���?,�����A��PR�A
�S���:������v2��Ō%�.�f�(�{Z�*�:�2m�1 �n&�� �����	��ÇX{N��;�>O�v��\j7X��2<A�s)�qR��@3�^�����̓��ɔ)o+�!rU}U����Q���_��?*�w��O�f;nd6��`��E�PCF,B�B�йd�o���^�h+�v��(7��q�CI.��"kz��O#xFc��%ى����@��v�1f�G�h>�J��PpY6P�g	}��{����;��¼���puѵ��Gw�L�lX��M-�?�K��1ԐL?+��F"���m&��w�U\����x���q�?��GN�Q��3��c��e��I:	(j�"Sͅ���r�\9�:d79�2�ytu>� �5��Rw03��ZD�ֈ�����o�ɵ���I���|a¼�|��<�����sa��"ڬ)
}�� v?s|)�d���5F�OA.����Q�.�L����dp\��8��*;��M��zz��p��y�c�����=3b0W�39��O��Q_�P�˳I���i-���!�<����u�=>o��(WAU˟���N�q�������^9�aX���ʞ�������<������T�׊�0S���J������N�i�b�\y,���C.�B�%�8 �a_4����h����3:�􂲘�Sa��JB����Pby�(���)`����2?�{��k��@�Q���m�F������<�VQ5��U��@��@�m���9
9��w�rX�������pi�o?u!�eG�XK�n����vɉ��vkØJ������g�.�f�)r�#=���9��>
��������j7��@|���J�cg���V�\�J�Ѩ~杫n'�Q8��z��2{5�]��u�������1�%C��dU)�|��ra�]�Zc����[8���u#�7K"ŭ���ݯ�Q~���~��Ә�g~{(,@2&#:�؎q`�c� �&Hb�?��I��( j|
Oa�)7��f�Z�D�-]������֚3�:oӳ�߁�uY���E:#!�����xұTb���9�S�� ���*�p�;yW����4�Љ�قr����ݳ��_.��
{���B��L) (��x̑uvK�η���b�M6w�#<²N� sY�5���2E��5��}m�
oi���(?�N�B��32�q;��,�%�&�{B:�t\�i�;�{"W�����m��-��
��,_�5���"�G6�[��p�"�*o���7@��Dȋ�5����I���Z�T7W%"��
�+�l����A����q�!��5�6<��_�+u�]��3.:5̒q�M� y�`"u����*v&�}�����,�(Rv�>�LL�n�ϴ����7.�B� �U�&������NQ/X���%Б�G�ub�*[F^J�A	:�Oq\cE 
��8	��N��(421|���j���:5HfqS�I#�gH���K;�5���4%����A)��n G�,c�$y�y)�v��޷!�:�\Л���wn�f�f�:{�Xq󠧙��$2Ia�tes�@Z�_W@���bo׆'�,��_�fٴ��Ƀ��.I:�{ÕKG5y8L����rՃ�[���(��}¹j���<$�7��T�<l�Pn�B�B�.���]L�����K�h���索 Y���`Ģ�����V�՛�^����� dt�UJ��� 4�I$պ��ĕp�D�V�?5!'p�d��h��G���s��g��,����<��!Rۡ8`j,[%��v�|���f�^����C�/ް�:"�A�頽g�ąb��?����W0`�m��k�h�[4>G	�/�zڡ��l�u�B��&�u��2舴�)��K���3G��<?��1��V�z�N�;���� #h��Đ��(���k#�>4z�l5 [��G����@N�<�	39���9�=p�"��D�A�w��;|�>Ǵ*qwm|�BGx�G��C�@,kѷ��a���q;S�9�v��pMu�=*���4jha����l<�an%y�x���}�B��T>���MU1Z4S�^v��X9�L�q�_�o��?��4�3L��7��:pr^W��]�_�FĆ��#�=]�*ﴸN��*��4�N� =-��|�<�^C�vOZƱjԦ��w{e(�Tk����l�����a��wPLB��@�EcĘ9�15X�
�Fj��EZћ�|��0y�_V@u���jnA�vR]G.��P��IM��~ʳo� ~~��i.]���h�������v�^�*`�p��%Fj(rK�k���#[x�h��o���dЋ��4m/�M�K"��|O-�6�Ӱ]��&mg��02CI�V��+Y�%�a�uU~��wܗk'�y&�	����^ћ�GqN~IƓ�$�9/��Y<	 �o�	�I����lJ^����D�c-6冶V�<D�n��⏬ݙ��?n?X�V!*ϧ���>bD�����qԏ��)wN�߆�#{�;��|v걁:�%�?qƙ=q�;ٍ��jo�|:93�v�O�B�:#5�l�xw�p� 5:�0(cÃ�R�}~*����$��J����K��~����9��[<�ײ�jB���Q��*y�%
 ��E�� ����tF�}uH����q�D��N	�z%-���r��x�Ki���H��%A�<7��H!���}UKXy@VVm�E*�y�uc�+`KA� �0��ֻ�z�۬�S4wv�2�Q++�ēXT>�]H�1���3�-	�g;Ȥ4~���v��[j}�`�UTX�u�׉�.	]��w"d�_ʡE�l���E�P�y��"�IK
����T�W>�kr����6�'�R	w�Æ<��k�~�g^c�m�\Hh���e�V{w._�Ƴ�W�c����q �x�Ԃ
!���
=s�T���}gŪ�K��n��a�T��HV�y�$���7�w0Q����˒�g�\K2b����v7����	�<�#}t�`g��ë�N4��18��D���`�E��V��x�t�Գ#���Y��1[�z,��ᣨ�Y��	��}-'AiJA�Ճ�Y(�#]���!ުT�u��@�|�g��_�gc�,ڋ�9�q����?ٗ�8�t�vڬ%����|&; s��GX�z7Eja��9�8��{΃�[��]�"b��J���e��j���Q� ��+cՊd�Օ'�0g#�?{Oh��;T�E-��5��mcXI[���3����%	(@� �1"�wP�Ex�b�J��B�����a& �ض._|`kwNw3M�%����Ct��G���I�����t+�ˉ\$:|`��`�e���[s��8BAO��D@_f�g��H20�[C
r9{�m�=۰���1�~cޣ��p�rd�	q�T�����y����,3b��h�(P���ux����:���/��'�|����������}B���¯߇[�����X@hb�$.�y_�yS�%#��J�H�
�*ZF�~�4\���=E�Ȼf�1E�lǵ�{%�]#��_���9�]�O����(}4�\�\��p�?�	)�К�^�^!0��x�,�
Ui�8Ȥf�K�L��+� 3�������w*�b���M*�j��7oK�NM��T���ѧL-M��y�l�4;�^�:�A9��G�L��ܯ��&O�����Ӧ��=怞�{�_�4�q�Y���as�j1���96��H4�*g�	���ؕ�+�)�/���1�N��jƠ
ˊ"������{�\p��9b�EQu�$�o���s$����q7Ҫ�
��ݷBӒUw���W_��X^`TxlP���cƙ!ZB�>w�b�[���U�K�H��i�pO�q�X1G	(�Y-����D9����Ww%Ƒ�Yڀ�d���)�oFX�8Y6A@Y��:�ے����َgz�R���ka,�L��қ�`�P�Ob��̳1D��ш]����D���?�uw�lx��d,�[��ԶUCG��R5���X*09K�}��lfs0���1:�>W8�.�N�������������(���$<:�;+�#�&(��5��3."ϠZ�Q-�U�7�:�q�����3�zo�̀EHC[��p�ݹ����8�U�O%V�����d_6��	�Oծ�{� �h�b{����l��V�@�b�񆂾��	�W�N}�JΪΥ?�	k����[oo9 ͗�_L֭>=ϸ�e�q��P�(��@���Q]Āb�,Y�#*��Y�ud�:k�cF	�#��vj�����"�#%��DC֏d��t�@�U��t}��KD���O�XCKj��y���q'���X��I��;�Ev����_&����[EVԎ���$j�- ��Yn%g��6��b�*��~��D��3��2"�U��7%:�\{�P7�%"}!�$��[��7HګxS��s]2H|�%��3��ptY��Kt[	�BV�����䋲f�*����@�3��"jG�=���O��Dj�7�����Pd3��ڴ}����ͷ�j���t좓o,��������JĜf���|�7�]᧥Q� ��>ꁣH���e�3	y����YX B��Kk�w�6,t�(�Leo�4N�S��o�Dt��R����I���nŲ�4^��g�o��I�T��S������:�c��g����/)�4x���6	��e0�~�2f�{O�1˅hN���d���&::��
7��x�bM���LJ�����3%����s8�/��a��Rs�a:�i�ܛ\�q2N���+��K��UN���2�sNQp)�i%��a�d.���V�y���YGB�>n���bU��	�k������l�ݨ���q���/���7��iz�$v�f<�37��l�N��Š�4����P��ޘ�x�ŗ4BԮ�|��������!����K�n����L��O�AچJt�o�U۾ %)X�\����,ez���x��@����:Lv�#�ݺ��h.� :�Q`�tiM�����?�'�VFb<8����(�X������ґ�2ֱ<�`s��Cj`IB�zq �%�p�̈V�l�a�/qgI�nj�!���PQG����e��S��UW`�q}jVƕ��*R"�z�o��g���$8��'����/Mm���� ��Pc�`�/�՛���0�Ҽl�%[����XU�ؚ�T�>�VH�Wm�\�w�8B�D|�
�w�{�H"�z�4��3Wb�d�H=x�}Ց�Y�X��8& Ǐ�]8Lu����4�8돰`�8�*�u��@��ϘᝢM�2ܮ`�m�8�TatO�-[��	N��1��Uj�&R2��Il��}*#�Y$�rq�ްA`B/��A�TkǺ����*4P��M�@��שֳ��"u��携�ٰ���0�cz��^�^��];zA�D�}��j.j/N;�P�*����5�ނ�2:��]�{�f���CA�v��YHy�\g8���sX�h����R�X :��32SFO�^����ӎ�f��-���!�ԯm��"&��c���pi�6�v0H�pޣ�{�~�}A�8��"�x1��M�$ͫw��U�̤�7~��� xn��'�el@2��v��M��	\(�~AF��:N(����	9��w�W�&MY��.�2�@�ͽ��G=ś��G�O��?U��1µ]�w�CH�[{�R����+E��E�L���3�ڐ���@ud޳�:���Gl��N��l3ox����.����'�P��-��y���g��L{ҧ|9��=ar�(��`�1_�[=�+��i�>^�3@�A5l|r�=yݴ����~��3���8�w�+1�BL�Q��r�E3�쌿�[�F��Y�]�=�����P�K�U�n��DeD��i����^�:Ƌ�\KX�p�g2�u��C��X=}�jw��(�?St5(��LQ(P4�w=Iq��.j���V	� 2�#�W{��v�{�������v��e�݉�4�4^�0���bs�A��KL���%?���oTY�	�p��������~9��T�	�/N=��8L�o��>�;{�!�Ae�m�Z�3��;��ۢş������,Lm��Qiv<R���MB�ʉ,μӦ�cF�X%W� 1��$��hƘ����G��B�fLb�R�]o���=?�/�Lu������:��~��i���L�+�(����٧�@?h�Q�x�Wx�|e�%�|�\����� ���ct�^5�W�>���ڌ�u�f�d<>��<��V�+�beX��ɶ�Ma�����N��I��-��Q�N�C��o�z�f !���!�0�S0���q���ZA�*�������������S�����]�9��1��7V����T ��Y�J���@�������PE��9�V2�̝�����hF��y��������8�j�4?�m�J7�%���sx�D?x&D��d:8\�
����䡠-:��c%����x��F�_�G��� �Y
���ֿ'x�i �(9���9y�"නH>�l��BD��~�}Զ�'�I� �<�:��v2�B�m���5^���
����k��'��ڡ�r�;��*���h�!,ܩ�Z�A(�n���j��r��C/l��<�k򨙪���	Q��}'���2 ���_"�ߥ`M���ϯ;��e�}��4"���?�����Pb�d���~k^ܝ��8���n��"r]i�W�S���N�1�[1nh���y��G\rn.�'�x.ħ�D3�d�@����&�8�+;��n:-l��hzh�K(
^���ߛ��;f��*.�(Z$!�>:y�+���¶KA�"�m,��
.U�U�
5c�w���̫��~iBW,Z�����B�M�0�.����^�~'3kZ����s���}�I{�|+W
{�x����J��X�k���0��삺;�k��3ȫO'��2$y{�.�(�$�G!���[��S�����k�LG�%�N�/�I��֪.�$�by�,`%�wW!ɻ�~�}�N��>|�9��~�#�������hO�{��a����S����ܨ�<Clk���?��7Zt�[AB�Kb��"��K�U��2#�E��6�[�Y�>Z�[O��d4a�bzN{������}r��j�~ǋ>M���v>`��&6�]��ƲZ����=]R���O��W������7��E��8�z֩;��p��/�9g' �i��F^�A��P�����>�Վ6����z�m�s���� k��%Wg��Ȗ(��mC�!�B��V+b�=��P&��H�:]7L�n��y��������g�=��rS��ŵ�!�3��C���{�k��4;|�2\}IiHڞ[�ً&�T�����:/�V���aes����#^�y�V�f�?^0/RF<�$��;��O�顥�a�Z?3�����>A��cՍ�o3]���eY�ٛ����3�UL�B�C��C���r���z���h�;�K��@-j�ra�M��G&��m�ZrNYP޶��4"k�ZmE�1å�1�(�J	[�5f0p��;�i��Tʔ�<=<~��av��L^���.d1����/��vka���H�,��Be<#�&��m"f�쇧R�͌ �KF��$%+������8�?C'�ڍ(ē�<�̷J��)�RZCv�4��<v��"��t�.���U��K
�ZV���-u�h�s��."����AQg�N4�X\����̿�����Z�y��"see�v�턳�/�Q�P�뼋��4$���S���]��qf)�R�1nҔ������Ѧ��O'�F��Q�r:浚~Z�ö.Z��#K�L��J4$��i�A�Sq�)_�uG;.�5�7ʺ2�⃚2S�8֊d�An>��P��ڞ㲔��9_b��b���JM{k����(�}��
S��Fb7�6S<xT[og��~C�"�����[:��4�'��%�a��L�H�c~'*ds�H�~�N�L�\GZK�,����^n�C�DW��'0��:I�V�R���L��$KYk_��6�v��k�n ����5L{UF�w��ivmF"�ۮB�.s�-m�8_��1��l�95�;6=؄�ޒ�#�Þco���7�%�//9+�V��#���K�����k>^6^X3r�C�S��9���M�O;�+x���Զ4vY!�&t$�R����]x�mUx��p���d�)�|��_��9�+k���R��q��� �������{���a�S���h���V�h�ٌ뿊�?S��_�C�@�4;�ۑ�wemF�~�Y�������2S�w1�D������Hڎ�ҝ���_Io鿰��B�l�,�2�Z�M�R�-L���H�F�q���ذvLv�:���K�NB焚VFIV��9
^^���l�O�3]��/��;4I�Olߑ��Ѵ?��Qo��"ϓ�m�D����6���� ���l��a�ShZ?�bc���|�c�mLmwQ,��QN�Pb�cF����c��zۗ�����9&Z��+f+��K��^MyN����
	������w�W)6�z1X��s�g�)"[B����]H1=�ca�]e��(?LߕZY�}-���ӵo `W�5���^�y�^�'�Zw$��8�5����W=�J8��7��������!�	a=U#9����ۮw� QS�I|0���x�.	��0�.�;��Q�)b�("�e��|D�7�+3|����o��&�=Qzp3˩5�Og%�{�Pf��X�9�O���g����zz@�_��Ci}��0�*#FHt�L��G�t��^��xsfsO�J�k)���O\M�a�u(�!11���D��[���}�#�����6�!'O���X9�\ae���Ϝ'�R���u�.�
}�D��
P���U�t)0�Rq��2D��K��PN1�	���G1jboUIc?s�x����"(m0�����uY$���]��x�A�a�ԙ�~[P�A5^^:bL��+�N�r�ĉ7��?e�{v$�r������s��V�5�?|ֹ9��Q��)�(EĬ���`���>�жKA�ڄz�b��^�M�#8%z����@�<l����|��{��q�1F by3}'?$i2��#��ńs(�]�󽄐��ǲ��gj���^��Aj��r���	��Yy��G��hٴxZj��.\[m'���S0�=E��#��;���nP��/�3���`�<��_|t���P���)�}n�%W�CP[/G���eP�5�)7��SM�?�ƮT��ǡM*5���&���5�8�!R��,��qʀ��䀄�S��C���uā.�i��
��ң:G-<bJ�Rr�"l�r�{�ھ��FD��t����џ\<�q�{�y;��Aw��Zz�u���X�)������B���TLG$_��?t>�/�>������7�da[5폴O�y�!�?�N�C�LU�u��#��E�q"�������Dw�����]��x�:�%|s/3='�`��q���\ɹ:=����U)q�/Ā���;�j�.�f��^:*��l���gŠ¦�8��]���k���G�`�Ͽ��ǳ�&޸8�U�a�<��s�,�	�X���J�רV�lN�*����cH'A&+o�aC�6	�k;a�P�b�H��Ԁ�#��nu�-�.*S4l�X�X�q�&T5���V��`F�pr�:���x=�ʱ�'&i�	ly��.���]7���/1����)��FUY`pò����ҟ�{V�b��!��o�-���U֎Z�kjv��67W�q]ѣ�����^_a]�Z6�#�C�3�0���Ƈ�'����a����{X�ҁKFH{��6<�7}�tC)�J����jF�gu"��O��5����y`F��[M,���8!�)�	�ǘ~����ۦ#SRSj��Y�þ	ƞ�� �w2gW�~�T@�B���3�F�)epqWF�GDX��	��T��t�Z�P&�g�������nͥ�n�+�ҽ�����ٷ��p���ʛW&k�/'@H�]�����U2�P��5�X�%Z�4��m=";��xf_�kt�Qa(}��<[��#��{�	r�v���� �uNe7���ʃ���ƅ�t��B�Jӹڛ�>�+��;�@�C;��C��vJ	V�7�>�t�*|X�B2�)Y�С���}���z�.���}D<��*��,k>����y�^0~n�8�`�}��I�^���ș9V}SR蟶1�����|�d�T �����eCa{-�Xʔ���[�^�s�7f���SӦ�1w@�}�e!~w�8��`�i�[��=�h3]�w�AW�j�������H���`�dp�<'�P�(�������Xѝ�,
=K�'������%�}�ԃ��������I�	�08#��c����h�,z�7��Ή�u���A�\(��k���U�����cd��*Ѫ_zR|SP�vg K���2I,��L?Tw11[�����5���3�i?{Ja�K�QC���������@���c4�Q��S�/��lu�I���+:�$<8�0�H'#����ns�-�'�g��H���bnu#��W�������z�t ^�I�v�P>�ID�'���đ>�F��w[9�d�\ɗ��7�5���ZS��ؕ����f�1u���r���	��d�����6LQ,���$CKSĎw@�_tL2~7�s��^�ȿ7���?>���RMi�O1Fp���0O��ŢΌlda뭨*��WW��"���(���]V�ո� K�ԕZD�3�A�e�����F%(>|��&���l��V���.K��K���@�{X�/�ȀypsL�s���T������ޟ{���p9n�I����T���sM�`
���==�JӺ�ӫ{�zRb��yD�~�����J=�i�)��o�3 ��ua�\�2,�F�ĉOe �{�8+�������x߲s/�/�����mq��/o^F3�b�iUtW��2���dy&��+�D�mP�(̣�p]�D��+2_B�A�p����3P�Tw��02�&��i���dx`�~�&�r�M*g:�"�t��c��J�1���\J22�-܏	Z0kI�[�V�@n8D�&�>X�C�X�v�w{�&E��}���IIW�p��$s+&�!BQKA�>�-ů�/�V�V
�{$�߼�G@��`ˎ R�m[-��"�1#	؅�U�b��Y�:�aA�~�򬲶8"ܷ��G��3$�����!}cf��h���b�	�+ 0�x8/�D+}ɵ�v�y��#�&���7r%�#X�L��i�q��M����C��!tc`� �i8�M@�ֵ�9��a�q�qçr�f;M
㹱��ru�%P)���	��)��>��R""�7t*f�KAs�%�l�)|� `����y;���|}�^���k�0�I�O�f.ӈ�,����7�w���.|�X���/{�3yEs���;�ȳ�mN�nm�ܝ�;�8q�ϨD��Q���\���=IV˶���{/rB����D�=G�'�5�F1���[��(m��ݢ��?�3�y�aA��1.MTQVH�7u�g���C�. Ɍ�;@CPbw��O�aLu�+ת�5U�(P�c�e��-DT; "��
��v��b�J6�`�'�zy .W�9���wgZ���;�ÿ�V�M��ܻ<��ཁ�R�Yr��s�8oï�(|�z��q�.p�#$Cǭ�h�� w�+��b��	�Y��[z�6���ͯ��8]�{������3�v�����N_�u��ә'\�\����� �����?C�"�1�fDW>PĚj�Ա��<ң'_P�L����t�CV�ڌ���|�[>��Ac�{��/�W�`����E8�>����EvOg��Z���eJ�Lp�А��UT����Ƀ���"�����~��(<�� �}�v������Lh>_Y8,��.�(�܏�b��H�R� +��+�A�I5;:��Q�m�ǹ���a��g�!w��>Z�uGĖ�2����u%z �0�H4�������X{�q+���^y%���o�R ��H��%9�����H�!镱J̅M桇�3�#T�9b6_��P��n����"^̶3&�a���ޗZĞ~LΔ���wm�rE�2wi;�5A��k潵�F?���(HJ��>3r&�Oh�7����p�h7;ZHj����d�[O*��40��7i�6�?���>��^i>,%�P) �)�I+��WLu�&޷�~^z|P/�bRtՅ��v������J	�v�v$k��E9i��9J̳�q/.xF��s)4�E
A}��<Dp=#�_�R��8��tB�9֛�=h��bC/�w@��?��$
�ȧ2�s�������l�[|d|Y�H-�����ٕ��G\��z����X�d7��ώ�؉����+�t6�m�?\�P��"�����0�N�L����;�Ҵ,h~�r��{�� ���l�I[u~$pW�E�a\��'�����R���.%?fv�o<x8�[��s9 ���f1#ib�禲;|P��Τ�>��	,uE� |����#��c5~����_vP[OX-_i�O5K�Gl��%j#��湍E���L0	1ʪ�9���6E�V䢈������P�/��k��'^�2��\He@6)�:���^�`��MZ��:>3`��J�ao�
�el�k:���=��$�.u%Y�P�"&@/ܳ+Nuf����Qϴ�ou�m��u��l���~y=��	�V�H��hL��*6˕������m�p��>Lx������CKBx�s��������n�G���1䴼hp<���8ܾy({7�+����aW��9��n����Hn}H�K�tu�K6K�ɸ�/S��t(nZհ�W8��ԋDM��w��ĭ��%D�Rp�Í�N�ȀG�k|b~'-sFc��po�b�x�j��-�)��&�ð���pf��� E!'�P2+�xUĽ�'>3P�K�@�= #�5��co8�i�W)��k��)��ht&�� ��%���t��c7��[&��br�r}QB�n*�ffD Q�I��R��D��yqZ�_�o��z���[Z��&����?� QP�e�+Sq5���n�kt��b�T���t���"=t��\\�
ɤ$H��k�*��I���}���w�,/��u�Nv��%��|�gp�(d��'�Ȉ����r�8�	���!%���֌".A��s��wF�C\��L_���;��o�vʼ(
1K\Qi�I﹥�j����U|v���誦h�J�c�\��j%F}� �B���*^���ďT���I����F��A�����E��3k�P�rJ������e���baD<rmv�yb�؅��Wڌ6��Ҥj1oϊ~���>��_`9�C(�����!RO� ����	1m�SF>�I���o�����6���o಄�kpaBF@�5����\7�i��k��B��VƏ}�Uj���z�U���7�^�|f�<~�l�	 CV8��#������ N�c��Co_�٨�)f$��`E�Bj�b�t؅gn� �$� ���']�����@���>���Hg��KG�I^D��1:>��@�p�ސh��@%�ᫍ��ρw���>��n�^�� �\��/�E�$�3�/~�2����LD�>|�S��.T�LK�໣��ǒ��^�� �A���\XF?���5u:wdM����qK��"�2[s6E�$���H�s[Ŗra"�T.�#�,/a��i3����ET|]$3�E����;�W}Ѕ��E�_~kj9��w�|#K<����6w&�����l�%���1��[b���GD0H�B���`�3゛�(��	<zr�wD�LОzF�(D]pΓ��lrq��u^���+q�'�L*[��-Q�����yz/FҖ���[�U�(k�Q1U-�?M���4�Ŗ�4���+�sΛ��M��_~C��f�P7YG�ˀ�1!��_�C<��LMrfc �!At��Os��G��	A�R�U?�ćS��H����=��T�����.ʔ��n/tǻV��te�U�Ʒ?���G�T\�ku�D��c7�&��&��YG$"}"h�R���0�z�<?E�\��Е��08���x��"����6�,�i����.!�o�[@6�� Z�!'gja� F.�Hp��D@�A�V����+�au�CF2��7�7�۩#�N.o�8m�t�&���m5���x���{�����~p�G���8{ՋXbAM�.�rem#/LF��KY��qF�,ZK5�5�� �΃mϾ�@���`��d�t2����r둜dR5e�1F��/e�����f0לLj+��K:��W"'�)+���Q`n�dQ*.����FT��]7gY�����}Z�`�:�������Q	_?�G������z�RII#5���k W��1�3�J F�Ja˼�g	�!Uo��IW,�O1F�nH���u���+�
���Wݸ�9�@@I�.�>C�lW1���NXS����	��F"V �:R�۱~0�7��[hv��L$����ߗ��:,�Kn��X���l%��S<pI�;���r;�9pY�x+[�ӑ�b�ɜ�#�W��/Ϣd|˸&`m��>V*�`�:j2�sp��7�ji?v�em5Ə��!J�f��m*�(A��Ȓ���
뙄度��c��#�Y�k9yFũ>\m4hW�gn�;��Mѣ�R�0?+`��^�|�#z�J&6����U?K&�Q=6��> /�F��Wr�?��f��V|���v�ǚwAux'^/��ܨ��8�Km�=�~�I!���6�~�tF=J��/���{��,Jw�>��o;2�/#�3dp}C$��Y�M���L"u��ƍ^;�I�F0���,��o5ʥ�x 2g�ugoԲm�cg��]�u=v����5�Ƕ��5�����Db��~y'��61�FMVbhq��C�ѱ���N]�$P@��SG�o��)b��vJ��:�@5�����pFy8�$F�C�+����lv0�r[_G�Әh�/���������İ���"�:v8���(�'z�j��R4�r�a !�௦���i��rPcAs(����Y8�X4lna*���@���=�HC�p~L�qCe��I>d�ni˙�:i�d�F�C��nWF�r��Y���0��T�'����'�g�u��m���z�[fi��dTw�uH3���7��]���A�������<Ɇ�|�9�r_���.l��Ǘ������;�4��S�J"0����=�Hf�a#4�л��!U�5�/2+����;s�\�Ŷ$�<%�?�F�5��~2���#��*�>�l��8�:�2/u�H"�G���j�&s�U1��
�N��_s�w�-4_=�s���["],��oZ��k�g����YWw�oc72jlǃɫ�e�8�cx���YH{o?��l��Bs�;�G~�Q�p,�PX�sSH�%J�h�C��̓���|�u_`�B�=/�8�^n��%ԧ@���F�j�;Q|#	Ny���|��U�.�5�l���L�ť��#��]�I�-����ǒ��w������{��J(��6�|��\ʦ(D�)�)� ̵�a�?��g/�,#U�9c��#T��_�ޭL�t~d��m�?�.��.��\�'V�����v	x�����N\�p\���uƦ���CaYF�V5`�6G��4�7�Td�j��*�-+E���\��!�M�q�������s��0����b
����U?�Z�?�c�/0����;�D�b:���/I$����q����IL�K� M�!ɕ��"���-ZsX��`�rUfAg3hL�����8q��u<��ZWP� �i�b��
�1�E%�,�Ѽk/yr{!L6j#1rء#1��*9�f�?�J�0�����[rYn1�/(�}j(�B��+�w���f��9���NDj���3�\�a����ʂ�N1�Ι�۹u���E�2`뻭��Z<�oh���'VW�ߞ�`ʌi}���sim=��>!2ݮ;BE� 4��u��i�0�����a����;K�4����$�	#?|K�W*L��OZW\��X؊��g��"�:;�:4'R�5�E�6�.Hq}z��h�3,5��������O��ee�����i�������i���k5���q�lѭk�(šV�&�e���"&_�FR����h2�fQj=�:�=���h��T� ̃���e7�yNB�'�,[:�<��X�ȍއ`>�{ޜ;��fz1�����M;U,y�����=��p/�er��I6k�&�>	����	6�Ano���_�/�����+6-��L��R\:,���!��T��UO$#�DY*C^�&�$"�4$��覢0 �����M�&C����u��E��}�M���|�)=FF,����z_'�ΰu���=�#� ��K�.��g-g��1��@�.���WWv���]?�V��)��y��x)���樦�!�{}�3;1����/�ɾ�["����Tn�97P���m�{��&YN���Z�	 o2���V�<�_�$��ln�4�p��`L�j-�x:���??�K����Q[C�?�9Kå��J��䮴�OQ�	/�U�Qi��B4��q�o�!۔��^�t�V5��}	��ݱY"���M���3'�0VeG�X�Fr:m�呒���? ��oK(��X�)�+�H	%a��^��Q�*&t2q�ZC��;��q_0�����e�j�W�O�_�"oH���oJ O�W=J��`�>4�ߤ�^i���Kf��,��u���m/_�Qx����[<C_�o�c ���}���x����ǾJ�V�(����-o���"*t�\�804F�;!��[��f���f�G�K�6hj��?�aa#�?V�*A�r�n���^<���մ|�*!}�,�%�78���jM���ɉ���M�������߽�4	�ԯ�:�t�wz|}�4�&\5F��9��~�4�u�Q��_J1��OWf�w��c���f��e��#(�!��E���'O�za����Ϩ�)B�����ҧ�R^�P_���9���30�x��	���r��1|�r�O�:�!~٫��S������q_6w�iw 6����r��������7s� �l��5����`~����(n�`@��sI��̧�&���I�����-5|?���s��"��H���y�8���Tz��NE�l~���ig6�=��Wt��nY��$Gd��r�@}���$4�m��0u��m���v<�t#�e7�f0�-�Zz����!{,��~������%-�@H���?��	�X�����s`��ZY�_b�r����gq�l=<��Я�l����׽d~���.C��!�wP��nIô�<�7D��k�G��R��|�P��.��>��}4��-�棼�U���pk~ʖ6�D{�A��V8(^����gD�B��\n ���/}��͘�>��?���ŝS!�uw�l?�Ia��ʚ0a,,�Z��ϊ��o#�=r�ޜ��s\� hd&|N ���D�U9r<|p��M
[��R�V�So/�@+�������Q�{����,��H&��~宪�k%ޯ6�=^K�T{�cgC7䅍����n��=��"�s_�V$Kk(*	��x��̺т�Nd⦖i�+P��m'-9. u~�^�ӶP_���s��,��VZ+�E��B���NWĞ����Gf�)A�Z�(|U$L��y�����K�F8�}	>��>���������a4�-�v��((�����G��KPݵR��(mҀޤ�C=������Ϲ���APR0��X��T�#X�yp<�*�����Pz��]�)du��(t�KC�M��	_���ԩ��Ђ���df�n��ET��[/�<� [/[đ����p�ʇ_���D�����ܥ�} �a���h�G\Yw�2�|�Ca����h��
�T���H�▾؎Mm��!�n�������v.S�/�&� Т��3R��o����|���!��O�Bh:*t�/v��!�⭞y�1�;����r53�K�x���f[Q���I1��9d"�in<���k3ޛL�>�o�9�����Kb�/�t�2����
���i�ҕ���i19��2	7�k/�)��VE���çگ���N���t�D=qHn[F��,��2�9����S;Y�I���يq�Ş�4��֐�j����=�)5Y����>n�?�܌�D@��t��6��zޯ1� w@^�p�!��c?�ռ�t�qKpI��5#�}�����|J6���7)29���9�=�!SA�)p�f�Jȵ�W0�`�+.|��$�H �$�IJ�0z�Ed��J���ȞRD����@W'X|_�Z���_��f��O�s\����Zt�{a~ L��a\bM`��_�#�Ҥ��/ 9R8�ݵƏ
"!k��="	\�9�aT����ʦ��W�	\�J��1�㙦47���|� ����y#� �� ��7�A�>��&!C=�%q�	�}.�@_?�� ��'�ކ��SIC�T������y�o,E��c8~w���h�����AA������ʠrv��(=���;Kߌ7����)%��gG��/��@��3��])}���s�<x3x��?�9�fhm
�G�ټĒa3���¸������g�����J�Vz����F�^fp�{2V��`H���z�LN�h/��Y\��qe\�����z�S�xSu�D7�������@�o1�����N�\��G����{��V�@���YسP��X$iPHB���]u!��z���M�K��	#�Z%��a@Ay%>Ċ��3ۼ���y�����3��ME<�&Ph�?E}��`Z�%g�e���9łV�.�a��M�H �-̹�S��ɝ��XS��y�NL�*�]׏�s<��C�1��� k�xsζ�D;����+�����Y�\��8�WȑFy�Zd�l�G-��p�U(�J��L��k��iz��_'-"6i x�-�T_�f���S�(1�D;��ݸo8!,�zW�"��W��
���Ɇ��ƽw�
�+���_�Ŭ����<������ǈ7g���2�Ƙ�]����W�F!-���MMɴ�,	*�;�E��iT�~����.k��&��	�OQ$8���β�|��ӵ�d=#��?�����>���d�vW�pip �	���.��&�:x0��֫�EoZnh����g�G�Z���ޝ����	�5����_1�r���1��Vg"]��O����[�-�$�z�D�,�vÛ�6Ç�:8�:�:���a�lB�*V$�MD�uP�N��l��2@*�fA��E�/��3�g	�_���՟F+c�ȷ=�|M�Y5 {x��/UJ��$eM2�J�M�z�V��d�$ʶR�O��z�V������9���,�� o����J�l��p��R"Srul���W���O<״L�:f��ǳ�	�����`�rI�����#�ʖ���������1����N%S>t�	��3��U�%��|�l���d�v �C�bo͔��Ƨ��V���UGγc��FC:Jޣ,m��1*��x�"��kd/��&ƽ��	�ؾ�I�"+�<`87���z�.�%�B�5O�I�P�ش��{�����]�y&we�QSQ�j�W@�~�@S�̋:�?�[� ���
�F~ɳ���5�DE�ǅ't>�v䔿`�G�u��"��I�;��6�3d~?�R�s�F��zB����4�#&N^)���2�t�C�����$�5��
7�<�/��s��.&J�@��_,W�%��f�T^.��j�z�`M��^u�U���#n	�Z.���+:�<�W��<[�dq�s���8(J�~{pA��r�I(١W��gބ�"�=@��e}Օ���D���e3{|�-���� ��"� D�;�K2Ŭ`�spa�QF��M�3�q�W\ V�$F>�i�C�}d�t=wRyvJ�ZSC2�"���`C�����v	���-��k��%�\HF&&����)E0�QT���O��}Բ�TPg��Aboq7�D"��R4�M��Z��b�is��h>��>P����Z��<�u�pۅ5q�\������?�ԁ�	N�"6��"���<w���N�\�߭��-i$w�$q��'󠱵�^TĘ
5&���k�8jW����/n�)�6
���sK��'�jS��.a!N�I(�9�=�ד'}@�>6���8�~��V���ZGvt��S�Oz��kTa�yڈhcX���(]�e����~9�ig|g�Z��w��9mR�����عQm� ��c�XL�!\�S�	�8�7��1{6�脖�q�����d���+˴��+��3�6#]�|P�X(��åWK`���4Fj����7h>�R·�v�Z�U�a�5My�t���R5��1���@���er�!�{O�>��xq/���<���Y�3%����y���B�d�I��?e�b&�1.�`�)m��l����U�H�&���T���d�ܹ��A�G�S@���{�4��A  �S����3��f���X�D�P_��u/4�cn���`��>Dp&&�AL�}��v�pG�v�ʼЬjN��|,+���+0�.����j��o���
�,a��iN4@�I=���Pd��*�P�̠�9'��@��K�FԨ��S�jݢ��3��p�@�Sc>Ճ��u�Gሻ�[��A��&�����p������/��dr���+_�U��"�ݥ�C�t�X\.r1���4�	�=�ȏ��D��N�"����*��-G�d@�m`O�9����Z�:�Y0���}��;����B�%2�G2v�!�x�c;+!�;F��p���+���j�)����#6�n_�=ΐUO�*<��߈yer�^�z�(d6�o5�V��nB[�ޫ�Ѭ�V6�G���~�96�ُ��cإ=��x���Mٙ�G�-=����H�U�q����t�����%�\9c1�f�P��B��#Γ>M|E�?�> �~��Q��S��}_����Q�z�����G5����}��xF�M��־�wW�)pW�M��֙�9a�_m��K�u%T��]
&RK��]�H�t�������G�Y�����r]���4�
����������������&r���R8�$Zٰ�O������)�b���Y]j@3%hn���aV���T�`�6$n�.>�������ڦC���OG�?��0��XЙ.��tV��?�)#���08�ـ��&�9�\2�S�@슢�49_9	���5��ժ��l�Ux͡������/��L���n�57l(%W� �ӎ�% 2��N]փ���{�ɉi�8�6s����z&��g�bx���L�cXT�i �Km������M��q-$�d������ԇ WD�������K�v� o�i���L�8�<=_C���>ξ����"(��:��+O�SS��B�x���kmzK�����zsڸ1:&�pP[� ���{n��%�f����BP�ҁMb��U
!S�L���S�.u���k��.�P��!�	/� `}���-��P�n��֜f}������s��@Q�[�*�y��c��$� ���U�{n���I��u+�6?�,����5 �q#6�SΔ�H�^Pl� ���=���þ�[t��F}�E�y�Q�)$g�ض��1@�|Q�y-� �Ux-YS��?#��D# r��L��Y<	�P�/�q��]��r�}����?�5}Ї�1t��:0>_���b�	��58�����rS��KEv��r�ig�e��ۚy�^I����-!.6��fV�'��*�]�X���k��l� ��a���b+-�\b�ݓj;�TH����OXm;���������4�P���!���a�0�V�<��I4E��-��-g��d$$�!hZM��&vw)��cꨒ�����(N�ֶ�����U=*́`"���P@7�C���|��� �R���ꗫÎ���nsYq��%�T���d����Xcw��{�"=p�A�tF�3���64W|8���_�Q.��n�J�?!���m�S*��)�^R��	L`�%�T��Doi#�o�e�NfNn*�`�Z�|�x��W5�P���L�;���.�8�mK�\�E�h�5b��Y �.��/��B�����O�S���K��ޛ��<��Hޜ�$y�$J���d��S3_z۝H����s�#$����@�BJ�����I�$^@�p"� 3���B�(a�bI�?��������g�����p@$$���&�҃;�������и�wr������!��C�DMZ��~D[�e?���OU���NM������5�ҷ��ӆ�NA[����S��x4ܷ,=�S�T���J'I�	N�ޫ�:��Sc��ec.�;p����}Hq�}|Q��>��òq�'�T�Z���+�;*�Y@�:�J'�h!D���;��P/<Т��}�R�rHf��?���T=*���a{2C>Лq�����*�N2�m޼,+�|/�'/ÂlX�%�u��3�e�%IDAA��U�/���UּKꝊӔx�z��@�F�-z�M�I,cq�ax �&uf�Vr {�BQVI5��E`
z��#�#%� g�'D[��dV�2`�	o-h�� ޑs_ܡ.iF�4Ҏ%ҡ��FϡN�H8=R<��j4)EJ��[���x��oC��B�n^E
�Z�#���p�(��ęh��24�"f����jWH��%���jکw<��75��5�T�`>��@��js��(74����tj5&U�;G$`�q2�4���Z)>��_JB���Q�d��H-��˦.)�o%Ӭ���)�*� ,�9�5�����V�A0��b>�)��ߗ�byI�ĉ��+��#�� #�}r.Cր/��=.��5����G�pҺ nW���T�o
Gt�&r�
����G���*>��k�k�/�1U�t�k����tę���#��>����'�R�2٤�U@�`Mn�?�:��Jo��_�@��_�/�o�'?��!TG�++�B3�({y��f���Ӿ)�ٶ��;b������w��\s�Cd�U��tc1���=u�-F���)� �����!��ǵ�+��-`�t���a�>��3Ȓ-�ֽ�cш�B���B+Q|1T<��v��[���Ž*ZLIK��Z.k:ذ('BN|j@������I�B�[��IK�m�am'6+6�ű�5My~��r8�?�^.̈́ۅs�P3佟kn�'װS��;Ԧ��>Y�R`y����P j��E��0��L��n�H��d��P��^9DI�UR�����N��z�WZ�Mx����_@S7���I��s)G}�����|[w��J�`˂�\���۶UT�����ʘ�jmd?g��qfx��՜�dD��!v����+p�߳Θ�x�I���Y��T��)��I��7(�������	nb��TZ�k]l�!�$6�^m���7��|� `$:`խ/�ϖ;�TUbs}}��>Ş�PP3,j�֋�/Lm6셞��?bI�����F�P�d��W�(����m�X����V>�mаX���޾�/w� O��RπDW�y��q�I.on���T�Gg�j��s���c�1�Y��+-;Nk'�{7E�62�3���$�	�/yͧ�c\00uⷮz3ͺ(��V'7^.�����$}�� ̳l���$:��/��|�]| �=XU�D��r7B:���� ����9���:ۛ�If�����N�=���_	�|�]��� ST�6�.Y���[�G;?$�x#-A�����Y�=(��g�.;��.+ٷ�c�Q7��(d%8�:s�I�=>��YlM�)�t��$��6MہYbV���FqQ�2X����wI�N�OA�=��Qn��mmI"g��b L�w8�b	���ǂ������T��߷���R0h�6���p�YZ{��پ� ������<�=�D��b�"*��"7����@<�/�8��KJh����l2Tw�de�:�k��х�V�:6���G�?&����S?����R@�� �^�GpW�K@��i��]7����p��9&��;~����L�c���@S8�&4ʼVg��}ޤ�,�?6z�
�E ��X�<��\���	o�L!P A�ʅ�7{x�
�/l	�ʌZG���|��L�*�f#�`�>q0��_�NO�|���!�v[�|1���z����@˛������E�r�;��C��"����N�粖h^QX�&���,���~#��3˻� ���!m�Y������E�@3�̟9��9M# ^A�]k��?��2k�<Ff۩H���՞���{��O��#��  m��Ѓ\KeD��Y���$�����/��w��ُŸ&���mdf�E$4S�C(J��/�cc�<0��$\1��J�Q��� u>b�:�z^ꬫy���f�jgHn4��4��V�J�rE��^	Z�/�ˈ7��)���3ݨ�Tp���{�����t��fƈ�ݓ�"]u������I��2�p ��˟��<�����7�c�ڰBM|�p�G�?%�YE��0�7-��T��@�*w՚E��SJ�=���
��\�T$�A7�������1�;��(.AQvr�����ҁ\s���ۼ9ӈ����<����݆Ʈ��/h/t��,����Kμoң�S�a���~����	�7�		�YnE����j�A�y��z�2����՘���&i��ˆ!��f79E9��k6]��
��d<�k�誘���Y�)܊I���3,S?��qoE�^�+�}7Eiyl)�D�D~#��m�Ft��f�. �g����=��)�u�� �r{��I��u8��*�mE"S�Q�
�c0��F0@?s/���Ji�i�W˂JL:�t{�\�i'G���P��G٬c���m9��7�w憑D�ÇWQ.�[:̂X��) ک�5���_ו��$"W�_ �4�ѣ �D{�gÑ�2��}��Uy
m��	�Xe?(κj��j�����F�*�|���^�Px��u�n�!��� :-� �9F�#+O�����xx��λ�Xs�9��,�^�:�B�~e�kW�H��Sa��4��I��=���|3��|�I�S�\�����5��^Rdys��j�'; Ԙ����6���b��@f��J�V?��8E��|��{��:�5�8�N���*����aȸ��{ViH]���Fp��_�c�lyN�������Tӂ�e��$�7I`��!amJ"#��XP+�9{�	���|0��H��ɹ�f�nK`=��0���H��<R��"yU��R��n�3�| ��*=9��WP��?�Ye%?8<WS��m�V�9���V�W.z�T��v��h����M��ɩɜ���	!�}T�>4���ML��"���ް�q;!����f�E�l�^L؎�;����d��St��J�+#'��ࠨ��
*��+�? Z�O�9����GG��q�F��q����F�ǁ���m�A� �ߺ5���_�3V)�@��v��d�Rt:s���]�C+J	�ۗ�,�:�r��?L���vgj*b�������E���pv�/�l�I�-�粆ѓ�����zڨb$c[��}_j�eL{��|�b�(5c�YJ�8����M��s/��Sc"�����㯙ߢAɦm2���P���$DZk�˦;@���|GXH�]I+;��~]K�?���g-�Q,�9����1��d��2�!@?����7�W���B��/L-�}���2(��m�Mw�~����z�ɻ8�����+�� �Y��p�EM'��`��g�X�L��*�7��}x� ��֦$޸��bo���d�.@G���b��D�@T�[��*�9:
Y����i�Gb�"Ua5*>n6N%gl:E��}��)!���-.�*5@Q�ms�\�y3��p61��G���i����� �ur\*�܆?+b�n0'�I��,�]�u�<� �\�F�	°N�aq��w�04�G;�o�kr��$�1?e�p�����EHܞ+�;T xV}r�zB�Hߑ������@�������A	)K���?؎���,����C����G�铽'�<�L��֭��N#�gJ$�/���^�_��Il�x���FF|^�ၳ�Fj�4Rk����+̓��!4Y�|9?�wS3Yn�/f:9D��c�Rh��ұ�:�i��kj�8NyG��qɗ�ګ��V��s�:<.��ˏ3�ɱ�C�����������ؑ��n��#\s�dpt^s>�8�Z?��КE��:�C��#�L��&�Jm��;s�?�QU�H;P��*���?�5���̊��\�ޞ����;$�L׋�"��Y�����ۉ�/0�,�����
E�9o���܎:��TN,&�L�.|�89���ɗ�D��q:�ߒ,�Po�Z�pπG��kpl/��ʷ.�@�^koߏ������7D *�Y/�';�a��'�leI>jYV�E�M4<e��f�~L�x׉���Yg,�l��*ǆ��3X?�w�p�7!vjyr,tǼ���1x�Ҳ@�;kN�����;j��b�W�['?�\;!U<�n���#���[���j�~(��g$*��w�Q.�pG�Uw�5k��y<s�9�"���5��j��~lv��K�b ��%չ�JE��z���#N[��0\c�t��qx��_�c>4ݸ0
@���g�+[,6{�H�J��}��YQ�0������%�滪k��p��P�ʟ-���س �H�DWT�<\������Ҍ!���U������U����+_{4��(^hB�I �kO@n�)�'�Z>y-�u��҈D��O#�\���F:�jmOԾ�8�q��Dy[\\&0j�6lH��Ŋ.>u���b|IT��td��Q4�a(f�%yo��Y����xT�a�o-+�6Gǜ����*zٗ�ڂ�@�ԧ%&�̅�V���fG�1[j CM���o���'$�Z>�(���JA�/�$�)gHr��Y��N&�Y���O�/яw�����H�2[Q��
����S�?�G�o"Q^n�Y�ԎD)Ni�s��i�{��&���L��S	��ER�L�A��7�v���
������w�213�Es�Ӈ��K�Z��[\�/�?h�{��|ٿ��+��YzϮS�n�p�wE�i'��^�m/w
q�b
\OG��OY��"b9O6�NW������*yUf|ϝ��됦�	���k��"ܱ��X��
���f�5��F����}Y���������DD����G���b6̲�Bm!ۀ���i����;Im �O�rD�s,�e���@��N�.�p���v�b����y�y�h�����0��xo�Z�̱�uN�c}Y椇�6+ j��Fy�ʙ"YF)�����ņ��m�1>�з+��;���>���6P��	%�-�V��er��iȶz䘱�7q�F�'"�_�Jbs(T.��
��ZU��{%��XO���t�4b�8�&�8GIT��"ֺ/ۏ��^�X��)|�|5ux�L�R�DN+3�,sYP��,#��c��zKZ��~��J�p-Jc/[c�����%r��u�sQG��gѸ���\^;q�ն3���9�T���<�~A���D����NI���N�zA���7?B"��;��X�Elt~A�`�u�$��K��۟��Gy�H�e5_�D>�~3���;�c��!���l�ғ	Mjd����E�ΑmFL] �m�J,��Ƴm�Q]����k�����=�j��YOA-�l���.��q����n��ϹM��xly�3���ָN���b=�]�F�xX���x%E�g��~�M
��9��g>ђ~�'pp�[�L��Z��/̍+����^3�()�U�
y�}�;ʏ�i��R{?�>c@�CF��>�U�VOX9̤����H�� ��v�\=l����i�q�a��Kq�V���1��_kzo	}�d��G��͞���!Rz����y��ck��ll���hS&ǫ�z'?8f7�]͹��Ώ�.��3���TZ�'���b�u����ܞ�Dn��M�Z��2J}/�kMoD�f*��Y���Ƚx�#�d����i R��vl�2�<�"���^�E�7k__�Y��c�5�5�q����d���yS�æȳMx�i���-Իi]0�c�E�/OH��|"��:�Q�&F*��&Up`�fsrr��cѨo](){o����PHC�m�m�X��P�;V������#~!��ݧ�f�T�����`��D �+���f�~e$�����X�(;�2wV޳3E˨�_�4"߿Zsg��. 
+T��)WPF[.RW8QT������@�2��~#�_5Y���z"�3�v���_[\��wO�̂8t��j�榀�%��|���A��`N�K�"����ͣ��%8>\� KSc1��!z--C�ƴ3`��I��*�D�G^i��F��Z`�R3�{�l�K_f��hT��U8
����#�Q5?��_K͋䅈�q%x#&�|��]$t�y�'s�T���
I���:J˿sU"��g95][mI-���>!ʃȑ��xm;q��7R��{�H��1��7���`c
{�y	��sI8����5V)6��Z9y%����*aJv!:T��y��}#�bi��ݗu@���66V��"��r���o��l����?/����������譂9����ӂ�~�Sss��MO�l"[q����zET/�"b��q��6"�{:,�Td���.��H��F�`�~9x����2˱���F�E�m�����?����f,#2��ʱ�p�e����N��Qy����m�93�#gX6O�s۵+�����!f�Ø�pww�����i*Q.��$��w�޵<�7:�$�`�s���[�	�Ip�df��_���4~����ȡ&���;ȤȡeģR�|�]�Ava��r���6^L�0�g@/J͚-�L�-t;_W�xC�l�q�'����#*�u2�u� ��:���]�H�������� .�V��!���5i�`0Iw$�x��~��� �$�fI?�N���e��f6��ׇ��9e�m�A���*Z(��>"}4����K���i9}��n��RUSw#�kut���O�� ـ�/OX�A9L]D9Ր�Kُ^#���AeHsn&)��Ő-_wi��HJ?X�a�^]�u��;+L��m����D�HL�`�A@����n� �ܩ��J(�KhSh�F�E�OT���W�!��>/��rMc�s���HP�������z'4��D&��IFwж������7������>��g/�5&fy�p_��ڊ��_=,}y�,K�O~�kB������=;҈�wy�Y��*l��knd�4(�-�4����%Dh���:�k?Q��FPoq*	'K{����UZyWrz�N�3�����P�ܥ�
j-�ӟ�U�+�M������L��<X����b� ������W����te�;�����O���kJ ��G�^��~xi&�h�W��]�h$uy�
��{1㲸h}���\f�E)_�4�(Q��1o5��6*N���hM�OW��
����ܫb�j'����;����M�M���>��J$��[�J�-��o@e�L@�;�ژ�1����:#�#tQJW.�4�;J���V�)���Ί2�[fk@|��uBwu�ѼTI A�B��5f���w�5���l�	<3nQ)�s����Й�4J�c�}gi�έ���Rm�]���֛j���x�����h�-׫~X`�{F����i�	�@[ߕs��^ڀ&�����)�Z2WԻ�.F1���׭/H�����v-���*�Y)����߭���|���ɔ�!�<8v([8�'��o����N�7�Ƹ�O�q���V�CC�������n�PJo��U_*P���4�2Qs�y�c=Z�����˷)��"�t�R_��@�\��0�����bDBlR�����%'��0�^^.ǫ�y(�R4y+��S�w�����#̓>��;_�kr��x����b��B��
~�	'4�������b&�/����c��t>�s�, ^�ȅ���.}��d)3��lB%�D��_r�G5�UQj������W���OL;2����s�A�b�s�
���\�Çee��C��s��Zn`�E4��*x�C�}�{͔ǝ��2Ej:]ag�(����e��/����kF2�R ��S�	�:'��m��9��"�v/�~�9t���ǊU�9������1��|o�o}����f�=���އ�~e�go���Ma��V���`�4�O|H�:b�;������C���~�}�}�*��YP�m�᥋�zc�K��V�
&`�4�J�mk�|�3���D1э�	kM/���_�Q:�!d���h��Q^g�Nԧf5m�o����y���y����<7�'}�(.U��}ێ�x���Q<f��3�a�h�<kw���u��ˌ����LL0��C��u^\��n�����_`�5�H��HFPk�Le8[����z�xa	�~�4$)�h�`"��&G٧D�66�6�#�@�<���Y$�jc��C-�rE����.�v9��x[�h;�� q�������=�D�"��:����K��);-���p�P�L,�pID��]P���C�Q��Y�J���yC��H�iRTؠf�F��@�NyUF�o���ܞtc�[�;��.Ն�i�y*�}�/�ڟ��bO��ȌW�l�՞	�ſ)0f��3���F�:��VM�t�4�f����4a�o6����t\~�ϕ��h��K�l�z�� ���37N�M�_��WWK�w~�����y�!8���ķy�N�W*�8ep C�R������yt��OX_�B��ϳl�c��%^4�-�$7h�γ�i��u}y|���I*�S�bz�(���g ��A'��$���h��-�A�@&Y3�=����6�j����bE�6Y��4��0�R��@Q}�g3�L���:	�N�^���&�� �����uH�{�������E@xj���o))�F���v�f��꼗��ug��&� �<<=X�Hf��.�Ȓ���&U��u�l��=����s�QL�s�ܲ�[���l����fv�����i�4B����U��1��7�];xmӪ�8e���g	�<�<*7�@nI�G�;vE�5���Osêr~�X~0�s��Ś[ v�(i3uf�+8֝x�~<�	��H�>TL{�<R��BT���4��k?E��0/��5%a�/*-S�Roa�%�n� :�0���s}����h����$(�.�s��!>I�o�uRϧ+�[�r�\�"�)�˳P�G[;��ɳGU��=� �ԡ�2�*^]��u�٫|5hŧS<�r��&��1O=_bV���X�i&�)`"����S�Y	x���d;��	��3b\��/����N�-�f��@M2���R} p��M� �c�L�d�'}�i=�s�˝K<؟M���St8�{�b�I�d��ˁ��
�v1zza�@��Z����sZ�G4jǻ��-ʦ��ep���{����Y�2�S4"m,��܇�Y�3��z[�b���[��=9q��%b?a��uWb!	��2w= Ao������v�<1�k��r| 8l^P��6�_5g��s���]Ҕy��s�'LNn#�&$7)`�$˚�o�������B�2�5�/����,R�=7]�K�b���16��;:�]P�0��฀a�.��Z��{CW�{��#��G��Rr�8��b�1�����e���#��)?��T�n0�V�e�F9E[kӺ����T�0����G� ̃�e-%����]%����P�_RD1GL'N�����f�h�2��'���i����`T����k,p<K���D��#	��@V�m�xo�0��6�D��B,��&���h��Z.�D`��%��*����{�#�V/Nx>MۙJ.���v *xN�`���{��"�`Q=�f�G8S�Q��v	6�_�s2��1�8�Yq������֏�p�R;L��py����ս���(��*����.Y���Q%u;K �:�pR�{ G�i��H�}�߭Xo�B�//�V�CÆpX�����^�h�f���)ƒ薷h'�F�ϡ�0����7F�).l��� V~���t�g![��d���x[V|��F׸��Mh��E��
�XWW�&A��`k��PXIW�3��ϫN�:	�Y�{��l)��-�%O�n���k4I�:꣇BNyL��4&;��N�B��Bor%���W��v�]$k��qĒ���\�}��(l(��5y�Xͦ��2$�;bi�XE�we�Ý/���1�S{]�ZX���5F@�řC���t?ʸY�t*ww4:>� �*_�B���%�脏>\Q�<�gG��k�L��p�N�&s�����,(���srF��z�zN�I!2��~�$�1��<���}K�U�W�AS���Oc�Nk`��I]TWw=�����3�Kr�L�!OE4�G�XD�n�&H������`
��gBo�0��Y�U5�Ɩ��jB?�:J�ſ@_Y@�n_e���ټ߰.f1�e��;֐Ou�,�
h#ʰK�R�B���T7�Di:�/���@v�ҩ�̭�h�$0QJ
��E�x�J��8�Ț	�0i\�F p����4�Ui�	��e����:�b�?��2t��Uo\�r�u���ʜ4*��T� ��4��I#"��a%�rR��Ӳ�]�6�8�ʐ�`r�2E5��;F�UFޔ��Ao�������d����6ŗ_����V��

_�������Å�ř[���
�Yn��z=��zR!���B�ku��}��3�;0W�@i�}#d-S�wGl	{yrBjO����Zǹ˭-� ���h�S�YXr�8ùyT�����DӠ �r�n���(�/�@������<#.��me�׿�X�q�>f�>.��_��n6k�J�V����5$������s�������<�WvT��:��P�I�c��#NCyפH�G�wz�i�*֌;��T(�0e�%�ۅQ�a)����
0��צ(����+� �|j������ R�c�V@8�������25ner���`w��ޗSG8���qgQ��VR��4�i�-k�T�aݺ_u9Q��9�N����.8�	O���T����fA��]��i-�ۗ��]hd�
����::d;%�0�d��o}�8�C�k�N+���̿�����}�!D���2;\��:��,l��ǈ��x6��m�et�d�l�!�y�և��Y�����x����2rb�)9�F��P�6���&�cP�{Ϳ���X��<�W3�s�ò~Aq;�\g�Û4Vy�	k�n��S<��Hn^�ܰ�7`0 x�]�EԾ��W��#�L�$�dD#+*<�7\��s���(��R��/����q����0<�L���Ċ-$Y�<�h�7&��˾<��IO�劤���Q�_|o @\�11~�(��}$+����⪐��O���cƕ�5�	wq�����I��jUj�����&�g�mw�E�*��ȩ^L�W�^qG��=ݖ5^{a���U��5ˏI�fn*���1��`����~C�Qr|���T$�2��fW�wUS�e r�S˘-.9�E'\����׌� �o�������s���8��Rb��!�X��Q(��A��}�w���dG��z���鐘�[�^D�P'�ƽ�>-G��h��R�c���"�)H����4��]�X��4�c�����>N�J�̕��2�<$EO�&$pM��nP�b�/W��s����1�I�+���;�=�g�;�{��
8��e�D?<ʕ��!���8��	W]d�5�����)�:l̚�h\F�<��&k�+�E����ˣѲ�6&T@��bG& H"y����-��\"MD�W�G'K8��~���v��K0;M�����7�##���C���树��5�]������_h֝��x}\�-�#�/���8��x>X�LA��/�p��^v���������g����8U:O�V�w�.�z��9�I����Xvo�WQSN�y�N�b7���g|b?T c�N��4��è{#�����ù�-�xLi2.i��^{�`�Cv�FG�qK�h��{Z�$>�9��ܻ ��ur�h��Z��Oj��W�[��|lv�og������+���!b��Q�)�]͸R��[�޴��aC�hߵVR��,*��U����W�d+?tAҟ(�� �#71�
��E��-�6�bxv��e�@��fه ������<���qǡ�js�`��	���>�l�����T���.�Mԫ�t���m����!���)TP^jVQ�����~�E��o�G��䣳��a0'���Q���#��m&���fi��({ʞ�B
��³�`�<���W$m����f�z�<n&��:֢g�؞h��������Fj_I���5'��	cT~��^�j�<8�p�������"��d5͊��K��4�ii��I'�Z���o�a@���y%�T��E��*���&�v����d�f���& °�x��6�L�aN
��!#���2��^N�~�W��Z6@�P4����]*��40Pj�aܐ;�I	����"TX�J��~�N[ޗ���C�ϩl�d��T�_�WEX'tV��- dO���AgX�����9=^'���>m�R�_��
H7�����r{$�4�~b~Q*԰8TQ<�'��[����B����[f9bϝ�q>�ȀQ�USƗLiZ|Ŏ��Tsz���3�!j�%SQ���#@��Di0j}���m%K`Q5ՔPC)��Y'�d�BjG���/��"��ؾ��������n�{I�q���Z�E!�re���Xa V?��}>��b:�oF���o�o�
��F���+#��������p$�8l4M��X®�@��G��G�`�@��m1H�������S���z�_5񚄩kraI����&��]fTZ�Kvj]�4�ʛ�Z ��=ց�ժ�C|�'  y�|ڃ$�3�
O+�2WC ʴ�>Q�i��ȳ�*e���,8��(u�d]礳�K� _͊j��<�X��x�cm��!x�bp!�o����3��'���wy�+h�rL�"�#���WD��;�6A*�U!f�/f��D�pZ _Y8����F������s���S�5�x̭�ܦ��L_f����3�Rm��-%1���� g�g���L3�`/g���MW԰`ځ��9���e%|��nd"��Ln{8;��&������&c�֟�)��p#,�zBӕf�H���i�����=��:���[v���#�k�7�`��{q�������9��d>i�;3�P~GC��6�����m���Z�Ӎ7\5/kc?ݦ�dD[C��pUQ�q�[��p�͎�?�	�*�wo?|^R��8B�(�����ZD�MJ����90���/�$��{�c�/���j�j������}��˻QXiG�6�z�pj �b-�����92tHg�Tj��b`��8�~���a�[�RJ��g^<����]������g���FnU^��$��t:��T�yFpa'�q
���0����80�dE{KT�� �E�oX�;H»}�: ��_�,<�7ֽ�^(1��n��6+���6�����.NP���6�x��#�K��������=�v��F?J�����D���o���(�E"��m�K����Q�v��D�䯵!�t·(>�[�#�.R���F��O�8�R'C��®�Ή�9�쐐&��9����/��b�2��˵A��ĝ[���X؂)���,��d�̻`���ճ���4^q�?K[��"�����.���呚�.��2s��a-'ܪ��=�����p+H7t���4~���Cp
���7�|h�ط�EQ�󬽩.R�)��M���:��󹾰��l;��נ�g�3�gZU&� X�o����3����f��͈s�@k�hZ�8�G~^��uZ�|�<����8h�3��9]$�w6���0�8�+&��h$@t0�ֿ�M$�߱�n����#Jl�b����E@�<�u�ٔ�Ԝ:��a̼f�E==*�#5������K���� }p��+Oa�Z�\z!�yI:�ov*�:��M�y^�q��f���T)v�o�RU����[Eq����?���{��ݝd�`�ݛC�BCAЕ��?�"���is8�a�.��7. ��*���v��;�pWV���i�=Gw��l�U�vM`l[�_�9�Γ�f|������CP���w�euc����C�&t�d�x����	\�r�m=T<�{�5��neIBS�J��u\(�u�4P� `F��,��E�M�'oX�siZ���� i{/qZ�w猨j1=�
�	���,B{=�m
s_�83�Q�0�gX�z�^�eKD�ϐ��~��e�s ��~�ޠ Lx�q��u6����S~6��H���dJU��V&b`�Plyd:13�6v�n��_'�0�b(>=���.���u��׎���� 0@8O�y*��3�+uB��ј�}tÌ�@����ď֊��%T��A��z�(�P#m���E���l��:��a����i6��Pj`��b9�����L���g������Ƕ��f�aת%'|�ڵXt,n����+ǟX�B�7a]n�/�y�LF���� fx�������A>�Ku��[a0O��?~�<y��.�������Nbi4Y�oաNV`/ޏ��?lJ?�bJ��7T��'U?����	�	�k�?_�4�6�WF h
�I˦�PN KJ b��ݘ�s���(#�Bٖ��Rr���_�b�@�n�;p�8�˓��׳� ����8�W'�%�4ִ�_*|��l��A��گ�︋��U;�I�G�ز���p��k�mǮy�%	��^�b��Fc�Z�ϖPv�6FS�*�t7A`� ��c�ݨ<�d7�wN�L}�ɭC�����Rs��Z�; �7n�����"�aZ�C
ݔO=8yg4ǿ�1uz�1��x���=8?��=u� *�ʉ��ɷ���z��l*++�f�n��g�h4x��E�&�0�8s#g�V��-�N��k�l'����.H���ܒE��PxZ�"��$�*�X��&��]�gr��kY�3��䢔�
D�u� g]���x�k�U��_�b��pA����ϡ�+��r��gڪ(�7��=x_��w;�f
>tt�w���(��F�gI�j���/�U���f�ښ�Yϙ�����g��q�ϛ�T8_qW!ͨq���)�\
��z���:~|~d��a0����+LgگʱQ��COW�3���8z�_�Ty��w7�]�P^��ؤ'���0��-Ҙ��w`�z2�O��z����YnO���c�p��Y��on!;;��JTZD�y �B��KA���7�B�=p��~�K����~���v���=� x���B��߃����C'�c%|_�R@�fp�X�dʅl���� G��u�u��^}ē�l��vU8.�S�H��-lȐ�%L} X|f��>� Z��':�z�e�!��tܱ�Nݩ�� �t&��~�ǉ{Ƀhv�Nd?!��m�HX���݈ҥq�(!�>�ý�g�����)=�Zi�1F|��FF����q�i��W�U6��Qi��o�h�L�8AH�;��co���^B0p��d�������.p�(�"�W�Ǘ):]va�[�5_׽j߯Z�+8l��^!�!��RQ�.2Vt�c����ě�����#٧,
{-�"n!�������O���&�s;����$���T����R/�j&ÈH�^��\X�כ=YDR}f�������&�ErUd���������A��Y>?*c̎����6�M�%�L��8�,�WǢI�w5�Q"1)R&��:ſ��c�l�/��;�<#V;c���
��&���Z���e��G
�ne� ˟V���PA�q���', ����ʷI�u�5�%#�^���l�z�Es3�Bq� |�'��1�;�.G��ӈ+�$��v��8w��tc/]��+��О7i���30��Û9�� !��!���O��ݥb���r}ȑ��F[�R�S�c��^�Z�S.��r��1���kr%-�9��b��G�l�9�qu��ʥ�1d{�qz��_]�Hg��+�G�j��mDBY �ȭ���p�/~�����2W�E��0%Q�W:�^��I�b����v�b9�<��/&��s������"�n��[�)C^w�4��ڍշR;��}�oƐ��χ�qw�9�Hז؂y�\�������b�F��ɓ=��	.��[���{9�*���	ԟ�/�W_����+�]8�]E�pIh��rn�m�]t�z���f�C$6Dc`|B�5+#3WD섭s�A�/
Y�B"V���P�%��}/��G���b�-b�_�s|Y�2�6�Wx�(G��zAq!a�$To�j��X����
^Ń����By]WH����4�lI��>XR"���i)U�Da����E<��y�5��l,-�uFt�
�g����{e؄qO���W!��%dM^L��rTj�=��i��!P��JS�iY�uա�iڧH�LN�M2U�c�K��)�a�el9�-/k�}����\�D��N��Uu�q>���]!��Ӥō@N3�;'�
E��EZ��XZ�ت0��dy�d!]��� �[������acx��r�W�}�K��� �W�/���t�sV����x���ɔ�{".�z�/=6\B�oub�����ƽ݄ws�Sp�Ҕ��,>�؛;��x�*���*;�u
���y.���
Go_���؊��d� 	��qS��z'�I ��L:y����d���⭮~�-��dzt�&�=^����y�����ot��w��[m�OG��01z�[&ߩG�C��A#�Dz�ErX%�Xi�]����W�Fp��y�?d��5'9��-Z_�ժ-2/����j���0Zj�#NO�)N�* ?5��Y�9e��Y�ώ�#-�G�m�7�<c����$
��Zg���4Y�ʱ���S�B�;T��gz�(�|����^&ӧ�Z�Y9
m�5SY�)��ȣ���?�#2��i�:��VTP�s,���W�ۗb�!��l`\����E�ͅ"��olP[����d��Ψ�����ٴ�D��8�v�ͯ�����Eh͘�����eۻ��[P�������!�ڡD~k��]��4��Q����@(Ad7M����z5��l��҆&V	��h��䕵So��+4��&��Q�Ń�[��m�7R�e�
'K�M�wJ��b��?��
�=ʎ�!q�Y���<�S��KXޒ'ݍ�B�P���z7�Tw���|�=�M[@aP�����l�������&�@~0�[Q�j�AAS!�܆Ga��ԃr�#6T�6�H�ǝ��fd*!����&)�'��q��M���偲����A����4�P{f�N��qI�y�ŉ.Nam[3����y���@\99��/�Q�*�j#*��֙FeN7�&nK�v'�՗������Z0.���#����W��Ќ{���-�a�"�z�3�� k���y�C�IV>��y����Y��Xa��ٝh������1���,�O�O�%��b����U&���T;�ȫu��KY66Z3\��8�I�R���4m=���%q�eؗ"5ZܮdR�gk��g�v�T�5r�"�_P��N�J�?�%�VWtR��`�q�'n1�a�i��m ��%c�{���#���ޛ�����[sn���_w%�wޘv�{�Y˔ԌKL�u6#�c�)0G2B1 �p.��՜Y>������MT��C�yd����[Z��Դ~}o���8pJ	`�4K�@�h�v�����X�%�b�j*�ՒF��$�Z2�݂V'�ӗC�<1��3}��/�C�eL����8��U̞�3���0��{n��aq�����݋���s!@��Cӽ9ad�d��tug��8�G$�(�l��?Ey ��8�
��@Q�v��ta�	�t��r���^�l��\.'�忠��\�~h퇛}�B�6��y�M�[�N�� ~��˖i�RL-ǳ�q�V%!�L@�ɚ���?N���a�Z��7ߛV���/���3�a=��� D(����tT���x��w�'Y���0u�X��L�<��Jq��G�m��k��q�̩4���҂�㥐�dǾ��NU��iQ[d!:���Q�Oc���)&�<z׾�p��ɸ��L�F,iC_�B�]�>Uȣ~*z4�f����7-[�}�,U��<T�S�U�����;s>b��ӷi�`C���̞����c=0|T�`���@I("s���5���bۭ�W�0���œr{� ����8 �_*,��n;�d��t��%7R�(���0Zpx������.L�/캄�5�(�;9��7��W�P�f��8N��k�L�+AN��Hhk1��g���I;+��F��F��[a����,藰��m���Y
�x����І����%PAs�
��6�8����W	�S��ȇJl�KZX�,;����;g��t,)cv�^��11^����׋LE�w{��)�{x��m���HC	>�P笰�����g�:Cpp~�@��_��)��vr��R�n!�X-;~Vl�����9�C�c�������ci�$���J�	"c��d��@>
_L{ �/�ؼ��d۠ob~=Ma�֦�L��r�Kg}mY���V�թPu.�-��_j�Sߴ��X�iwG51	�l~D'τ�^껅��$D��eJ-ЊP���f�SYT~΋Ap�n��WtұΥ��m$������WX�#��/x/�n����a��,�]�E
HT,T���%n�>�ӊ>ya��=?'������;�o����(2��(������+?L��̩�֢I�s�F�õ7.=- @�9���3�P�#���,[{o��ڧb��7)r�����婈/R'�����IXݳ Ӌ ]��{��W�Q�.�����m}�q��*��s�;��S�))����'�������S	�i)H�˛,�����h��C���r�T� ����Z�^�kW���8�Pa�HO����w�Ѐ" �O ��8�:�0�{�_��3��7a����|�ȝIR��ZI33���-�!�ޚAO������/+k�I�AtP�
�b}��]���C�J�$Bv���OJ%�ˍ�@�,�,�Hv���*�$���<�{��]~��'"�6��1gg>R���?،�3$����_EoH���f�.�W���hभ��	<��R=7Q3%յ�Ҵ��;A<O�!V��B!0E!��ZwM�ف�s1G(/��v}G���(<�1>lMMi�m���a�+�?�[�����/'0��o+^[O�A���A��H�w�.ϯ��p��Ȕ���9d��8CR.A4׊��ݡ�	���i�"���TC�n��R�Z:s���9@ur��W�4����)���`�Kv��F"d��zJ��k�T��`+��f�O��׊R� �t��_�o���M��(K�,vC����ډ��H����ĨB�|NbX����{����4D	���k�.��8���PC��)K"����-�k��:~���	@�3p��|�g����K��[7���j^Sh���/>�%�)r�i�TT�E���M[uԲ���g /jk��y�i� �ݲ����8���p�vY������N�4�S�}};U�P:��̚��ڗ�z i%��#7+0��^ �\��4������!J�+�Ï"������+�i�aϷ406�Re�¸�G�MU^X�{A�����Is���,������Jx�>���<��/��\��:��`�Ȼy��nP��m'3��qi�"���i+n0�6���-et.X�����KDjO��G� �T0��"2U�J3�ծ���B]k"[�4szN<�~��$����X馑F�7#7z��w"xsX4$	'����X������T1&��*��볧�(p���u&{�O��po�6j�ţe�>M�7�.5%�^�t��Jze�I�	-QO̙�C���)=�X���	��LQ�cVA�< sh�FػP}���:�鴖��%��g��Q} �$�V�����vSk	��p7��@;���g��wo)둎�a��U;9+���k��ኵHT��
Ti����Ċ��`�]=ڶ+C��|�WP��V��͗�hxP�BU��1F�c�]b�,�:0f���8�+w+�#��(d�B�S�k�!�!d��{���p�����S�N�7P�{�k��U{��H�}b���1,�Y ܂�	����g�`��N��`Ӳi�ʮ�� �>i�au�~�˘��z)���ҭ��I.bG�6}� �L�����d�YJ�S�����&��5'�p��
?u��P��U�q�?�}-��R�sU�D	��Q�!l�:��%��A�ڟr3MN�$��ɄJ�TX�5ћox������|v��,�+c���&�tj�j��E��kj��7�R�	y�Er���"*�Jx{�;a:b�^f�6�^y��
��Ә��yRa�Ly`	`��|;�\mHmE�*�k�|ʯ�j���~X6��)����H`'��;����b�d��
�=sn��؀d�s��1N�A���Տ����!��A�!�����^���w�ڴ�h����*.}���Z1���)"��*��j�t�P��)����5�3�q�IE�_���cw�g���)?3��Ng&Mw�M�����J]��3���tQ�I'Ӄ���G^��Xwh����r-:a-�����+���?�3�s]�oq�{<�+9���y���Y�I�[Xө��g��seN�v�)���l����m���T|���Kl�C끯�oƥ#j���_ �wyA�`�Ʃ����}�����w}{���,)�9:�Gqk���1[�ۡ���R����i�"6��2�/�q�P��κl3��gz�8P��ZZ��D��HZ>gDGO���3g��vu�5N�g'SCSX�8e���F�ZɽvMT,%��ټ�x�	<�n��fϗ� #I�MC`əb���L}v!�ŜP� /�����BXvYG`=�VnFS��v��:���Y1�[��o��t���
#ӳ#�SJ}�-N�ܐVX�&�Ҙڛ�����*�@b�|�	�D�@~hj5v/=��nH�Y��2�gn9��'{�x��=�[�4i�M�e	P���}�]IIL�4�PK�>5B
�=y՚�O ˽ݝ��dr��N�@��Y�NU`�Jw�G�X�#^R�
_YcQ�V����W���$��!t�����x�k�P����#��B_���]+�=�ܯ���;p~TO��s����Jn�i��Ҁ���L�-����w��y:�� �V�'����~P� �q�N��f���@����޼l����3f��Z����:Wj��~��6�\)��6�C�<Ą#9}�ي7/�LV(c-���\�z3Z������G�{-�]�K�i�=�J�PG��jN�W.�-����d�}���4���K_S���y��6��2����c�^�3"��i��C��<O���4+E�D
������wZ���Q�I��Y�ƥJ�G���	�n� ��3���s(;��(!�U�9�̥|��)��H�h�	��) Fm��g����F��]*-��2�^x�Ug;h�؅���)p]c\�����KF?��P��ț��3
R�%�����C'd�Z5k��y$��`g�dm�L�!��ފ �>���5��q I���!5���h��*;�x70#q�q�N�g3�N�5ifچ�Q���O�r2�S9�,:e��Y�:�r�q:
����dBʮa�f�V�ѝ�J��[��C�Ɖ��D�
j�4��ञ���N�4��4{�\�v	�o\c��sqB ����|#�7j{��a�ń�cM�p�.�!��`m�ʳ�S��H1�����A�����)SKUlѾfQ�t���b��;Nl�`��(�
ܒ*2�Bu���{�Z?0å����݀MI�s��1�i2��۹֠4��u�����WR���3�vGe����Lz1L��,��;�H�,;��dDh��]K�-b(7&j���V�C*{%�͑?��S�u�ہ�M�u��C�'�@s��(�k��y@ES#�!9x{���Vz���0
�%���hfHHx݂O��]h�G������T�����H��&u%�8@L�` ���~`A4)��؅@��~]��[�+贇�GgxM(�`��5��t��B*'��e�SǺ������~+��S�@��7��iX���b�'��^�2�ǎ��+]�:���/G��e^h�R��o[��.��6I:�ߘ�)���e�YW��+D��G��	��|p��053�vX�������fݯ�-	&iCʳ�O"Q(�x,^Z���K����� ��f2�ZC�{�K�'W�L{*�/���O��+?_N9f�/�W�|�~�x��(����~?]EL"�q2,��T\V!n7� 6�,�l%����B�ܩug��ǔ���,V�=�yt���β���+ࣉM[l0���?W�xF��$sh�ž�/��hN5���0��A=�%j�&��iޛ_6��bս�$oh�� ,�u�8��7��փ�M��D�͏�$����7��������*L���H��}�1$��8t�U�0Q�>�C��Ӱ����:��=��  3���j�·/yŭ875ܿ�d�$�_�Ȱ|�qZڕ�Ê���<b�R����z��h�"N���%/)��=X��	�F��$�ֻ�ϫ&��=� -#Б8�e�hL���z	3J�脿ޫ/�ChƖ ڄ���8T�l}K�S0 �ם:���A38�9N�C��c��?h4D{��ݠuO�V�m��FA��U�&.�����������(�Kac"��fN�T�`����5H��¯���Ae�C�Рy)I&��x>J��A �iF��E�G�kh��_ ���u�S����3����;�	%c ��"0�.q�븙Fo����ƣ`%���eZJ��a^��
FAP�L���M�[�s�㙭��V�P��͵`]} �J�;k]p���$�R��bJ�þ ��M��j=ɗ�V�b��a���q�Ź��Ϧ�7x�)��I�V�Q�C1�,��Z���'������H����y�����9�qf�X�Kl"��<���4)�h]+9;�&ɲ�l=���v.n�Hd�� L��v��>�D4��ai:)�����]���{'�"}I��2(�E��ͽ�f�=d�$�?8љ���_�wx��Y��[�F@�����������:E!f�����9uA� �Zvd��a��*�?��$M�s���z��8 n���L�aQ ����R {7�)T���t�a��*��@�b�4�����j��=:j������ds- ��e�1}�!�Nf����Å�qj6�� 2BL�F��#�h&Q�B��k�^k��ks�r���w�b�d�E�6&��` X����1"�6�jR��1,Ϊ7�~zP����.9���t0sf��P�� o�YU��� �[�x~"	@$k��z��5��$|��?���5q��ʤ�ސ'Ņ��k�t���a�������)~��c�}4V�`���#����@�W�VA�9�=wbn�D��X\��y��_,�J���*��{D�0K�)���0Tʼ�܃��ʢ' B�R�mV8N�ݖ3�.>��$+C�+��x�%"�sj���C!1��N���i�?�Pޤ"�V:QD>zy��d?"�E�l��S�~X�Y�����1���P�'�,�é���!��Mpa*�#S�N�I]� ��#!�n���ݍ��\��KX$g�nB�dϟϓW���<d��<⚗��ya�)�=�dH�KMP�����Jo�'f�*�.�'�0�c�H�N�h+u��=��TXJ��%qZB�����_�9����F��6�_��y�v�H%7�\ �(J��B�>�7�t�+�"��d�Z��2���Э�q��h��<�q�4X_��?qSV�a��B:Ҳ�¥L>��|�b���ɭ�#���ǻBeL��g<Gm�xa	�>�Izacm�蚩J�MX���Sk�(a�Ǥ��`_�Y6���-��b�1��-|�-9�i����*C�s��G$��0���'�ٙ��$�����[��3^�w��hE�I0����j�:�� *����l�DJ�,Ɠei"�H��X�Z���m]�g;Q�W9C��Կ���#��˭Ń6{K�W�B�Zٍ��%���D���/�8�f�w��b�/ԃ+t�J�i2�=IR�������ʎ�m�"� ��
�3���r._]}���w%�o}��.p�F�0�"�8��}4䇤@�j��,��.G2��r�/�:���iiTB����2���1Tnңf��+�q4ʁ��Pq�.*ec�s�@,���t��|=�3?5ՌQ@�f�,J�j2��Q�i��r�|�"��9f��b�y9��z���6�v<)'�	g�H(�y 9.6��F���M����MMEN�'_h����I���F�q�3i́�_�)e�g�+xC��{���8U� �r�Ui�y�Կa�@����j���(,̜&_>�ͫO�վ��b�Yd��Tr�Nб �!���ܐ+�N��fuCY�,actGq�e�hJ]��F,�޿vZY�+��i=��o���g�&s��Oz��c1G��EDI�j�xV�u���qrP��5������W�Yw�fh�C>)UJّ[<��Q���{�����Do,�{����f;s�}�egL����0���/�x�  ���2���$��Y�ݎ��%��'R�ۉ֋��-e�=�,����[rѠ{O�1�\���6�7�m��'Q�5��G���g�I�����WC3W�҉�%���o���6�uo�U��N�*�Lg]bXF�n؟�;�3|�0	8��'�&��^C>R�jj�r��zF��"���TD(=u�r�v�5�{��9�3�8���Wբ&�v=)�)��/��Mn&wb������Qz���,N�^+.w��zF��u:����|F�e�=���d=��+�ml�ɓ_��~���(�}�k��ϱے�
����T��s�@�ٿ���Q%MkQ�b�4���D6��?H!�N�W,��^�)�mW��&�G%9��hx�(L�������\�*�b<��p��q�<�'*�+8ރu8��{�K�ڿ0��Z2���V���k�UƎm�$?�	flі{�����v���t�r��ƽ��(��\�yY�2����p£f�C���^|���
1)�b�(�w��~�[a��X�ƟN=��f���{*_T��@���Ͱ%"4X*���HZ=�$4*c�C�l��!FJԽ%�(�:}.<���R�yĜF��L+��H�F�k2�m<����>H>�9@�V��(,]L8E@ᆿ�Y�l�Kq�<�1�>�v@ ���3˹1�zE�D�4�Φ)Ir�,���A�T���V��MGV�u�z�Q'-�m8=���YER�L�{�E�Ӹ�ّ^�6�,:��aN�ٿ���r��J�����]�$�<���5��7.5-Bh\����;a��C��|:$�٣
ï�N��*u�ө2i颭^���I.9f2]DV�@�����3�18�ܪA��]�KP3�=��a�`Y1���dF�mF_)���*�u1��й��K��5X�ULsDv0�(��QT���ᘵI	�>b".ޥ|"���y��#����;%��/m��`c�j#D�O�e@h�q�DF����ʥ�:�W��1QbYQ��f�h��x�cKAs�L��H}��Vr>����H~Aq��]���R��N�C`�ډk�a����y��f5�m*���F7���K�>c�ׅ��䏢����q��V����ZzᩱFD+v"����z�1��(�\��H�����x����u�����P는8�Ҵ�UFTd��l��m͢O�#�oCP}{�j�Ǧ�vt/�JWB�?@��ʋ���N�/[�J��Zs�X6i"}�T�������dy�{�<`+C�%<�k"��.�R���+6¼L~6�����hd���-"G�1��ڶ8Y�ƅW{�K_"��O#5j��|3w����u��hW�!���	�<q=��و��b'��� �]����2�\�De���#X^��p�?һ�x�M6 �oO��r@�FlVף!��hRֲ�`am&�[���g@�1��G0��p
�'�HuV��=����{���(���9Sk��$U��˯�1�����Ƚ����>�^�K/��gj��Dyf�Pto�mT�⠅�$�	��DC��~��y���B+�Y��i֢(x���+���OO0�.���騥i��$,ù��9;n��O\�T���nRX�V߆p�	��	�@��7�Yh4cؕ��TDE𭌭���,���f"E��������������� ��is��$W����<���D��A{_���n������>�xz y�
�n��h�KM)�,AG��y"�H�۫{���6p���nG����c�=��r�.��ԅ��B�%C����~y�%Q�,Pm�&m�i���6��M�±ch���~�"K6O(S#�o�u?b3Y����g i�Y��.h��3om�⿺�|�ϫ%�����]?����iL�D(�=�"������b�U!�dkB]e.6T�qT,���-�GLS���t��U�����H-����Ԃ �[����W3���/��D��
��Y���c�F���L�NǢ���o�}���p��!�7{5��Z��o�e�������:���-�dͧ�{�O�f�)x5�R�A&\�I�6c� 1f����	�[r��f˫4Qzy-����0ʦ�N�z-=+T���vv��p�aki;�U�ٔ��w��:q����\^�Z��M�ޓK<`�1c�~��������Pd)���N��=���8�S�ݏ�az��F�G�ވ��I�XJ����D��LΩ#��v�d�"S�y��Ō���	�ݔ� ब��v�ɡ}�o�>�7�"�P���S��ת����^��b�i<R$��&U��h�ؽ�Jc��Qr	�'���h�L�U���U/��_D�N\��3����탄i�?��i��k�c��*��s���F�9x��}��T�K;��?�-�+2B( ��Ҳ���g����]�,^���Ey���W�o��8��Ai�WP���"�_�n�j*��QI�Q������Io ����x������	�b���0��na\�F�W���bz��	�
�Y�$W}M��M��c�7ŦF-=�A��`d�ԗ���(��%ͪ񔀊kQ�Y� NlT�(���)��os,ug��F��*owq��?�?x���
_D7�Ss��Xʚ3 rM�n�Q���h�m��#������͞��8i5Ɏ"3O�{GX�V�X-�9��Ԃ��ɝ�],6ZS{�M��SH&�ѿ���{�Е�����L��O&Q�<���=d��ߋʣ�+�V�����_Lp*5���λ2@�D��^]�!fG�q]�ۗ�+M�,�'-f!�p���0��W�I�'-�#�e:�p�7�f� �h�I�;tW�ѷ:�'?����0�n�Z�M���\?����).�̀��)7M��/�qH��T���l�ַ+�����I��N�{�7������g�]������r`�ǫ�b�O���Q��mD�������E��r���b}�0������Cc�$�����@���5�u՟Ln�#��t Ɨ�uӖ��Z�YU�+x�T�o�C��G*�c�l��Q�O����t]�c�]7*Qa{�Q��G�C�����h0��a �{�rڑ>U�$h킢�8`��tS.u� �)9t��8_��T�)��8�{�r� ��l]���|��i��@�e�}����i�<Hwr-qw���*��1�⎱D'm�����٣"���r¬���oB=��l#���d��GpbU#�n�$�C�D�׽��K9�؎iB��M�J���q��I�GY��Ì~w$(�/�Vۗ�FR����8�F�
���-(���Z�] ��k6dQ4)�4�D�X�M��d�����Lv`h��^P+Jr#w�%�kC�"Q��D�7v%�8��B�ot�#'���#��J�q��z��x��d �����&�7�[����Gj8�=˯�N�5�g_��G�E[B��`�&װ�AO֗0�#���A�6j�����3��1̲
N��N��ݑ����l����O˗������QՓ�L24��u7#�Y�B��J9�N�|`��VH��L9;%~ڎ��|�X���,% 6�� ���z1p@j8'H�@�-�wf�����|�%�h���%���I��i;��$Ⱦ�9?S.�T���u�҅�|�C@'4^W6\r��cŘ�	���R��#���"���Fo�����G���d�x�l�]KT3����!3of\��s��O�y��ZH���O&%�"�Qu�@$q<�M11<�<C �M_5�_�U���4�ke��)��쩱�
��HM��M�_��z�nՆ^���f{N��c/Aֶik"�"?Ϭ_���-��B= ����銋R�j�c�4�<i����p9AFS-x& ����-��+R{��Ot�wc���7v[.[/���;�ik�� J�}2�D��ӜKQ����Wa��|tUZ[K�t���I�Zc��I��T�M�*�P�{:n[��g�n���)�H.k̀b3�.iiawQ�.��4�������݆ɪ�N�+{������Wi��)�3z��X���|�n������c���j6<���@�&�X)��eC�l(�A"��k~`���Bt�}O��ɖ���ϓ~ ��(�ٙQէӪ_S;HFS=�qW�s��-��Vw�bڷ��������[��JCs��`w��ᆔ	�=�H��d�-��A�(P����*�q�t-Ң!�b��lb��K�\�
,��q�&����R�D&wc��N����#�2OB
#[��JT �8C�bT����`���	�[᪫!Ђ�*���"��e����oJ�	��@18��O������7f�݋Τ�E�5��L��.�'3�8l�B���C��BWuV� �xkn����H�:�P���l��Twu�c��U�jwXck9zv ncZqE=���ikD&?(�׮�&�h.3KE�IMԋ�����8Ha\`�x{�E��a����1�g�Oh��2	Br�@���wf��q�󍔏hz�x���=��A�(����ηӨ��ƍ�=(neB�Km*������i����avu�=����鯆?��B���Gs�Փ�A����*�E�0ٺ5�P�+?���%��9,(����*Gw�M\Um�a�ToU�Qc4Y?uN�\���LT�xm�i-����O�2ב�.���zi�a6�6��)�ф3���_�)\A�=�ɱ�9��Qm0�?�k5ő��s9xl_�վvf��9���b��}� ���rV��3~��ƣ?�=2�%7�J	7\2���d6y�QjO�t�(�Ҩʱ� 6���;�OSG����!�S��T��1b�Frs���)�ō=���"0���3}^����-�O3��� ��t�1���y&HE�i�0qѴ�sߜ���)B_	��B���܀�;�D�����Mf�SWfk�a�e����r2ё�#J���e!6�����)�� �"���@����]N�W=j���\��.Rn�A������.��Ȏ8�����!Gp��q�͠s`|Re�&l�����8\�z(��"l�������)c�� v�8DSݛ�S������o��Ox��}�m�0������%�4�K�yԓ%���@���JO9~哨 ���_OK�"@�QB`��������M⬲�T�[C��.��7#'�
M� �J�.��;�N��8Hu�s��N�2w����A4	g�-W*'5�a�+�D�Z��݅��z�ژ�p�{��� W�v���͜��O��+G�x��rNV�h������+�"Yfέ���u�9�s ��8�B�����|��cV���vc�o�.�:OU��Ve�W��m�)ܨ*)^���-�&Y%�DK%�����'��K���ʑ-8�$Y�����+8��i�+�E�Q6����
B�S����Ȭ���&�˾�2y`W�6�P	0�Йyf�DUI�E<���+�F��~Qúv����eq��A�_�	���y.�
��r�k�%��X6yוL��_���X���:�_������%#�05�ٱr]2��~A���7�I�!@ƭ����:����ƹ�ࡳ2 {9�)���|KUl��� ��}���\��*@�:�ʹ��Y�=PD)w�0�/��3�V����k �5n���\��̱M=a��/��\����@I�3�A�md�+5�c��p���r���,¹�q+�X^=t�h}[�E��1�V�[���Ҽ�F� �'�w�g�cEL�u;��w�����r��h:���/:˹GX{� �ԕ�%I�B|�n���:�-h���a��z܇�$�g��P� ���Mz=��C�^-�}伽h0#/����#�'ePhbf�fE$;��u�x�5�e"1�I��@�b�>�.}�6����Ԓ�;oe�?��2�RU�$��0�%���x�y��?겅��ՖmW�^�B���=�g�M�3A�e�G*������ V�A��Ϛ\o�&\�nwa>��!�ӎhd�A�Oi���_�o�ƞ@��|@d ]C��+tʨ)�PCS"Pl+�0�U���~}ҕ/9����T		��U�`�Oo:-EM�$)�1|�(�i���ђ�эU�0���� GODk���������w�]�X¶~.lJ~b�d�4
����)g䐏�7�/<�s��\��A�
����F�s�Ȥ����Wr8 ��Τ��l�Yq�������ӕ�/Β$|��vh�+�!����K���!Z�Ϻ��=�o���`�hַ����~9R׋��u�<y`�*�[��h��з8��F�F3��o����@���D�9��qL;>>øv�h�wһ固��wݡ��+�j6���mʭ:���\����T�ˀț���=R��}�<^��9��(�ﳦ�=+����p7/�qt�"��v�/�B���/kōy]݂IF;o_����������*ox�D�s��K�7���iF>d�V���,ڠ4�A��U²�5�a��^]C8[�_�0��\H� �X̄�B��N_m8�dkL%1�X~���[�c�r���9H-�)�/��:�aa���:�QP�!��=)CB�����^ �V���x.�4P&�Ia�`֗�=��#�����N�~pg�Sܜ��Uj��}ܶ����ڰ(H 2V�Ul�i��>��e�?kK���6y�����sv| ɵ�>z�`:�N볔�,[��A�4����wy'�C��0%cQY+H��,I�A��$#;+L�(�`�UXE^5!�[-����A��
iC�c�I1#�S���n�b��p�AKً�0A���d�������
l� ��2�P/�#���WfBR<�T�cX�m.��O�����^n:AwF>��Y�~z��z>���0
�T������DIc%��4� �{��!l��A�s6(يs`��4��!	���#&r9*��ͩ��6���n��$��K�b�#"D�x�{��mB�Z��l#��;Trw4M-�Ot����Ɵ�A��"�զ�3kǿ[�k�|���Hu��*9�ؓ�� �L�:�������R�����aI�z� ���У���W59��<�u�F��\ma���@�Z�k�#��5���Y��v�]�������r�-��+�5A���ɱ�}j�a��:b����JC��~7��܊�������^Q�Q������!M|6�]c�������Iʃ�hz2���+��ݑpp�BG���%�V���5j��n-|�Z_��7�M����`�1�Ъ[P�_��y��BF3g ɏ���2�M�6����V5�zR$6M>&x��0� �j���V��M=��k��u�I&�5���F-����O��|u[�+	9Sa���ʟ:���i�a>t���<�-�h]���ϊØH@4�B�OO-�����n"2rX"Jl�o%j5�9Đ��P���TR�X���&��|���m_pR&�E��[��kFG1<WB��VZU_�r�Rgsݬa%G�������v{#u���*q^�T�e�q�6��Y�e�eo4Lp���TnM6Ϯ��'��D���H۞+�%0� p���vύr�uz��̄ͶҕYl�/ؐ}b��^��6W
�-��̿��x@�����*�'��h0��V�R�w�)0�ͧ�����U�Ѻ�EvxP߁�)�im!ICRO�?�&��뛿�MN)G� ������o�e�**��n���w{�SE����+�9�X�m��b���B���㬲`S��ׂL�@r�Jѝw��s�X�|�KJ�@�q�ok��ɚ��4"�E�F��W�.�l���X�d'��U��/8K��\q!��H��=��~�c+YzsHcQ����ua�΁2Ge�_�>�u��NB(��T_�QV�6�ϱްtӑ��oM��l`L �q>�-*BF��e8���M��>:�sw����	W����3�0מ.�_� eM/��x��Z�t��Θ^?d[����M��:��A�����Bq%C�E>!��tQd���gk�7�3%~uY�:��iX'^�ݴ|՛�H���ȁ�D#��{�_�C98๩M$ -_���F���սp�Bpl���l���������܄�ٲ21���"wvK��Uqٜ�P&!w&���At�67�d^���z��o��|4j�Ҙ~b@���4�������vA�V�*�����W�H{�`��w�:�Ëh��� u��%Q�;6�| �1ck���&^�[ʙw���y��&�g��haM^8
\�G�J��(��Ǆ�M� ��Gd�&��t8�h"�Aqx�q�l��t�4�{
u�_��f��	5��) �[I��(G�Nj@�r����a�u�ȇ #�8�p	a�Q		L�Ah�㕮=>R����=�$�����3v`�8z("O�ƈ���	�c�1���G���e%�8�ƭ�ƍ��:�~Y<��S:�T3�}	�ֵr���(�m��{��M�Ǖ��~�7�8{��i�Sr'g�!��U�u�j@D���Nϥ��W&'4�|(?>D-Uqu�L��lH2�re?��9b��Ξ�dK�P��WK�[o1��R��|I�u.�B"�����o��{!�b��S���8�G��b��l�í}춲Y	c��1�ІVT�98=RI�^����o��
��;p�e��5���;��)~��ܸ���{��_��U��AU5Fa_å!ֿ�ԷT%n�9��x5���Ȇ�y�]���}�:;*��_���Gنɋ7�ܸx����
�����՚���פ%�O��k8��)�+�Y��	��Hֵ�nH0j�l�)�*ͤѸR�.�8Js	�����s˸��y&�6$��1�t?ќ�8}�=��Y�b�r.��ҭt�������̾��]��7;��<!�c��FC�ik�����p�+! ~e�ҟ@m���B�+pkτ�R*]�N.⠳�:<����O	�	�����P;�ڦ�q:Cu�l����l>��h���.�O���M�u�U��;��޹���*�Nr��ɵbq�`���u'�XYoh�n�V�����)�ld������|>}��D�zfa|5�[n��U6g�~����Dz�Q�i�$dRߝ�6�51)t�;|�{�s��4v��$')IA�G���}1W�z�FmT{��u#�����`1q�C#��i!�������/�	e�T	x �=-��$�M8.e�c���&jN�ԏXHM -�	Iw�!̅RE�MB�ǯ�#�����(���<�k�d���VN!��E���ټ��\�ʥ����B�I8������u�s���d�ue1��댏ٷ.)�	�	:�L�n=[�S"�	�=�z��)�{1��6᎑�E?�^R�sc�a�W̬�8D[N#���yx�n6,�Bo���7{���?k^��N(w)UL��M��R�99NěE�@���2���V�w+�پIkW��2H�|`�E%O�J0�)� �3sW���p�DW�t_�,"���!"un�kJLb��^�s�aWݽ{ͻ��l������=��g�"��M�W&je�4��(o��%DJ�%����M`�ѥ�\x]l!Urة,W/#d�!��%v��B��N1��o�[#0�NH��|L
��� �[�[����^�4f�YM:A��c���7 ��.w8/w8I]�.@b����\�Y_T��W�����6q�S?+�GyǭOqe-�˗08���Fv�@A�nD�_�_��G�_��?�p�K��׋�	���s�P��NDֲ^:lyKZ
9������݇ƴ(�{�ك�䀟va�V�jj���gW� N����澈(�F�I
�y Ԥjj����fb���i�� �p;�Q��>D@h��֩�b'�Ez3���HDe�u^�Y��`3���,��>OH.o���~��J�!�M ���4k��Ɓ��Ȏ��aĲwfY\��6Liz��/�d��=7S�8��~]#O÷0V�����\d�]% ��}�TN-O���[�E�#����&�T9*���]^���H4ϥ�;y0�~�s��qH�"#��(�ħ-��2'j�yKp} �9:�n���z�;Qε3��{=\g��5���x!)�_���@^h/�"Dv��|���gL��2��ְ��.�����+���Yћ�$�F9E^7C�+߂l��nn6+tG���i�Q+<���X�Rͼd��^��~ (3?�ي��1S~?��w�%�x$
�˼��T���T�*��*İ[5�!b�Ț�e��=L�AF"���8E[g�f�e��,ŏ.����Xd�#�[bm	ȃ#�ϛ�5%���Q�(?�ֈ�D_U@�:U��|U�݄| .l�=��5�;���`XI�?*HB��v������_![7�:�ۂ:��R��"��&�^,�p�0�el@���,+Y(W��[GW|x��>M��s�+o�u^�q�5~���p�n��p�0��O���r���T����Ǝ̳�"�j1�Sa^a����m$��p)�}=P5���8N����X��yY�w�=���FP	N��H��H���7��O}�o��to�;L��¯!�gUw����(�ɵQ�(�7£��NP)K��OP&������;�37�2�� ���F<?XO���Ts�1�J�$p2`���fK�4�f<��wṿ.-^q��8���d���r��(�h*��!�v1p��/�K�E=��0�<�h�-�N�@7^��k��>�g�u�V��#{��*N��%�-6_Ÿ�Hţ�"H��d�1Ķ�!�Rj',��U��pK(��+��-w(���<@�o�"祓_y72�UK���﷬s9�D���ag�Tv-sT_��A2���FF�5w#^ݬ��5�*�OĲ�s��q��<r1L|RG�����~�&�d�A���JOj�i��#��R���o)K,�6E}��ﳗ�T�H�W��;�䴁��	Io[���w5L�ZN.���8{�z3�;~%��ISP}�/
�<�`?��%�H��Q�.��԰ģ�$�"#u����y�rl���&�Ydr��<׳o��|�KaX�z����գ<I��Rj��8���n �8�(�u�O�G��Fe�D��6[������1���R����<����� D�|A�®XV0��g��
8d+ۼm!X�ʱ%>i�Z����S��s�'b�I�'����E����b��Ƞ������lt5�����^�c��JB��s���������-,&4ԶF�<m{��<d@�u�O�X��l�')������rkS���]Q�G�g�u�-����o{�NG147v��A���o�x#_:�j���6o:�Ƶ�&���n�n��e�H�+�Ŭ��رtD����Ǻ��i07��Fy9;`�x%1�f�v���7��@$��a	9�bۈ|���՚�!��|2^��f�J���# 3���ޒ/��DwaQo�PF���"Gt�t�q1mNhİ
������F��k	y"Um�͍企��%�L����g��ka����tF7�U6R�d؏@�bE�Y��~���}BJ�T`Hm���@�c����<%�r}�2VV�w�g����	��U��^����͇���YVd-姰��n�Z�Mr�Hr��~ӳ�۲4�G���RK+��s`&�.�I�>��㼉�`/* l`�/T;/��_�O�Sp�m�z���ç	�y�0Oj�
�·��"�R����Ss�E�z7*SF?J��n�П�&��U�Mi����}^��\ns�K��/R���d�5Z�4!9��aDWX�v��~����ʥЍ|�a���)�G��D��Tx�<m|�'����	�^BWF@�m)>H8ǽ`�~�s]{@�%� /�6q!��5׎Z]��.�n���F	?�\�Q@r_}N�� �2����#�Z�P�����?��gZk�,�K�- ��8�V�CE��� ɿp�#o�~�n���l�/r9��w01��F�F.(�3ؘ� ��_�>�^�H�B�L�?�}��kE�{ē�G��[�%K���D9��Z+��;;�zD�Mj1�tv�ꢒ0E!���^���25ӄ��ۉ�����;�N�A�}���^��x�Q+���/@��9+��cB0��Օ��{d��H��0?;)n�L��u\ � W�7�_U�]'"tv�EH��P)?e�y��۾��B覠"t=�2��{/z�-�L�^�j�QMN��l�c�RE��~��-����sa�0<j�ǣ������9DDQ16�;��g�<ât>Us��P3��j(��8,+²\Q�.���0��|�~�=�e>��OQ�z�+$��31��D��H^���p�
�w�@U�^�?s��"���Y!3�5�t�[q���˲qP��-�����8�>�+�z���
�c8	�qb}��%^u��g�p��d�{W\�f��|�1�nX�C&w�hδ� ��
׭��#Y�?��_�\���V�vtV���i[����{�ERK﬷N��A�jcAX��n�G.��Xbj�VY�~�Vب���:Q��
�w:>��E��ә�e�����>?k�g�tI�E����fId�wPoi��X�]�`�;׶��j�s�(��mx�Մo�I
+6i+Շ�t�]��jY�mv�7T;X�ct6Ɖj�ƫ�}�[s������J��`�|�p!⠓
e���vf�����yZ4���_�c{�j~���2 �E�Ew:��g��8�º�Ӟ��R�u��X�7-��=T/�}��1۶O
�%�m<9�HVX(��4�w�բ�5�f�>J=py'~��)��cMb��G5�k��`�b2��D��O4�UL�'H��Y�(�e�Ǟ�]�:e&4�-�|bN�+�0���9-g+�������~��j�17�GX��'�-F .��f����O�;g���aF5��'�,�d���M9S��R�x�Hd�b�5��Z�9�{"��p��&vq�>�ež��q`X�e�i�'�i�p�<&gd�F9����E.������(K0MY**�Έ~#�]R�D��/�s�)woI@!A���c�u�:��[�׭��8�mZJ��?�%	l��6���J�c����s�о�l���0�×t��>b��y��d�L���2���i��m?�Z
�E�[����@�֝*��5a@iYо�c8�E�ؚ��S�:��dL�2	C�/E�P]bj�$�3�ۥ���(�o0柊p�ȡu��n?�]��S��.xN�����L"<p���P����|�j:��~��$���'_u�m���P��e��;��R����߸�'�UA��>*���TŇ��U�Oc��5թ'm��Y�5�ߧ/04�%%
���n�4�^�W5A�]�f�|�߷Pz�)�3]�ם�g��i�9)]OWR �3����;�8ȯ����wT%,w[\���/��T�:����pSVV8�!՞@��l�Dƈ�O'� h'�D·Z��t�l�3�@xF�c
[���"X	�7Ӂq�b.�et������v�p;�,|�ܱ<��z��f=��%��V�]��a��E�ǻ��+ުv�wq�<Foۑ���""�ډ�|�w��T)��}M<�Ig��}Ⱦ#Pk$�`B�A$�6�R@L,�c`����񎢔��H�&�Э��J�_��o-t�}?�6v��u9�y�~�����(��`����#_�_��Pn)9�|��c���h��=��0&t���\p��Pa9u���kT"�1w�*R-�0����K�MQ�&Àk!Q�E�a(|�Adh��`��b�Z�Q��",!x�{#� µ~��p�6h�V��u����qOu�s劘�At, ��h��!J�[t�eMf?^�mQ�T��`�dw!0�k�5�� Z٠�F�s��2Ng��;�qT�#�˭�ݖQ�<>�/w%/[y4l�M�/b�VwH�[`J5G�=����6+]��=��ᠸ�P����R(�D_n�;���An̖J���U���b4U�t�>��Q�p&6��C⌤o�^9����,�
�u��iv"#[�0�i��s��>��[
���rq~J��`��W?�F,�[��6�Y��J�_���Q�M�刃O"��g4!R��C�5��]�Ww�$[l�0�N�����/csԕ��)=�-;q�\�����M��`ˈ:�	qG����3/�8i�ʼVy[ʰ>!	ŷ�@�G�'賘��.���g�q�,2&��y�'����e�G���BDsC>��X����4�I�t��Qʽ�'$����K:H'W*Vi��?�ښ�Z���2#��\��b�/W�]���I���$���u�3�ԍ�!�����JSx���\�}�P�+FL�PZ`�O�?���֘��Lf���̼�j����]�g' ��CC�X�X�0zLb ���"C����}w��)�"7je����j���م��+����P�+;�aUq2���ϥ[��!��z��Ec���"�zmr�wJ^ۋL�m���Y��"�#�}�C�8�3�M pC\7?^�A��0�-�K�f�zzL	�)R�$@�^k�lp�y��_�sПF�ek�SY��˽�ßk*��/����4l���R2�;�,�$�Db�K��ʌ/�<<�9/-ڹ����c:%H}9͆9��������MAe�0����8��K�P;�Ug�A��dM\k%~'v=?���6RN��X�~�{k{:�׼%�z��=0|��=5t�r���7!����m�.R�_t����\n�!oSg8�m<[½���B!�*��*ҫ/�l� XI�^uޜ+�♧���$����[j?�4�68
��R��=����0_�HGK��n�G�W	�*ͩ����(u��u>sY�i8�p�W�!��@}]Hߨvj���җط�_��vxp>}�������[��L�0F�i�.�S(�E�'�$�-����߶rl��*vn��^�U,�� {�����t���?'�e��� \�a������@�~� �޵���af��=ng�FRU'�7x����v�^5ˣ���cT�$H1���҉���d�7�f��C��cy$&8�D�LܗV���}��m��G5$�A�5��Lۉ�h�2�+*���M��'i�Ch�@��l�Ome�p����T.�C��RlB���gq�"��*�tr�`�[���+�!v@sR�|?j�A�x)#���܁��m�3k�y-�:��G��5t������|�ʻ�. �":\��lw�|С�}؛٪�q�u���-�`��;��W�
+~[���7>݈t�h��N"Dc��a(*ko�~��x���Yhœ1Ԃ�Ŋ��.`b��rCͅ�O(�]���t6���ʹ#g�
�ga��<T����y�-f|s���!��z���ˈ�_�}���62%-=1�:jѣ��e3Κ��;Bpp�s$��ɪ�X��3]Q�(��'{�Z�#M�ߚ�L��;�	P����[�v�!'�#[ H��K��؄:���&��\�^j���I1�J���/���eD���\��|������_��GZ�p�'�VPh���x?{Ix�p��?ު�{l�[�S=w����ഛ^��~qp�,8ZO�y\���Ũ?��\�J ��H��"m�Og�֓:�n��/4���sJ����Vf�ԃ0��L���mb�|j��:��;u����RX]�����m:HX�&e���Ȣ1�a��⼣�)�i,�E�gݷ�!6g+�)���'���Rx��V�0��Ge8�]X�������gX�n?�=����Nh)��	 ��k3V��u�����a�?f���-�4!�*����7n��g�Pq�/<�0���G#�����b��ǩ|�0@�ZC�`��hӧ��o����J��.�q�Uw�@���s����~M��!�o�
Q�b��R���-���C�JٔYO�x흎�S\�f�?�������3��������Ґ�Jd�jW�ec:���E1�iR	O���$K���׻��j��K�����a�~�#H�]}U�m��x�jwʴ�;]����oӛ'J�J~r�.�Q����Ș<��H�wAU���1q�D]�@��u��ɧAꢀ\0����=�/�E����/x��TiۧH
nڳB`�P����2s\ OX
�L�`�*t�l�#0���E��I ���
�}B�q��p3'�Ƒ�`lT�Y8pM���8���(�9�Ep�4�4�k1gv��R�����!8������f� �Y���٧:ةsy��^(��e�>�ZL3�TV(�	mkV٬l֮Ǽ���)�p��E�
�k�j�)�����5��j�/�1p��T{������5�i^T����9�O�s؈�`��Ls"�`�-7�]�]�È�U>�uf�.yQqs��e��k��|��b[u;�ŀ�nUCt�|i��I�X,��s�3}�a���ŧi6�u5Xl�;V�X2�'��%1ğU"�zrӺ��8	����E�XR�����ή�:4n]D�{}��v�؀��`H�b"�ɘ0��U�%�����1���Uފݞ������-���!-~�����%�zp2�c8�?MD7� �c?w�zs�g�=�̋L�
�M�TvZ(	L�;+�&#��`�6������f�"�M��>��{����00l�����>=x�rE�[3��ۘ0"0ec�G�����JU-q�	��Θ��5L7�S��/���II�sAl��tW�n��.�ӌ��t�l�d<�_�,�I�����ֱ�����?�(rV�&�9 óJ�|�z�Va@����f���#�P�Y���7��(:��;�1`kNY�
���v�0!����۬c�,��
e�M�<Ww�x��+���3R�SWt~c�s�̾�z�H�q���`�)Ē(�
��W�?d�}���W�x�a@4��K����1�9�j��G�"�r�+><�@4L��j���k=o�����H���s��N\�r?����<��מR��.9PKPX����!m� ����Я��m(E���,`z��= o+�3��p�O^(��^���S�b�ߗ�}
e��ꩱ�"�@M�����-�$�`2j�6zU�7�b�=V.lȩ�{�Q�9� ˷@�̀r�$dh�n���f<L�?�!�&�s�y�"�L��t>)݂��#	L�k��<Pg�d�uFȤz�9�����6Ęº���9܅q�S���DK$�����&'��~��2a��4�ru �5wGƒVQ�:�w���a�?����o��%�VpR�phE*�Sg��=èdU��+���B]������$j�d�A���fu��@�(���Y^���y  �z��ՏPR����}V�,,C X������W�㎭�G���r2�R�O�R�~�t�LVE��
�0Q}kd�V���/�r���D���f.�m��&?-!�C���K�y�F�)^�QѬ��v,����-Y���J��-��t�f�Mx�$K���w�Zˣ�W8�ڟ��M��7;1T�m(d��26F;{	�7-��{I��o�>�r[1��bsB&��Ա��#���Z�]G��iZ��=z�i[ c�&��t�&����4~{]n�&~�l�f*�2_zwm񶽏9^�Ι�9���,��a�S��~_��R���"��0dH�]�~��� 9F���ˬ�	��tm��!�P�mE5�n���$�z�V�Z�Z3���{84Ѷk�}�n�G�� zU��ξ$%��8�7�X�=#������`�sl�@�El�y��yx.).\Vz����J���)�4鉥β1v�����a3�f��G�c֤�l�#
Ջ)���!�xa�1��w"�{<�\��V&!���/��*d��-|�i�	S0e/���s�	�����%�Љ/����䙽í�M9ᅎ�.e��Q��-�oL��%��!"{���W�DUH�gX���g��	~��O���y��nm��?���g�G��^e)���,����!����I2��'Cٔ�m��!����P%�´�=�*9�/�5��Dp���q~���Կӡ5�P��W��5�=�W��� �X�1:j�D�N�X��/U&��G�`�V�@��$яt�tzq�B'�a���.���C�U��5�
��KN��p?$���bv+_J0�*o'PZ��Ɍz���A�ϡ�����4���ި'�d�o����p����q:+#	��P����C.�Z��i�Q K`����8V�+w|;`�#'�xpE��4�l��o��X%h�O~�,�۴>r�� ZL�����:˅m���BA`�^D��p�EL�)����!��I�lVK��2<���3�#̙����o<���lY��_�����FLh(�Z`�@�R`AF���Er ӭ1܊�	H�sE���BsER6�*k�ʃ�Z/?����H���=�0�I�]�|%��ߞ����-��H�^%��1j��) ��"���﬏?Bz�Ze�z�b6V��P���� �6g�&t�),c�������oCZ�i�o��F�@J�o&G�� �i1���:>/��q`Gj&zI���Z��0����Fg��ȟ��x�؉��b�����$"�@N�P�)��4���S�۠>uC�L8����A�-�5&.�q ­��ٛ�"�=�j�P�Y��:ߘ��g��M?$��Յ� ~l��@4Il~/��[.�7�*/`�圶e) ��<^g �k�w�*H���x��2��qj�ѺA��ȿn�����5A�3�J�ױ�c�J��"m�Ω*�/������3fJu�9y��K?��l���#"W��h���*/2�Sq@�%�PjbST6r��ű�w���D���~wO,��xN4��0h�2�4��
c��,M�Ð5�����weۢ3��;)0����Y��8jTp/�D�xo�� �r���`͐�̆wA����6�`$|۸��W��$%��>���\���Mg>��sY �ig���
U�}��pԦ<��1>��W�{�WDT��w�C�?b��5��a�H���,<o�E�	�&�Vkڜ�b�w�K� B���L�Ϗ���$[Ɏ"5K@�t����P�f���6c����K`�?�=��랱lW�G��S�7��$�:0ȫ��So���Ω�E�o�u��|H�!%�M��0�����!<v[C�����D���ל㄁dU��3U�h�:��jA������N���PBIn�.�S�p�X	EE�_�G&��A�o���,+-4{��3X��Q�njN�r%+�n�o��qEε<��X���	��DRm�A���XU$�hcj\�"�RH@�~$7�;�Ւ"{�M��� ����w��K�-�~��r0�w�[��n�ܬ('��k��*�� 8bn��­�7��٠�P9�7m�M&1��H��a�ݻu�A�Ҫ(q�N�zkwݱt�0Y8�JŶE��#�u.��\�~�Nk;�<�?h\����Fӏ%8x�X���ł�f����\YN�O�F����Z�j��u���;G�㞱�I;d�f�/A<�12M��^�#�h�۬!�3P���Y�UH$�ڦ��V�1��D]ι#gb2��y5F	;��|��aj�&j3�eKN�ِ� )�,��g��RѷZ4Hjs���32����+٭�r��i����U D��!W��%�o�S.ƿ��� F<[ǔ����f���NgUu�J�׶+�+'����1��tiTE��{T1� ,������S�$N���b�S<�c1@ �r�`|!L���K7?{���������HPm��9b�W'�A�S�vhr#dEb��KI]�O��!Y.�x^��|"��a7�᥮�<�eq���u��6)�Ѻ���uT�o�c-���L��9��qWDc�g�5EvL�I@dn�p�G�s+ ��+)J�#C��Q�p��}K<.�(ѭ?&�4�0�H��	�㆟+��k0d�� �G�B\���*���;���Á�32�V�l7�)��25l�R��aX��ԗ�=�S���������X��q�}�ĸ	�=u$;�`�V����6ni:�c^�`s
4�������w����p�\�K�Ms�2�[;�����O��;zk � Vu�^�Vʕ������dU�SI�C�=H�i��'�~~��϶|��ތ"e���S^�pp�5o]V^Y�o~�SHk�|�����Y����Ϻ&]��&P �y�5K��U�Z�����ަ� �����(K�!��m�a�%��>L\9f��<�p|�J7�vᤀ�T��^?M"0�<@���6���#��kJ����W� ����ȑ�U��_�J��l��	"�}��p���i?6E"�E��E\�F��b��
]�����F:w��r��
�eޚ ���I�y
���qu��|a>�bNJM`�]��{J,��f�Lb��C�kd����,� 6���;�����8Q���Q�R����Q{���z�)�%�ab����Z����m$$����*A�p�[�_���cy��4e�8��1�#�������0��q��n�A���7��M�|B.W�.v��B����{r?�9kĩ�)���>eW E��L��D'�J���>np��*�U�DWi$��U�Ҥ�w�@�#�C��V���Q�Ӈ���1鈜+}�o9��?�qY��<!��p�R�^�~$NE3�9']ĺ�Jfr����`V���ٵw�`�^<�×���$c�O�=$}�Y `�{�z!���iZC��n	�~���Tk��� ��Q�\�n3|���JD���Yvs��#��c::����p�2z�\W3��]�
�Gf����$�b�V�râ�Y�T �@���tz}��J�fG��d�<�-Ĩg�Bt�{]c��8)��y�E�l��Q� �H�v���*��;���ؒ#6�x*�볊A�88�}-�� ,�_Y�L�g���W->u�7����̄V�v_}�7ʕ����C�2-i�h�|������5�`�1��S6D��{G������:�P�?ہ�hU}��� ��S����upp2;��*�i�\qbY�_hƓ�WwscnK���9t����Ԗ��}����f�g�Rџ�Z��H]��>Q7M�d�b�>����t�*��:
�>9��M����9pE�i��p�?�MX���N9�7z�$���,�hB�z<D�������[�X4~�B�AՅ-���~�\�W-���N�|�{r�z�\�}�����k1Q���ȱȾ�������9ᠨK3.�\�\UϤvV�AY�7����V�c:-y���/�B�Y�1�o��&�!��Z�@��0��m+�����B0����~7m
��K�.ۮ�l�}�I\$7�P��'�0���6j@9��?�N.D�����d���_���2�	���]KG���Gar�]�?|�_WoN^�<�P�d�]'~�܄����Ǆ馆��	�����PE��k�����B�I��ڂ����N
��<��ub��Y�6p�B�}����^/�O��a����p��$Έ��ٹ��d�>髹�l�w���ʑ��|�����ʶfb���N�^Q��^X��� �t�)�\P vĖc<�$7<�5Y�/���5y���@yuz��W�%�&�r���\�8R��(���Ѡ67v^��>�7��[�{f~���,���;��KD���Ҫ�8d�/DP�D�JO+$7�0�!}��s05b4:�`V��=��ȷ��z&���T�}+-��[�޲���x��ѓ��6VFuo�M��=��\�1C�,=,�+WbtS�^;�51(ɶ�f��3�R�)��bQ������D���K��p�b��w2;�U?~���{��Gb��9WP��M����D���v�����:��ժllb5�2�%*5���Ӣ�1{��i���9_5���Ü	X�klp�@zaG��;��ڌw�M<7݃#�b��/�
�`����T�Z��s
W�V����څ6	F�OTEI�Ё� Jl����l�'�qp�M�j�t�����V��N���^Q��r㇠�'~=�{yc�5�������]�4�Pf�P?L�5��r�y��B�w���:�o�:���¯zEZ�s(=�H�?�U�Ƞ"�bO��Ŕ��8 �u�c@���NeΖ�Sةv⹣�Ɋg�s4e��k�a�N�F��,b2?���dA��vl�Q��U�UH�Ű�Px���n��:��)><�������t;Q�!Ѻ�ܣ�KX���� �$P��i����7��:����&q�ic	f�LJ��DAb7���������Y|�/5}��^�t�ܛ��	&L��s�>��t����FLMs�z6�ǓT{{�����|Y�]�G�1������� lY ������;�Qh����\8Lջ�ҝv��V�m_Є�]��»2�F�x:�ԼО�0����"ƬM4dR�K�Z�*��a�����m�Ǡb������_��5b���j��W��_����́�T\��"r�QVI��֔�yrg,��4��8�#N���b+{q ����*���z���
񃛊<�̛�F�j+Y�A��S�n�x��S�s�V)������|���_��>�:"}FUj*/2k5+ğ>b���]��v�Q�8��p�F�t�m�}����_��@PV���;������꣤E�T��`6�� ��-d
�ߎ8Gn���ʞK�����Ji��ʛ�C��do���zx�̸
�C�o�"V�	�ˊa����j@J/��~Y]p5�`�;ko��i��c��(b�3�e�G2��|���>#	���~�z�"��olFy����fi��2�N/�3E����l���L�N��W=����}n�L�YE�5	�e 늇�L_�H'.���L:�Ҟ���V���&2Q�4*���wnT�u�;�Ѿ�9l�("L��G�C�-�}c��������4Bڬ����+�[l�.N��0X$�+�^�t�U�SzƦ�:�=�vg�E��W��XF`Хsl8~����������{
\߿H�,9<Jo���'*I�c����v(go^;R�#����2*B?^���p�Υx��Q�.2<��ãk�c����� �*q�$�20X���ǲ�r�#�s��9mNs��/=�{7pR��(�Z�ι�[p�v����o*�Jͪ(˝����Ms�:$�t��G���&��)ϧ�A����7�� X���I@��&��)��;�L���o� ���1J���*a#%o"��-��T���e��d�i���a�ǜ�.B����[j�x��?�9����.���:.���h���ϷCE�߱YvF�$`��	���B�@w?H�T�S��q��ّ�r�AD���(�;k���B�	#Ѿ!�7�^�)���&o��m��2Sу ܔ�/�0i�8�ob~�w�]�~ji���� �ȣA3����u�n�Qx�W^�%��#q7�U�]P��O�Q�R���!H͡ċ�T��u`�&�2��C-T�h�����3_�
��x���������3G��1���jl�N�V��+쑸y/�ш����)Mf��/`�ο[�^)(�E]�P�.����	��6��	B�
�G�k��o�!�ẋS���I�Tt��H�H�b����jέ�Om�E�� ���L�Ok����g,��N<;��!$^�\�u��,��V�ߌ=:Ն&;CM���q���M��ļS��.H��$K�S���P<E++�4��T�i���^kl�@��r7�`�Ib�I�'b3��;���7/g�8=�?�.[��}��l �*1��
#j���Cg����_��b��
4O'��� W���E��֮�{jȭM�3�|��<�1�`Ԃ�)ENZ�đ\F8�����2#��8�	�̊��SK�m8�γA��\��-��6t7Ӯ��hx;gS��o�
���b�O��y�d,�U���r�s�'7=�3�5�N:�y��cz~-Ӕ1��4���ak�@#C0���mׂU�@���H,Ɂ�kӸ�D\of�B�} ��%0����o�7;��΀K9+i�p��C+��HH��I��CO
$)����=�\�`7S�ξ��5r�w�/c��n�_g�QT2��*ߋ�C�׆���\.~��=k�r����p�Vc��&gX0.+�v7|�����H�2��*p����	cE)��~F&�}�.���q� ���-A���0�"���~��ӧ.����\�)��=�-{�J�hn����E�y[�u�O[��b�o�nWBa$���J�/����t�� Ԍ�,y=��oX�[@��2��$���o�7�hP��;T�*�wbY���Py�,�^��a�0������U��W�dJ�$駧	<ߦ��f�~QR�:KF5���gl��	�)�����ƾ�/:iYz��ў	b�28��ϝ��7��L�D�M:�Y��92�΂����)O�*��E�y��U��#���#x:=�$�g�/��-��qz�rOf�}�$;s��C�+�O���uN�g������L+'�P�xǬW��?͢.���17s게ٜ�zx[�k�@U�N톋��r�jv}N�U���f�t�	��BMOO'�C�\Ր�/������1��K���2(ʉ�|�a>��z��	�H��_-0��	��h����x�CT��ɩl`/ea�#�<�w�X=y��}�?r:���d^���5	�M��T�-0��*K�pK��c�·3�����)GuZ���.�,9z�t��Ŵ���$9q�0��x�G/&7�3:m- ��E$��}F���sv�7jӚ���zQ�b���3�e`Y�q�g��v�
�0�ȩ�l(FBz�{L:-}!�CK^g����4<��xQ@�H��]���j�P���J�e�@�%��x�=B]�ny��#)�*���5�pگ��b���:.���fFkr��I�b�XA}	@����[`i�c	n�|/��5G���鎥����e%���0Rj��B%��e3����I+�vP�E��%޲� �/#�H�X�䕳��ѷ,�-�(_�f�bQA�PfI��V�A a#�<�&2�t�{}i~��p�IɌ��ܸ5��Zr�,�*�����O�����n*��q��)�&��W_����t���Pe��c����\D��&�~��q�`�&B��W�:��p�P���l.�I��JΧ�7���}h������`�.3dJ�{��Q�n�Σ��r�g���F��ς��w`�%$���B�o�C�ZѦ$�⭷#��j�9R4^﹍��BS?�e}��i�����������J�h�8�͋-���od���ȩ�9�L���	z&���
�J�u9�N	����Gow�4�X�eus�A�5��Qo��q�G<r�u)�Z�^�0�ULМ�O>�;M�w��i���$fL��ݦ$��(a�z穃�ah����b��f�;
���6*u
qC� iU�|�>�$�hy�\&�ȶ� i:�/�X�:�� ��F:.�N*���$��g���u��!k,yi�~�H.LP:�J)Ŷ���@������w#�F��n�\̶��@8:��~��>I�'i�ӻ��|��;�n�����*D��b�j�ܛ����=M�11��Y��s��+.��0Db�s��V��6pD;�;ؙ`TpV��zp�%Kb��7�JQ�xXy���q��� �j��D��(,�Y*�{�Pˎ����z��PuWv�(wY�Dy�16�T#�RX�^��q����`�#����13��&(!�=N����E ������qNhտ@�c5��>�#�Ӷ���e��g����:�m<J��x�"�������C�;ɉ�z_�Oһ��&|�w�:h��̼���9�������UlC��z�ܗ3��i�+s��iw̺0�1�y@w�1��~J�;�c���QQLL.P��1z��P�Q��=X��V0�q��_:{0�5���|(�9s�7��.�J�s��C�nB��'�0Q�����̓��a�znl��`ЮOe����vF�~�ǝ�2�K�h"Kډ���<�c�6P5A��5K0�u�5��8�&_���Kɢ(�Hp}��)���<�� ��P-�\r�����`��۫�"� p�G�Y����X�����d6����S�}(o�w=��݃�z;%��kt���b����潇펷I�V��q��-�e<)��kX$��\O���kc�r��VQ���P���5yG�57��R�ቚ�_a�\��bq���'�&��P�:w����jk����	#(p��\�:�3������C��i,�@Vj���゗s3�L���M3�� oE�Uk���Z�(rS�7t��Μ�vq��i�<���.�� Iɟ�3����|��[��*��Q�����Qm�6�'ԡ-�h�8�Kk��FV��V��8u��@b�D_l!�sݾ��3��j�3P��2x{7X\M[�OG�g9mX�W�a��p�^�Ѥ���|��b��ҙ��2[1��Ƌ{�Mu>%ed~��]x+��~���n�Խ����|(-)D�RDq��e��������P=pS���0TC+@�h�"� 1��yJq�b��Et�� 
��LI�	�Nݞ�ځb.���_,&獽_v��ᶄ��� �Q�(/<.F��kKSssfaR7����׃+�c3��!߆�6Z�湞"�3%r<�8���۲�,6�Y\a��5/?��S�R�5c�!����'�8��/4O���Po�����CNGi={_�4��'�܊���R!��Y���^V�k�`5Y*@s�mF4c%txqt���`�����o�e#���D��0�b<�P'�t%Lo�9v��֫�pߧ��H�c{��檨�l#�鑟S�-'݇�q�6Z�҂�S��@~۸�o��<���@/�¸T��|���Gu)�����>^������[�r����6X��D@p�]$�G�ɥm	��Il%X�4�?>lO%�xt��9Ak���_i;a���<{�G���^��-8������B���o����+ J?��=���
�*-zD�1ҟ``���^8����.�iW���x���ٔ�s���XQ��>EB�X�Ӹ��^��-�u=l҇iu����;1��j�qaB�b��g�5��a�yL��N�pl���-H�X��E��X���L#
*z+]�r����zq|�p��
�s��j;�.sEJ]���� ��|�{��o$�IG�m����P=��۠^2%?��R�.~���O�#��H����Kh���̸֑�$6�W����*f��g�<��-��XQ�'�0ұ$���k�&>���Q�>�v -�jK�̙>�L�����m�
�ޢ3��z ε��p��r�����yY�bx�]�v<�ݖ(��.�M��X�	,K�1<�|{�y�z��#f�US���a}��C��^ J��q |o��G�@��L�i��$C�8�|!zs)Xm�Ч_�.?/ ���_4�_��RG�V{�����,��J���y�s�p�$n6 �(<��y$e������:X���Fe���K�V}��@4�0{\�0|u�B��R?��C ���i���(�QXq�5����͍6�`�7<��C��o����ă-�w��@����CA����,Iv�~g�w�y�c�߼B���i߁_:}��D�@W^����4�!��Z~�����1���ۃ�$��,=`7]���xi� ��[<9�wj�}��]%�zH���=c8m\yD��U���y��t�/>Ն',Ě������~O���-/� ���ď�J�ҥ�꒧(l��f��*�/P�}���V� 7J�KWm�����$0�d��h��O̙�9~�8�P�;�#�*K��w6��h��ȕ��)��{��1�Up揸�҈�$&1NmT4��\����E=��\ա�&<OH�v.iLEh�j!\k���ڂ����`���U`�t*����5�jc��������Y2����ŤW����3j�$�	o$ܭrC�Ff�	�T��[ph�z0וq�d&Rx��{j�ʄL�{c����&z'�w��`����ޑ�X���_rC�*<��C{#�ȳ��f-���{���%L�Ȉ��g�q˟�����f�FLl$1�g�M���!Ə�ʹ���`��8\M�4s��[��Ȑ�o2Q}8^@�O�,ޥ�hހ&��"Lиdy�n�?�ط_�u�'Y
��R����	�m[u���mv�����R����UU������4�fzLE�T������o3K_�ճ����ɚ�1E4MHe�ID�g���g>���9!�x&�%��Ѧ�S�y>ny2ڲ8�V!���6�ƫ�oj>f��5�׾3�(�4�8��	2xEޡ��-Q��_D�+�s,j�@{p�*�	�J;���X�,�I���~#�O	u�x�k�-�<����Z]!��n7�쇑������n�88��j������� ����P.p������������h�i�?�Ꚉ��v�<"8��O��<��i
���6�q�s�u��0���h�e���Q�>j�+2�c1�8�X�9H�*�$I���r�����>$�3aW�2��i� ��z�/Q4���\]%�{1(���p+ ��}��F���#���]UE�E�2�ע`j9EC��k�%�g�͘Bٵ.�$�`�\I�e"�Ȯ���,՟,�M�ʆ�U�f,.As�R�/�6�����W�	Ep�,�뫒��qGqf>m��6g��E��]�c��2#'r̲!��P����������nr^�6������|���k�&S��?	��Z��S�*["bR��:��	��	��ʪ��\'��fjؘ>+}�f�.5��v���r�,���_��GZ֥�.r�x��ɥ�p1��mUs�ʅ��!��s% �6~�!GX������{�eګ7e�%���x8}���75�TMMJ�a���-�q�ny����Zs���l�]-�(�}غ��I���(�eq�B31B��D��>ƙ��(.3��=#�Z_�i�B
m����RIcR ��:M�
��b�'��Pv�L9��@�{X��)�g�ِo��J]Je��זݣB���[*�퉕߰  �'H�EX���O�Ȟ\*J*�Υ��no��pݡ
6�N4I��;_"Q�0F���"�?�.�[�.{н� ��e���p>
�D��gH�q�2�KJs����;3cÂ[1}�C��Os�ԃ��*�d�6�C�71C�9��jVv#ۻ,�������Ȫg%�t�>�� Q���WI�*FB��F$���J@dZm�8�K^r�4��%��o���I|KD��2�̯|������z���T�Ѵ*BJ�ѭ~������e[h�?7����d�bSP֗O�H2a��/���%��Hf�Uc��$���y*������u3脨Z�����p����z��Ed��AWŚ\����m?_����CV`��}AU�mfB��i��U3�7����rC�<)�aZ�`������qC��#r�_�؍�����z5s�AO�咅�w�z�)�0~����U�[�Ul��3dZ�Ԭ��p�z!'��0 N�S'�Bzp���LC���2��KDV�;�Rx���w*��by�!Ik2�K�A7�����2����k}{dDP�V�i�����V�M�޳��I�z?	�K�@���u�O�]׾J�6� ��9����d$��J���gp�Z���u�Y�+a�S\��������5�Y�et�eȟzL, ��;����q�ҏ��Ikb��rkw�)�"4�7=��/��V�9�8�{-D�@�:UX݋���"�	kmg�P"����}'-�����'��U����x���m��YW�-%C�����G���,'�b�0�椥�/�MF����N֠���$\�z5�NS��>=�_����)���Kw�y���A�8�P:!�,G���g��`NyLs���M����0,���,'�$�x�D��] lG�B�Vr���4'�[��
�r�QnXf�U�Al�O��c8J �H~N>z34
I�M�6ȿ��s�V����g�P6pF��ؒx0���Wr��s=����,�Zڍ��^U.�=��{��Ҟs�FU� �����X��BGh愱{�ĢP�Ku�:�
�m<o|D�d��?�՚ъ<|O�0��Mo1�ǿw�V��yk�l�ǂ�T�.D����A��*�&�
i�JA���[m�r���}��QCf]��9i)̇9�ΟY�`O����D��I��7~�c�U�DI��.i�p�<b�F'�� �tx��9�-D�U��,�5�1����#�h�:����6�g�+f&��@ ޏ�,���Sh�z�ë3�:����b" '�U���W'�Q�A7�	���$��f��-��%�#K�a_��oW�N�L�Qu]�N�46(�45�ôx���1db}�����fr�n﷭݉"�N�'��FF�{	bz����~]�C;��7�s����<%�_�o"o�n�_��ȝv��D�2�Y�� �) ^�C��j�?�e�<��r6kd	Pݽ55\i�A�	q��*,#�%�`�� F3�����V���T��jѓ���(e����4~/��#9���'����&3j����x�'4�yX^X�e��fuA�X��X 㢿����\�E/�,��9ҵlo3a�K��cv��Rˣ�t�yzy�P_y�����z*|��&k&�=Cwm/�bT���(�5�q�9���DZ�ks���i�nN��{?{��o���ʺ���.������aꈭB�O��/��Ґ>�`�����S�-�=���3TSl	� �܍G���i��aME��-t}�K��vl�wS���q�Hp|�����T%�:���6d���0���K��JA�B�?ҭ�k�]gҶ���:��pS���L?+���Ph�nl����u�H��t�cо��~�:ã��lլ��>��!]	|���V4���T��6�cKTҍ�1��(�.�ոW �����AI+�֓	ϝf��vd B��}�<�̭7\&�6e�����/�� � ��P�����f@�	�s�uJ4~�Ǔ�/$@ԡv@'��5��?�Q�Ϭ�d�?�Xњ���QTX̫��9���i&Mlz���� W�J�c��ǉ_�K��8ap,&�*�.���ثS���4��73�n��_����ROě\������ӳ�hmE�P,��X˝�
t">�Ay3'j�!P���(�$��lJet ��PP]f�	=U�8G�����	��J
j�G7�x�-kns�S���w�i�0娔j�@<b1/VA&��aKM�S������8��?�,OMJ6k�{�|A�%��.���@H�l�Q�ARɆ��a�nJ�o��\{FmŦ��j�Q�X��`'3�N>�R�'�-g�/���&��5��x]����N�π���OXW�/��ݮ|�"�m����Ie���) #�=r@�MUQ?Z�x&�����$���~/�%��!�U���1e,�XJxY;¼�O��ꐑM�Մ(����.�9���o2Ra^E��B
o�?���8�#,�|�c����c�< ���,�Bdl&Ҷ�#Bj� i)��C�����IP��$�Z��7nv�u��B�Hmj����!��Pt�9����b|����$"J�2�s�E��Y������ �
^�#j��F}@Q��ϊ�P�-�|�p��
fq���p �	َ��p��?�䆯�I]d����-m�0������էrs����V���d����G��j@�Vy�B�1�B�mN�Z�;��̕CD�gP��c��cʽ�T?I��_���^�%ni�t��f�7R^�R�+:A��><��؆���cb�}�����"З�����qy�S���'m��{�ơ�[�+Fn!^�3µ.7
��5����]%�QѸxĄ��� !�̣تq
s}}�(-����ٍ\�A�0e�A4��;���V�� �2G�T�V�Ɗ�N� ��`܄*�A�b�u@N����O*d_����{�bY��T.���'@.�Ηhfz��A�ޜ��Á|][GZ�di5��Y�!ŞZ	l�A�gy��� r��f�J.�������1lx��n�(�g���x��5�,D��6�N�5�Q?>:NMw�i��1/�F}�܊�w�'�W��3���hJ:h�G~���6�Lq�z>�(K2IPS���oN�ZBոނi;ͮZ.:�����^=����,�K�t��v� ��	�����\��2ܲb�����|�
^\D{T�<��ljݴB�e�s ������"�1*?�e�у� _���b�V�E��ϒ7�:G1�
,���B7k��������ss����ʉ7���ѴJ;�'�#k`�O�����KN������LߓWt���1;4W��/]#ӊ�l�d��U���Ռ��|s����أ��D ���z�`�!���e�~�D�\|�[c�3�<+�b�9	�p]p��Q�˛���w0Mui��3��>����K�b�������o����k�Pc����� ��t�qr�a��5�h�o��"]E���6�T��%����}����XLuL���o�zF�*e��A^�6�c�����	��U�^8u�M|�;�w�,
?�m�T���O�Aja�[ ��U~IE�m�k}��3��t0vM��(e�Q4��x]4�Ι !��	�>�cϤ�˄��G(DH���tY�����<;���[eeʠO-��ݴ�Ffy����4UE�u��;Nc0Q��oc�h<
D���d���z���;�$�4,�բl���ғ�aGq��sS��r*����ZvV�bƓ���b5+��y@�=#Q��G���m�01�+��>��Wvç�kZfYl�aL��/��B��{�t�1~��>G�u4p�<#BLIcE��||G>A@�\+i�Ŏ�3��4TyJ�|m��C}����*���A���D�@ҥH��e�$�N��b�dX튦���vt��YUL&�b~�$+����( �}�s�!k����w �.�7a+gGh��T��N�Zj�8����y���g3�	�z	=�6m5�	v���2��$�Z5�6�I�r J����@��`�<���%%'�J�����9��|�i+�!��7�<<��l�z��T6D�t��lpˤu���Pυ���[>JĘ��,��T���]�6�@3ޮ���$��G1�=L����y�zp��R񊆧����%�j,Y�m�g�Z��Y�#�v��$���Ô>��*�޻������<��J�N����h���:�Qx���,Z�h��8��ܕ2��.z��ա(�p�b`�<�K�fdk�dn0o`p~O9�E)�8�-!�~Q�Qz���4<�I�冸e��T�L�*��Z�/�#p���rFBgsK;a����xX0@�Mv�Kʘ�4��>�q$<m��a;[��y�"bn���3+��W)1nS��527�����������/�M �֣�zZ��������к~qa��<��_�^�ʗ�ۘ�x.fM�9]��m��� �@���jh��'N(J�-bW��PC�1�h���LI"jE�A/ok
0��u�L��X�tK��#��H��>��:�,U���3-����g�����8|���aU�=����4���R�]EY�Ŕ�1sa����+(���瓳�I��j���$3�jw���6�7�T�9����(�,��y)(k���'�:�Cm��&� Y4CM
�� ��~�f1��Q5���pJ����su%�~�	!��"�s1�~�]�t�m�oL�p�վC�p�����F�[(.�m��nXOJxse�?� ��!}����S�a5�$����b���G�j�!!D0�L�yP'��T\��m�_y��^�.�±}�{�wΘ����Qz(�uӄ��p�B;��w���2��v�
�%�-׵EE��TԢdG���ER���Ah�F��=?f�:U����N�#��t~"Yv���o��r�j����v�Z���_��-B�+���*��]�9���F8���\���6�'���HZ�q\�1���5�Hn�% ��8w�wA�.Zeމ���R ����/���A��EF�p����43��-�Հ�8��*&�N�%�_J��!�E]���a
�)=ExM�ە�.|���B҇�]��8��i��J:ط��q����1ɞ�UT�Sx.��Z��/^�G	���� =�v�[2��hbN�&loq��	پ&~��QI:����1➶`����W
R����d�H�s��.cl�%�V^��	��t��B68�2�.�'�����-B!v��a�Q��$,��R8��4�����!�i����^4AH�g��E-�`�H���ǀ�}n�g7��t���=ۖZ��g���t��GCӻ�g��~#�n��mme4~�z{�8��TVI&���q��1��O�����}&Z/��u��[�S��)�E_�&g�a3��dqE��+�T�5���qN�N���8�#�̾+�h�����]���p�^��M��KuMT�twG�=Ù�Q��)3�TCP��hbNeX#�Z��V���w�D�c�Q���O s�^�us��𺝽����q9I�Q��y!!�?,�:t� F�<�������h	b�$��5��0��$U��v���p����ڋ�P{�/�J!�b�!�'e5�����������k����D�M$�5��a����lm+��@ �Eѹ�i&c{M)�흆��������Pd؁����wh�Q�N?���ժ����� C����`G�Q=�uw���Q�}oе3D�������fL�d���;.mg7������i4���0V��Q���$<�+D'���๯�C�:���I�U��s�{�{�_���x����}oFR��)�_�}8�J�Ҿ�{u0N�2�5��^��8���.{��ŏPS�@�����ۦ���G1z��V[Jq(lC)�T��jZ�%���@�2�Q�o�aF�|?��tD�fƐ1TiF�ƚ��]s]�k�X}r���,Xj0Ox��(�Dc	\!8A5�·��}n*�zN��H=�Y���^R�O�2gɬό�Z�5(WU�9,�nz�0~]�w��I	s�t�u��h{۔��4�fJ��<DMhq���|S)����##i~�;~Yi�/�jj��i�˞g�|�w?��p�bC��]�,{��fX���+BK�Ř�Q:n�I�gZ{
֤�[�	�O��[�$�UO$��S�� �iP֎�!X���KWu��%\ڽ$oDh6ag�^~�֚�4����Ih��u}v�]�i��,mt�)�k�9Ad�yL[�u�b��H��&�1]���O:���E��Q��l �w�Ƶ�b�TK��1}s2�!�&�$/�����FxN�G��ے�i�&�8t >C�X�Ϯ����X��r�$�r"Ke�y�^�,'3>�/���ƌ�ң�}��.d�8�m�F�'�T�7'k���2�s�<2�7+%�}bf/�h���ߕ2֔ݥ%%/��Õ2�m=Þ���L�f5�c�A���;��yO�܄ �{Z�dЉ�"����<�	�uP:������c:_J�����ӳ�!�GK��";Nq�8��#"�j1k�L��d}�,�D��r�,�@NO��!�0+b�L��63 ���c�-S��%]�ܧ2N��G��5���\z��*c@�%��!q���X3�{�;h�j,+��1��|��LY~��F�8i��>ud(rΥ#�^���[孁�X=cu��흤�H�Bm�P3]	f�ϸǤ���z U[w��ގŦ[b8D���k)��`m	4W�e��)�ځ9�ڡ�;���#����B	1ǯ�=~��o�o$�z������;3.�e��^�4�_N?��q�Gv��Bp��O�v6�?w���'�n��l^�e�Dm�R�����ENdH�̀�o�t�Y*"���#Q!ap2jغ���8��ހ�c�=�4F?�{�)_bQ�9��L��i���}�Cҋ����l�;���n�0&�
�.���U�>uD�6�NYK1��ɂ�N�L�&�M��(y����oW�5N�`�7c+{�^�+�S�i�Ă�2�*�?�0ež�C!�/>J)��'����g���&>�X���;�ꑁ�:�w�}�@��~��,(��m尰�aS��	�:l��<����{7�X�T��D��Z~��2~§5&�*�!�L5�
kc�F8[���x�[Ǐ��L�$���{�(�_�����[��|�j�����!^�%ɷ �6�Gĺ��UWG�)_�:�A��m����SBx�f�c�o7�z����펝z�9�r` L�+yT�u
FR9��a���Z�]���VN��,
�RO�ePK�A�K2��8�!m�}�ȶj�w�إ�L3���[��@-�O�CN�P�qHm��c�>u�A�6kV���:�4^��K]���8^�,�W|p������#p��e�R28���R�g�]��>����#��M��>��EVCb�8'XR��Iz�ܕܦ�4��MBb�׬��>�v�ZL����.�s
TZ���O\Si�>�Ƚ��~��p=JxCM��ū�O�	�M������Q��	6�̰7��lo�j;���߅�n���ņ%=�/���w�(`�Oi%v��h�ڮ�1#��,>�h	^*>A����c��Q���e��g�G>	l���0��@2/ٽ�O,�6	��p'RhLP�{�@vD���M���Mp?O���{�)�N}M�񖆤��MS>��1��((�eB6S� =�κ
yE0k,�y �(E�ϸa+��ZU�$]�)s����rE��,?�?ryC�l-n�b��~�N�d!�/�u`BT����GD��b&�Y��v��t�d�����)�&�Vv2�r0�D�|�J��*���/�p�!�ޝ�Vu�S����#Hl��C����k�@��g��e����)x�|a�
���|��Zt�� �
V4���eU{O�t�f�%h)�R�D�/���)wJ��e?6�d�4��oS=n)R��##x�*,�KI�(@i�[��w��"F\�=�.�E��F��n�%W�:���qt��&���jJ��$��ϊ"A}��9�i��#0d�OR��3�9���d;�x�(�h��ģ=�|Zd��bi�L!D~p��D���y�;eh��xs| ���v�Z�>7s-���:�Eݭo�~�F���H34��v���L����?}x���>h6� ��m�����xc�ݣHۑ�{�3��?�)k&(2�*�;:7o���	'\�}}�;������X�s"j!7�j�3b��AڧF��4�v+ޘ<>�Q��)��f�Ăe�/�!��Wm�f���;m�G����/�W�� w+qx�ob
�e��:x&���=r7}1W[x�m�7�FB�k��F�4�Jļ�rS�C�J�t[� 5Y"=�̟����ݟQ�)̀�\� ���Ez�@��Z:��O߭��E	>в�y	Λ�yv�1�Ә;�2o�6Xs6 D�" ���sY��+\��#F@c�-��r9r4�8��>έ�]{����DC 80^��k,��5Y�xl��Re�q~�q����/�g�{h:�5�`�t͸����"rW�<~�X��i��O���)TH�O|��wLn#PSg�?h�&A���5�H*0]�N� _���A����\D�Q���d?n5�/��B���|,D�O"%� ���rl�a��.��M@��	"X�9��P��N�X�y�Ł�]�D��Y^ߗ7�z��`��Q;8Q�Uҁ�LJkC��r=����")�I����7�I�iH:s��sЛ�I�F0�#�9��#֎�Ԑ����Kc%���RK�S�]{u�֮`�ƥ���uWW��=j�?W�iVK�xm<Ka���@���9~�3m�n+����z-�o��8�JG@�3v�wr�5씪���Wv;��n�KKW�Y��XS�1<,��I��*_�A~m��2��� x�ʍ�[���<|�1�߉����<Oʹ
�D#t`{z�
È�{�x��;>����v�=��G�(����:'��5����?�)
]����ɔGZ�[Ñ���9PiH71&+��:l�:�;�xj����gB�D��n0Xs��yV����G���xtLk$ �XZ����U��fy��9������t�a0ǖ��s0�]?ɣc7��Z�Kᚫ0�ڮ�����z��0ӻk�Ny 2�f���xw�x�S7M$ ��ۃ],�?�+�\G-X9E^��P�򭝾�]���l��,_,N@����lt����P_'G2 RwRI���rV��G�h!�
\����/-�����q�A/���s�(׬Z"�\AG����w��h��4�n�nSn�Vo�Hfg_��c���M�$��> ��n&I���[<�4��4�������"��ϗ`3�~��� 8q��WJ�C��]	´t��}��������D��]K�'y�  F
)Cy�5q��CAR�K����ͷ�M���>!��-�G�g�q�i㰼�q�ٛ���D�z����1w.�(Z����?%<��&UPI��'U�Alo��rO�����,K�?=>z	�`OL�E�E��؞X ��'�2q��E�.M<�%+^���݋S��í�ս�>]2�:m�� 	�<���0��V��+��N+`Č摿C$�\Y6[�En
9��@��X�"\�"�3�
]�@�p˩�؎�Œ�n6���H�	�{����A|#\��E��ǃ(��o0b:����o���923�XlO��c����ͅ���K�(x��p�Q���ͷot �}�l�%J��&�bSnY�Y�L�Ol�R�]����P�I�1�T����hx��(��$��b��;+�]����F�b�^���"y ���w���:F�v�	���0�͒a0	�?�K���%a���^�L9׹��'⒰q��V����9�5G�d}�/z�߹��4�Ηk�.��۔�~��?!ƥ|�pR��8ǈ��i����\y�fsB!���2���=���"$7�K�*�㶖���q�
;hq:�����Yxq�����H}d�G�bJ赇%1�lӺ�iZ��R�n��:-vO�ix�.����\�h��G��-fVs`8���H'� ڸ���A���fp����mB\��`�L��v#��XV��:O �Sf)<��e��=����������zt�-���V���P��uk���-�T�Ц�p��q������=��c)�v���|R+�!b��c,W�a���឵������K���Z��PM���Qi$�=��"�i�o3��QbP�$�#�o���W�t����θu�2t�﷿^��퐖�4�3����n>�ͪ�u8+��^xW�`CgQ�i�r#�]�+�b_FJR�]�1/fՈ�Z�"��뱴z]A٤�er���\���y��T����1ڧ�c�>ȍp~߃R�������TN�ȡ������H�&d�>ݛ��V�7�%FE�6�_P���D�Ho��� �ֶ�����Q�R�J,�E)�T�cO$s9A$� �g�m֮0=#do�d>����G��;3�L��Xn�{�,E���
X/3�ݚ��u�T0h�Et�[�����aD
p�<wْ�p$�_i�7EVS	V�K�Ԑ<��Ye��w<}�[�����03ڃ ���ָ�
��*�a�̉Y��ѓ�b	�2q����b� ������� �z��J�7��/���qu�&[]�	d�_�USp�!�gIYd-ja�=���v�*��H/��E�"��9�9�-c�$djn\YN]h~H.�t��*Ʊx�)P�7�^^;���`��%
��`��fy�L����eZP�����2�6p���XY�!��1<�>�ik�V��˨����X��uF):QS-�ԁ��=:R�E/��M(��G`8� }���u�NaO_��JY�e�;��A��`�S6*�ʇ�-�C����:�ߗ�q��v;U�\n�;Ҋr�[Tc��at;Ȏ�9�����z���R
����*��g�b��x��F�G^�.B=��cȤ#�nMN��B���a�:�%�|�q@k����y��uQKr��l�%�z�ke'l��*�ï'����"��9UG�"��Ѣ�X�?����S�(�-��Uz�n��D�(��}_�͏��oK�/��Ve3�K&�v�.�:�M�_f@bH�)��q��6l�'�R���g�����߱��?�1i����T��Z��I{��'3�N/��o;�^޳&z8�������c�(���ͺ�,��MXϬUe����aWa�T�2�������̎� �m���E�^�����15x_�R�ܗˣ!��֊��Sh�D	r�{��A_�`�}�=)�O��wk�s�9o����ώ��Z���u��̓����Zb�Q�7�MBph`%���Y�k\<K3�Y���Wv�H]�q�H�����GO'~��f���/�_��h/H.hp���~>a��f�E�A�8�X%�Q����(�}�wf��鿤�..Ld��2�,�2Ŕ�o r��m��4#0̅��IM������b�Y���@�.���޿�{�W�d���8v�V�J��6o�>@�-^x�cҦ5i��?t�r��V_BO�Y�rQ��f��أ��2��ٷm����=�Ʒ��d���XvE������a ��.]{�'_�`�]�ʼ�$��,ȔI�`�k���g!��O���Ð@�Z�TpLڇFt��X��#g�BG4y��G:l�I�,}�L�zhR9yE�֥>�v_IgV+��]�Nf��ndo1�tL+C�n#�KbCwPe���Tq��������J��,	c\�V ?g3$���jka��EqS�p{Kԡ��NO2���� (����m(����K�uZB�����s����v��7�۝��p�Ž��0��G\$(}���)^l��o�[��odT�c&!�T�ߕ�����a�,"E,��uU��;��\��,��*�uG���U|0��g�-ОY�<��(�#ٷ��h˽ǭ�	Ir�ʟ�t�1F���f�m`K )����
����;\4;�ϙ9���x���"$YY_���!)�ݻ���#6�*`��T$-b���_B�֔������90 �c�,��M���Ơ���`D�p�zˢ�ʷYb\Js�#�
�_ż���W�A��F��Ɨo�ݵh���K�'�'P�ʫ��I�8.xl��$Rܞ�_=���~kx4����l-��/���(�e��ǞN���R_�qU�Y�wS'�e-�'�,ty�Or���,���G��?S�ƃ<P*J�I�s�eB�2�ܲt���սk��ei�v�L[)���C<晱���0�V�<��V��?��]p�Bp�Y�Y_'�ڔ��8,|���:~J�I�u������Bt��9<�)�]r���	�($��A�2����EǬI,��=�&��4{���߰?4'Un��|�b��n'oѐ�~*�����v4�PW4^�<d�i�:8�\;%�@�Ǥ�������r.w/��� 3��`5�P̶�n|:�֌�����S���9Z���`�8�*��^�aa���X=��jS��k�����;1��T�_n8�r��5F��b�
ڇ����!%?ô[u����7h q?���Bڈ�ǜ���oE��]��Y�n�,��H�M/R>�^Λm/�<�<�?����h��A} �Xtz���ڱ��m�0v�.�Wᮧ(3�ڛ4��_�`�OZ���y�5����?���K,�tO= -�@����D/Vq !s�Zm��Ci��7�����5?2+����KF���oݎ7vJ���p�v���U���<y
�
�U��(k�T��O���֬ĜpaA��Z�HU"x`x�K�Is�P���bٹ_��<����;�A@б�@$ڒl�{i���5��b�/gü~�8�z��'���|ʹ�&R�S�f�d���O�ӣFR�����j̬�ŝ l\m\��z!kG�����&�?�����͋]��إR���O�p�f��6�����ۧ<�����s1驁޴t�J�@7- b�\�w�[tm�6�>TF����`u�3���.�b���`RT&m��zL��s�5,��s��l��\g�I`[�<����{����?6�����۶���.�N����q_@uu1��TH�n�e	��L������J1	�)�e��cw�:T�o�Q�3�1{9W0>lQ�r��|�C-4��EG@��3/�Fm
���5h�(*�U�9��8�>ju0��h��)�����ɜ��e(�b��˖g���E������>ǀX�".�"
��UjD��N?k�G��LElk��(��O���M?������*�T��Sor"A�7l�"����%p�wfS'����O��i��|�
������-am��ym��<�����Pg1�%{�PӐۤ��!�
�b�L�`��N�ߨ�ԧ#;T/��x�b�+z��g�$|o+t��BE�U����?��}�Fڮ^@5z47H O��[�$ ]�Ž��X���P��,W#���O�j�������b�T��F�Iؾ��Y'�
:�!c(���.|��U�~��y��JY�(UV���y���Ut�������/�.�ԃ2l���.�����x.f!�kj�HTTeDg%�k*H���i����j�����&����+�~tt��EIm,���6R/y�R�����L��*�7W���M���$��Ue�����g�S"�1W������X���~\l[9�>B���\ywr�r��TT�0H����<7�YS���ޕ%W�T�jpݥ��:&=��>W���elp���`�.����"~�j9�[���j�HW3���f����O��q�PL�~�V4�+�?���y͂��6��HC5t����o�{����������x����ߕ��*>K�wc'g�e��wV������e �7@����)6�����4�������? Զ�\��gn�J�6�뼷��z-��CS��Aߞw���^oR�Bқ��P�[�����<����r��)�ᑚ?J��S�`% �"��!=� ����"�� �3��Hd�ꣵo�FkB|��67Y{?$�i�/�p*���M�� ��q��=�[���q�l3�/	y0I+�o�t�L��͡=�'�U��/�9��{��kh�'�*	��\��{ �]�oJgS��������M]s~%-  D7�Fc�R���(��Z��F��25��6���0Ɔ�D���Բ��=N��T��ZiϾ���)���#,��A�ּ�;}	����lD��/.]J�Nq���J���ށ���#y=����.[V�
,"�V�Z��x ��n���9FhM�e�����6 �(v�k�vRs��|
�)�,�f���Q��N�˫2����8w�j�mG�yx�^�2���@V4��#W�����9�TQ����:�	��h���M���� p�!&��S��0owz��ǅ��,qrpu�?9I"������Ih���]���PgB�>>F�+���W�����%̬�[N���9Kw@����A>��b�"3��Ǟ�m�jJ����-��VZ�ؖ5e�ըB$�!�k���̢��K��,zj�ez �'�nщ� �Dܘ�&�.������ȕ3�$dꜝAX��_�Qg3ZE�<R�p/<©�W+�3�b��L)�\"�*���N�1�?͒?R#�CA�����:�,58�đ�We��2�%���3����Z�^��Uz���u�C�!	L�����ul��7�Ep1�0rs���"�ʝ�������P��"��u�TN��X��)�މ��T�����$@c�:�?�-VKʱ��$����g���XQu�W�F�t�=�}K`��nP,P~�:����(庣�s���a�Љ���Mè,�p��|y����!��7�'pm�����]'H���Ӂ�2��sς�PAN<��q�»�Jb�QP�k-`�n*��L��'=�I�PV�lG�o�Ka�x��e ���B*u�u�*�Ð'�����$��+���^ʊ9�/[ҫ�t�hC˃Z�@�����:��Q�>UBU�0�z./~�;����x��� ���bw7\�zD!��P�-f�j�T��*����a(Z!������.�h� s��=ˑh"��w�i��x`�G;�mu��~��h�g��Mf&�e�aHT�/�J��O�����}��KSb�p���fjb՝T��y�D=>�����(�| T�/
�g�.�ś���l�eH�k��R�}��%�3��<?�WN�{m!���<��}u8VY��tst�ض+Xfu��)�BQ�����5�^k}+%k������HQqA�\�X�"��Z+@�"U���B��rX G
�j|�`�����mL\�(Gr5������W�����������Ǥ��6d�vڀ��ݖ2"/�i֒멾��Z�d#٥��2�!��>�ݸ�M��f��K.�J��=hȽdIBL�ڿʵܣ��C[a�m�b��aj��OG�S�[Z�_�3���/���:�r�]0��.YI}�Xf��܏�T��O�@�&tj��-^j��bܰ�u�)�9��!�sL��d��p�����?��h!�;4��hOP�/�w\�J�w�6�	���ȧXf�WQ�����<�)���jt8�գdΡ�NG�sf���i:�i�������2s).�#��3��E���N�� f�1�WWpyr�����] ����gVtSmgS�|";a.,CL�宍D+m,�C�P�������x�Xd�
��Z�^�q�ϻJ���E`��v�o񛹿���WJc�w	a8�}[�\5S�ig���Doˌ��~țSb�1j��]���;ܹ�;�8�IɽØ?�ã�×)��R�IШh .��*�����c����#�fW`Jw麮������N�#�h(1�,~����(��̀t�i�UHW�;� ���9 ��؅MCruto8��=�����vN��l��	�p�Ǟ܈<ֳ�b$�8j
h�G�8r:����$A���;Ճ6���,G�PbY(L.��%�� �nU�^��a�p��om�+��]��������K�@�h��ϲ
( �n#�sh}T])+���U6�,	�
�rE4){��B�: ��w�qg$Ւ�C��%��q���1������!Eu���o�r�D�	7,��)6Xί��٬��6+%�M˅8� �q!3Ia�
T�����3 �����|����T1O@�Y�Ӛ�1+�(���$�rN��-����Ꜿ�`n���RB�ҒF�������1[�|�W����,6i�ʐw�݂J����L�Za�7������UV`a�����1GW=�V��Q�N��,R�O�u{�'j<42x��@�`��h��[��rI����>p�*(1M��k�K�b	��V��~�1���q |t����?��P��t:?x�8b2��iƲ���0�ip�W������=��3=����U4Cia�\�����y��ܚʳ;�I�"�z��\� ,�M���f������^m-�jp��h1_z��jID��>S,��� ����<�vm�Q�G?P��X�ʂ�ڔl�����j0���u(��˵J�������L!7y���~A�}��Cs#9'Q�x7�S����[��</waZ�4���MP������g���Ij�G;�1O��(^�T-����3�_K=Zg���҆����F�b�1��)�uX܀��\��F��7-�o6(��ғ12�?���4��c�<�]q�fAE��A3Խ�4=Z�^����u�9}��1���" �U��f�d�@Ս&����&r1^ztX8Pw��}�V�aI���/a.�uYp�^�_|`n�8՗����cEKd�p�N�����#�]�+C����S��c����1���t�D�J+�*V��p��#�?W��gk�*0z����'c��=2�d�]G���wz(��'q���S���0�M�v�n��8%���~�9v����p�%��cOl�7������qE噹 �[����~��)��H��� �pvVk��O���5q��N��a�;w��6�?���9ʔ�""�~%���}�":z�l�$E_�h���2���+�\���l0�U_B�W �!
�� 0�K9p.�s� V	B/�Ş6��=�y$P�ӑ�ֱ0�GT����o�]$I���3�Cc��[O�+�8�\N�'[h Gƣ_a˸gs��E�~���J�$ے�x���f�*�WY'�r��?Z>:�] ��=�������Z>ȢS+��~v�
���ii�lD�wC��SiQ|rD��&���;��E�Sn�5�뜁
'e!vGgt6�L�:iT[�έ�n)Ȋ|k�w�'p|���N\�Y�Eh��7d�p��"�	[����`�������@XO�y2pO��3f��	E�s6P!A�F�_5��w���A`z�V-���^>���\4�m4+
	rP�}���&��8���>�H�#(~��,:"t��:���҂��Se}�)��Ĝouh�mØ�k3�y�jN����-��
��L�?z�.��'P�R�e���Ϡd�-Ļ��{b��Mf�}�Z�9�>ۭ�E�G,�Km�	�2��H&hJ��WJEK7�1}�[O���/���gb�@�e "G��;U�ds�z�us�u���m����֘�#�X�2���vl�3��|�-�b4q�C�yb�N��:���?S�ڋPNO��}j&��S:Km��=�A4k<v��� �8}w,	�s[����,E\t�͙IA��C����`oQ���[��=*�u��Ɛ9�Z��xR#K�|�`�Q����� i�7�[�a���BUXf�XM7����@�rw`�1����Cw_+�3���V[��� i��h]:��:P�tR;)\BE�j!��Ds/b��W�G/��'�Ζ5G��4wD����i�S��X�Y~q��J5o�@;��<���z��躄a���'����#�&^x�F�腒X���[r�Ƶ���j��_�P4���K�$z�>>�y�uQs�����L�k9UZ��Y��v2�.+�W��T�G�[ʢ
�t0��|6x�j깼
͖ӌ?�"���T���ʹ�z ��Ve��V�?c�(�?��E�B��yJ�8�� ��~A3~��Z�F��X��D:�Uu1� �P[ZZ-��XXڝ���1�k�9�l#��JJ���̿[���YN�s6$�Q2���Q�tfd7�>\�5�j����>��k3v�wZ}���Nm�52����P�9����[�Z��s�%u���`�q+x��(�J�[�l�(��	�{�D��s.��S������u�,�j{��<o�fq�e6a��PkC�r*H��[��",����XǍ�+��03(�;ͣr?�r��	�K�o�LS�w�w
Ø[��jP�U��ἴA��; �Y�����gGzIH#4KP����8�S�2�������6ZP���.%�qW�d�X$s�r{}��=*]����	�&�;l���(��6h�jH�cl���tb�O� n���r���Qc�p+'^��0c$X�S�
��.h~�2c������1x7/�t�'�0h��cOx��Pi�5Z�q�O��,�V眍E溅�T ��}�[�~�)T"�𱌀��8���X�]Dh��ww
���,�KP>~�%�3����b�e'��6�tl0ceV�}�e�n��!�7������ X
�]57~��5�ل�|Iw՟�ϧ��?���%yoz��~,K�Jx�S{�9	�@ͳs���NZ���ۂ��g���]�������xة-T�I����>�'������Y���f^��^��zdD�7躺�{_X�⛚����~f��]>M�y����� �Ɋ2��7����	R%�:��H˟��s�T�j]D�W�\(X	���Y�	�>X�2�bA^�Ѓ�ׁn+�d�S�����x
�sQ��!�N��=D)I���n#|�1F�{%�p�86kﲺ���LXg�R	Yݏ���I/9	�#j� D�$3�z[��	��PO�q��K�UͧL�&V� ��FT�&��U��vk-`�����2�Z+^o�g_L����L$�	 �q���B������U8�Hޮ7��*�=��U���M]t�-J$�5\7[���hi��qC�3Soǌ�N��/s�fF�b�M�#'��y���.Y����&�铁ƽVUr��W'�j��2sAe�3U.h�L�T�L�0F �RR�0��?��ڽ�����.Z�bdd�Aa���3rI����6wA�?���&)�����1�;*��d<�&�9�>8Bh[ȷkgO�Xb �OF)��� ��Zb��Q���S��4�D��a`?���+?��EG�fnu�0P��M]� �~�5��,�ewIt'��:���M)OA;S��Fa���A	�gӒG�'s#�R���A��NL�u6���(��փ�h��N����5�|�y����oR#O(͜L0���l-�Xwg�#^�׻X�H�; �-��IO��R����'��
h}��wpF�hn�����϶���c�����E�:��d��޼�y'��@��c;�eؘ�gL'Fc���A��a��\���|q�U�Ӫ4�ζ�Ob1o���*�uX�y���Q.����|��˜�"�X�
Uz���.�`W*$%��2������{j>�1�����I���R|�d�8O��x�Ĵ�}̣�^$|�Hz�B^8~�.b�'V��
���b�E+�!���g���rsT�ޙAuS�ӄ��Sk��?�?�Uvo��7��!8!yb��v@�s�!h]��1�܊��v�ZwT�>0
��9T�Y�ʆv�U�4%����[�NltB%B$'9 ����;��.3�I��:��Y��`_!]u63�D��֋��ଆ��i*����F����0r7�:#���{ӆ?U8�0ƑɻƵ������f��-N}fM���t65���qR���d�#�V�i��Eo܉�rvp�<�����4�)����E��l9ׇ��4������g}W����]�����_6M�e~GP������a0��3��+��<(}��`�k�eLq�E#L��&��x̐�Ʈ���ɭF~[���uΫ��Z��;7��s�I�՜�
��V��d&E,�~835��W�?�x5����b�p�j���v/�ɂ�&�J�_�7E���k&6���ػmF�⚚�X�̏�@VX0��=�n�:��z]�v!`a��b���J����x��mԗ�@�Ĝ�`�7C�2#N���KJa���{8�i�h��!&4��`�p#&:ydY�"�MJ^ !�& d�O�+�F� �	d��+�� *+���
�/k ��O>��ߡ���_�Ҙ�Rȇ���;��%R�8�&|C�`�Q8I���"q�f�;犸cRX��<}H)8>e(�rW�9:�sL����[��ā�%>IT�
��}�Hrڇ`�z��*�f��/��_b��O��ž���Wi��u�}	R����W��O&���"�Q�^� Z���u��s/I��@������\ę97�w8�f�dG)�Ma\�*Ԅ�<���l Lء*�H�L�tc���(�{���U'x�ǴP!���ع�x������S\��#�*a�],!�'��ZSvB�������C)/�������IT��[�oY7�N�9��EA�$(��9%3�.��$6��ѭ��]>	o�eO���rGDzI��ua[��}~�Ig�	��P�Q���|��p(0T��u�'�'�ػK|CW�nDsQ<9=닾�n8pW؜�0yyH�$�M��~�?H���Rr�N~c��;���5�T��3����\�Tdȕ��ϳ�`��d����HybG��b��ǰ v���上�]8Ӧa��!Q�].+A����2���#H��un]j��B�������#"4�T��VM$��y�|�)�ǣ:��A�7O����V�?/�")Xſ�5����H�<��; ��)!�|�^�.?���U��]�ɽ`�G9�W�lt�#�v K6����F`hU��*å����5"����q��@|!�{����G�ܔ|��E(§��?��nl����9 ��B�ݳ4�1��c��Ue���[��բ����^��<�O�)Y��\�e�Q;U��D�~A��!��1`�ݴ�FӐs�Ю<�� 6��ΐ_^�M�s�z�<�_!�ڋ��=>�_d�y�ZKB�y�"�:��� ��:�t
7��`��ޮ��`�,�3y��k?����t˝ҹS��{3�� ��͞R�OY���8�T���Y�{v��<	���4)�A��p�����M:��I�= ���fJ.��
2F"��c�����̀S�!�)Q�sZӓ�и� ��'A 3s���2�Wq9�{�kq�mQ����.�xQ�x�G�L�-��|��	%�I	
2&tm����V�����X���;YZ���rP�^�ϡa�|���A�b���E�z-z4�z�iL��%w]F�;��!����]�K�n,D� ���)-�{�����5�{	�C,q��p���`ܬ�F�v_��=�@џ������/,�w>���u'c��҂�.c����D���h�t��w�~:��Ϋv1d����kM�H�p����J���`o�51�^�Z��r+*Y��ycTg �� ����/�0dne�\�Ϣ��&y�a.�붚C�����FTE����:��ٔ�\:)+�w#�Ō
&��q^k�w�*�|���/8)��
�XoO�ǽ-��˰�|�%�Ҁ8�y�T��&���~��v�ͳ�$��::�;c�zW>����3h��US#-��/v��,jD�tF��#�������� xs= `xbp"�g9�j�s �$�)� �,�x}V(ʇd�PI��q��u�x($��bX�a.�=VKC^���ᎋA��%7,�6��-V3�r�J�
�l}���T9s�Ig.�yE/�,�1�Zx;AvEO�{��%ۈ)��� ��E�D�!�4��3M������6MP���	��7��V+���Tr�hN�F����)���?Հ[C��*�E?��G�]Uܨ���t�DhF��#�*�["�8L�D�*�R�J��l���_��c7�D�;2�ǝ����!�������Q������.1z��,��}���8�f�ƛ�DC	)��r���\1��4��P��{�۔�����÷x�Y��rz
g��j|�u�����auȘ��͐��BM0�*�����@ՙ�����e��0�-��pLp4�a��s��U܄�3�ܡΆ".sF���R�ߦ�z��%��;ݛ����	�%��w7oJ~�˓�EZ&(c��g�\iN� ���t8�y��]Q Ǌ�SwO�E�4�L([�������u�_U|���t.�-}pٯ��.gu����"<'���T/Z}�z
Aq���z��XH{���5W���Bm����8V��I�K��;��B����3�*�V�9��B;���O!��=��Jw� Fz�2D�ۡ �y��Z�3g�8�rn�ޮ_���>�@�Ilv�ݽiJm1&E1B�ZlUTZ�&��%�Eo
eZ[��ą���(���-ߤ�X�����v{S��o=�l���c0W�y�@"]LĤp��d�$ӊ{�蔐	(�pD�M���� "=�/S��H�F�H��j�s�S��l�Z<{+�ES��&2/�(��.k/Q���z�oc�d�{�X�u*h(�Ӕ��
t]�v�A�(���?'1 �M��̤�_,q�=�$\O������oq���M�#+��p<�Py���)bR�T�2Y�����9��F�50��U�0��i8B;�5�̌^b 3��lr~�C����r��A��ұ���V�q>���@��֏����<x�&��6��ɓ,k,�V���{���}���3�:f@��pm�nM7&���� ����<�(GDL-3�G�eYđ*Y�P�h��0wV@I$A�Qf�v�)�Q!�N ��tn�*�Ʌ�Z���o�����W�*����(�##�L6������vOr��=cU�<q�<]���>뛢���V��'��*xکKl�$^vmM��ћ��Q�S�>ʐh�n�4�E;a�_��<!�����<��$ _wY��O���Vs��VI��.����O�\��9�h���q}R2�A��ح=y<C)��S���x��q�`\ҍ�����[��5o����y+�S�.������1fj�>�`bnH��F�;A�B`Me���!�T�m���F�W���L���:@�u�8�8_�������/�}S�����j<�SX��?�AQ����Z8��Ia�<��j��7���ɭO�T�\�7�Ԯ�Q�9�}liQ�n���_1Ho%�)ݟdO/GsV
V'#J���j�[<���־�9Rq�)�M�!D�|�1�|b���H\;���D�Ӝ+>�J׃M��(NK��v����1��+��Q��Ň�9!��oگ����� d*/b�\�RXU�O����f�/J�7\o���N&�c�lo;Kɍ%��U	��}A�3�t�ɂy3a7޴J��6	�C]��8>A� �H	��ge��T[V˨��}��I����&��5�1�HN���!G}�S�E�(���P6hM��«�*w��S�����J6Qg������Y�������i���ԑH_>�w���(5|"@�ހ�7j�ıXP��R�2��� ���#���� TX-t��g��|�Ztؤ�d$��4�3 ��~�)���S=A\���K���M�_Y�MR.�QG���Y�K��ރ��P-�~���P!o�"� G=U�oߒC �M�+�~��t�j��"d��+3�,86��_��8����K5i۹�
Q۰�������tX9�᫵ܕ�����bP�.����9�᳣il:��l½G�mp�9k�@1{Щ$����.��L
Wn��͐���?�OO����	��cGΗ���w�!L� �[���>�;f|�4�/��Mf�������x�埮F��X$]��#�]����VU�t�ҥ�6�AP	�yR��7kE>�%>&�� ���q����Rt.2&,k�3qt<��t�bԆ����a���&����^fK�؇�zI'��������,;����Ԯ��<ʛrL�j����Q�w�i�۝��͖n;"�	���F{�~L'U�0�}��(�^O��;���-�a��W"	@ʤ�#hG�֨Z_5Ör��j�AUWv���i39�_��*rAD��X���X�= ��V�֖N����=c��=x��c*�{�4�(.����-+��ӹ^~,���i'��v
-ʫ�y)���X�F҂���e3���0�'����Y��B��Z&8���[�a�ф�� $�MI���,�@�H�&;�(��0�N�F�=~i	�]�X��+�L>���y+��K�?������&�s��\:�U�Kbk��������!��ڮ�	O���H��k�"D�H�,q�@��h?W�-��A���m�N�#Иc�f}9�ή��:���6��g�ι:?�V�hF��,nN��)����ze��}臍|�/�3���3��4V=?�>���S$���M�rѶ�܄��}����,�
P��*�S��x9$��g'���ֲ&�����0< ��~08פ}�R���etj:�F(7�
�����f�=\fś���j�S�;�M���[?H@"bX6v�T���p�&ס��K�FJ�&:�k���xi�����įi������^^"��+h����d���Lę+�n��)��"1����Q��9[�DP�}k�Y�-h���v�5��½����̇r<��$'S��tK�S��[�;�	��ěg
����H��s$O3/�C��Z��e���oQ��<Rп�	�9�p�c���܂Hh#�#��в�<]����M;�
hP�~o5;�6�c�rp���qX�4�(Ε��O�~���}��Ø'Z0*P�/A-�`d�!�$OH�������@��W�8,\�t*7T�}��4�Q���N-�q�e����BN�����/~ �k��"H �wg����mJ��j�P.$r<�b��=���]���wV����C���έb'1BS��U)�	���kj���p����]L�O�?$U��5���([QĲF��5T��r/����Bǆ���O������ߪA\1�`$���Uk�ň�o.Ov���cǕ�K��Q���͆5�zL$|%�_��9f��A�Τ콈Y�Et(߫�����?|u!G���G�� �G��qg��eBH].�������p����>�����Q��wr�$K���"nd�Vq����
����{Q���3 3X0�n��"���a�u�E�;��Ԛ{=x��x�Z��C�E���!�A��;M��Q�S�3���R, �C�Ԇ��@��ηILʾh�5k1N_����|T���s@I�[�@�ȡU>V![x�[�~��s��T��*H`���q����U�}��/�"��5��}�	^>�]A��C���I��iZ��:�a���U��L'�(M"s]ۘ���^@��u[��a$�{�hw�.Iv�(�3�b���I�Y��:#:�	f"��7�W�z9�5�|{�U���6Q��\P�P�^/*��s�L\Y*l� ʜ�+��]i��g�f���0�֊���g��XТ� ��z��x4]��Y�ݶ � r�ʘ�l��Z&������R�s���f���
��bwr����>�J4]vӫ��q9i'�K�����3��;���*�
����(O�ʝ7�,�^C�3�S����X+I:�,G�S���:�&�m�D�e��r��}u�6������៱�h��P��V�?ǑַQr��Huɸj-�1�P*މ;"w�״�gx��1�x�!��X
�r���nZ�3��sV~b�w������`����R0v��b��r��u��\�fuE;��pآ U�>y\e����ı��%�<-ɔ֙(��mG�8��U����0fh�j�o$ު�Oݾ ��tX��\	�	!�a��4܎0h&��q����_���D��]B������AGn8��[hT��迷:�бB�<^tl�v����PumZ���@x2���L��p��m�[��Փ�}�A?�ɃZ0�:_V^,÷�4;��c3���,W=�}ޒaY��fy��,�ƌV(�U��dLOfd�3���C���H]:v��5�S��6��Q~~�3�d	�c���,I"�Ȇ�0��+)	���R�2$�',�Xn���1�(<m�Wjc�	jRX�c��M��,�گxS�3d�����4�^�����>��L@yb@�c�C�}�o�y�t-�7�qk�b��b3���ɽ���/8��^�� ?�_��qRp��qU1�;S^���R�#2�t_3�"�T�I�J)��J�7��v'�x�+�Et����G�e�8%�[� �Gh.D�J�Q!�!������Z�J �>`B9�e�Ͻ�H96��X�	�{� �!/Ho�f<*~��,K�M��(˒	?�0��1�¼�}��.���랙0�#(g�6�=S�O�x���C�}�8���b>�� 4�2���w馮U}@�e� )�C���p'�ti����w�2?O�z�&�1�޴���M@g�Tְ�y�4��5��)�N:3�m;�d�5�5hJ	8~-`��Ɔ[iC]HlQ�B`�C R�M^��M&���]�=�:�C�«�uK�G�?���z�gJ`�륙�3 �C� �/�-�&L�la#�:&����ޮ�[M�~!jy�Z�sÄڎ��̌��g���^'D��J�����²E廳�r�O�޺0v���<�Ó��~	 �|���&	�ə��F��ld��~���j��b צx�@ �O����� #�I��E�<��K�7	5q��b(��4	�ӪY��Pu��#�E8Vc��C&���1�t �K��Ά�G����⑹��I~&I��\��=L�:���P�N?aSe�C�a͟�W��eU��>���Ī
ZU���fR�4,GDD%'��&жz?������oyƟ&�ȾͰ�+,����V���(1�r�_otH�2�P����S��"2O�)��(�З��J�!���䁺$�c!om�燡)�:��{`��С�2o�'3E7�Y�E�!�$*w��t����?Ș�m^�׺*�v�W�U�.�b4,C�����o�J`|5�P��]������Kl5o��,�~)q���6�5`��˫V�q���5SsVF�C#�4�t05��p�!��:|{�vh�����{��O[z�mi[�xw�G0/�<�Ҫ�O��9��YR�'�d��W��-!u��B�+������b��S�.7��i�v+��j�/���uN$���x>yI'��F>�d��"}��~�>�����4s]E��[���0���Du�u�E����m�Nq<�Z�v����q�U��xޢ;�~�M�Xp�U���Q22(��eבՅ3K�}�}o`#���?_���y�DvO�uz|������?66��O�N;n֬s>��v3 <�KHqI��zE�GG�elp���؋K�/w�M���.�ԧ�8ڻi�+}����>����ki�����e����!�MK�j]��=Nx��vh�
L>b?m}�N&�A��9g���#'�*�+�bM�Ѽ5��Mt=��<�U�`BM����1�����Fw��ۅu��2��������`��X{q~��\Vq1���臌�����&EƇ����!���匶z6"����Vދ�e�e6����s�QJ��C�CF����'�>����撰ޏMy��@K B�5�x~�2�D�����*���J�k����&�������$��u!rn�-�����WT}yW���#�R�|�Z���3"=� I���1�k"y���������/Mh�
��_��d�x'g �&����n���`6(��B;I���gp�iV�P�q◦�Xk�}e�}�S��sI�)D�0]� ����+=na��i9��p�~���_��HuB�%I�I�:����΂a���@]�b���u����<�z�	�t���l�2��jF�~7_C�Υ�6�5dz����@'�>��N�᰻�d3���%Y���F~��5����ȸ��h��h�;�y�_�;���
를�A_��C�_����KX�|�_г/J��"J�a��� e��D��]��P@��wdH������F����Ji��xh��`��\��ۡg�i7
l��)/J ivӒ�#C�ns��m�&���
�ᮮÛ�KC��C�1��fⴏ�=]�2��C���q�|�)]�u��f��"��#LTX�+����X�>�T�yo�"F��1�l;1`Ζ����~-�Lg���`Q�/p���'�.�-��|Eط��+'hwT3
�F�&kJ��e���w?h�p)�S���줏����a�z���A0#��L��0="Y[�(��tt1�W�X�6<߀D]�y�	
��U��[�@8�cI� �O����v�Ͷ��q���PӆJ�v�8^L�R������;�y�_���:��OB�7�h�]1ngV��&rAo��'������[K$#�>�z	cj��<1��nw�?�:��q���� �E�x�s��d���ESe��ev��O�Jg�-�I�Y��`kuf/�X�ܩ/�ߏx���V��!J�Y9�Jp[z�[��y짻��L!��cو~�8�_�l(�4[�)���5��2J�ՊR ErR��ޠ��h�k�9#Ӵ��=�"b�������̙� ^u�����M�K��xf	-���U�(�����P>" �]+�<�Z����+�g/�!�ʨ��@�k�Sd�`� ��s8��13�83p�/ ��� �/��4ˬ��B+tJ��bָ!1b���(_��%��/�[g��r�p��r8�׃8E�'���빯���{.��'�'F���䃀O��w
�=��9P-�����J�޹p��6��Uak'�C��'Y�h/d6B��=�SPBR�=�#(�-�we�sfTE:�s���k�6�3�(��H��(d�ĩ��a��˄�@@:�V}w]z����Y��M�$��;DU���|�N��eÇD&�A�o3S2�ⰰCP)��S��<�5���g����aX"O�����eK��C���n�{5�ɐ]܈�kr����ܬ�~���hfQܗH�����m��$���Kޙ����rw��l%Лw�~�p"6�f�l�.4%,�B����h�U;ʡ�J��L$���[a�~m�����x��O>��"�0�J<P[͒ۛL���j𐟰{5脲8�ҋ��i�)�ମ��*��M�����d�,�Z��Q�Ж�yM#f"��G���;ϰLmQ`cYxx��iz�d!I<���sSN�ێN�̖)t�A���'p�0OӀ�?��F�)Z��\�[[��� �np�g��mZ�(1�9�������f_T"�p�C��r��g�Dh��h�)x���2u��˗l|LI'�|������i�W��d�`�W�P	�i�V^�wg�F��m{��!M&�=6(� ����^&�+7�:ϑ��[��
�/�J&?�����;_�xq�	n�b5�Y�W�A�N��=ah���_�8�		����:SQ,ʤ�u�[�I�|%H�l'̶icVE��;k���.f��xtl�P~��O�������a�)���01�@_5PZR��
�1M���#�q�'
z0l��wз�!��c���Y�D��w�Ο�T�^�9�n��WHD�,%�:��d,��`Z��J�9Z��r��ܢ<��d���j�B.$:���:�A|zyO�F��Ǥ"QY����C��@%5���e�$�+2T4�7���ukWc%��\=?Փ��\�Թ23D�T��[p޲�[�Z���{T����M������&�Gv�
�f$t�#�f�(�����Cy҈	k�^�o� 9dԪo��&8$o���Q�'�m��J��֫���,e2�������	�M����I5���J��+{z��l	�R�ua	�Ĥrt��:E�L@�R�N�Ohy'�KWW�ʔ�C�Jnvp\čऴ�؄_{�V>x�{�9�
�m$�f�: b&ZV��l����b��f��.K�]��:n.�_j|JW?P�(2��/>�K�19s��vQ][͇
�z�-'�L$Ý5i����dZ$x�(ZiV�Wx՚�+�O�.���w`�ܪ��2�3��Z��tbz4�h//��1e9e�p-�0�e�4�����Zݰ��Ô�I�V�S��rs��5�����2Sꢛ1��V}�e�$�B2`�OԈ�J��I�B\=z��!��&�E02��=I���H\ ۈ�B�.�yI�qhoʶ�iѸ	Kһ�#���`�#�� Q�7�Xk�-��ä��)j��$�W�&L��/_���֪"��#�k y��#"VM���1Z	�]��=�����{s�61ap�#�d���s�k$��"̭k�����i��1Ʌ	>\j�~�v6��u�X��8U
f1�X�4���J�O\�)�ٳ�59�y!T��|	�����u�����X�x�W��܄�X'~�>�~���Ӑ��͖�[ʂ�@��GO��owPZ T�እh��8Aw�'V�|����zʺ�l�ȴ�-O�+�@KS*�
�k�������Z��W~������y�qw7�����C��ln.�}�f�f樘7�	�1�����8�x(Z<�K0�淿H/b�������R�:�K����+A�����{c��H��k;�����"73�~�?o�ş�sf�";���A0���]1�Q5�:&/:`rC�U��)�l��!���_b���y�� �2�R�Dq�r^a�6M����v<���b�e�2�� ��. ��ڶ��P2��*�0��KY�({[�Բd:�6F����\�IJ�g�}�6C*�ԁ�O> �gz��D=�a���ND�^��� ���]��7��,���!���O�0#�%�MJld;;=?&��X(&e~n��}I9
[%GiR�W��GE�r8ܭ��5�W�^�bw�8��G�23R���8��r�.1��c�$'`9��f��w^T&DM3|*����m�0EBi� ����+�7��Own��#Wqjn�}������CU���e�̰6zu����!R�sG��\u�f8�!ok�!�����T�Q0�I�B��>��i�UB<�`77o<m�v�x���q�a�(��zL)S�j�t=�][z>_b��W�x� G$���c=��T��y�z�ǲB���F^�	��4e�К>��xT*N�AD��ΛsN�|2�˶��NF� �5.Ak�Oe�����G��mЮP�b�m�T1��BF�@�	�6��=+����Tߋ���Ѹ���StT��S�s���MEZ���٤�_kڼ������������VA�������$���^�[���
��E�Cd���{:+�R��AU|��'���]AVx�i����h�6S��i��u�ۚ�s�M([����e=s���' C��Ƥy�Ug�'g;.�f�h?��
����r�楎W��E��7H�'>n#e��pC@@�9S/�\�Q�Օp��c��O�ӷ�1�Ns$?�Yz�XG�e�J���ᛚ�f �:s�7���#݈Q�5��2$�,0����}u�5C�B���f��(��X��b@2Sg6(�M�1
��<�t%�r�h�t�N��FM[J��]���1{���_N����+�f/ d����F�t�y�lp���#��o5��ُ�9)�5���6�B�y�˩[t��BsL���=m���b`������G�6T{��KD�F��ړXi���G��J���~蛨OC��:�c��WVw��?�_gq���+�q2�B˷	��Ye����A��~|�3;�K�1�K�u艒�<N$n�>A��V�%i.�i���y�@�})�坑���� ��)̊�)ت��=�VC����Q:6E�J�&<���\|��~�V���Zs�/3����JX��#\�3)K�q&h��՜�v��h���atg����G��]����Ջ� ��܂ɠ3k0˚<[�!��>_E����	H���pj���~�<y7�N
�S�� �D��#�V���q�Ѽ�
i�NJ�7)<L��d����c��HM%�v��#��s�M:�f<�d�C ��g<9��ٛ��Tń ��)��-¡3m�[I��@�.�P^���
��"�X1-μT8!E݈ITJl�0����$�ǚ�/�2F�6؁�����N*�^����,E�g�d,<1�a5-��}����<����{�K<֓��AM��4J8�]�*B5-��'�+�Ƞ?2e�(n��7_g86�	v/6߈M�yN��{Ն�W�(��5U1�(�l.�ۆ`�Ca<��-�HO���}x��G�B*�-;)�Z�O:���Ө>�� �S�6��#���|��;Q
�xT�Q��ﻢ�I_��,!`rMh̤7-H=�ژ<gf6�͎9��yHɋ5 Ɨ
����b#Zxxj�T }��ݙ�Wv9G�n�M���~6:�ݙ�4D�.�������?�rƀ���/��|X{���b�v���&6��5Ʉ_�*u�mC�v����C>�$�ʯ�����b�LT�eu@TL�(�X�~\>_�ٜ�5XT��F�ǿ�-M�f����_-;��h�)��t���|�G�M(�A��&=o�����Z:�{��Og9m=��ŧ!���;p�������>g�t�܌�Z6�6O�1�1T��ì��xn��gԀ���jZ>�[&6&��|��ِ���<��m9�±�Bq��s��UP'3+%�oOȕ��f^�E���I
���%o[ a�>��E;I��� V��Z0���;����h�>��8�L)��+�A�u�2�]��5����ˉf���?������}�z,N��hi�J>Ŧu�� �v���/�Bž�4�+M���� IF���ꎾ^����H:��r�%J�<���X��&��d_�.���x���S6��8�iە���M�@�#g��ɱ�"�F]fEq5��#�U;H�3�7t�$��;W]��7��Moa���]7|�LQ���B���0�`�a�P��ew����1�-r�6�����`j�3��LW���q�G�ѫ]f��x:Ł���E��x*�.��إ�����t��׽Q�Ȓ��e���(�bU��drp�ie1 ���Aү��:���R~I��7��,�k-�H�{ӫ�9�)��[��@�7�Pr��b� �Wa�#절S�J����5o�g(�(�\/|��KFM�I=G(z5�"��x�1xI���C6�L�=#W��>o㣅�����Ə��L�h@�	.���_}�E��g�x�λ#�y��p��)�}����e� Ľ�H��"ݗk��l�r^ N4�4e̅[˵p28��A�q�U�Us��S�A@V[��H�_N��l��8JIYF	O\ ��Ҥd�������~� "Y�b���(����h4ؿ�F�)_-��+2`�Z	�PjrF�����o-xo2���ҟ�V�<]a6���O��Y,=∦�	�؉��!K%%\G�$����Վ�=��L�M@uq��7�5֭�B<H7L�e��@�����`k��ųz�gP��O/�d�n�'�Z@�z��ސt���io�3�'�6��6m6
���d���Uz�[�;rǋ1�n�J�׷t��g�� s̳����`�,7V���>��O
7#n�KVegu���ˍҭ߃>uI���t�%k��P�~>�� }S.����'1$��fTO� ��57�F�M!��,�M��B@�F]���{�`�"h"�	f�PtQ&�tE;wF�P+=z�	m뚘� Փ,�W��$ U�C~&��s!����G+K6`�ã��I�N� �*���ʩ�I�z��,��Q�w�ZW＂#T$��g`��rÞ�:EM9m�`��k1-HW���ڰ9 �.����� �5�QJ&���]-�{V��C����z����=j�U5����3
������w5p@�m�\2�#>��2Ep������p'((n]=���w�,�`��X�ܝ()t�U��F�B�rlY7TF��\U�d�?�:S/l �V�w�
�U�G5ve%�`���ͭRr*�D��(��4� ���jX�^��n/d\@aZu+�	мi�_�l8]����t��x�V���EvW)f�'��a��}h�:�6�/eS��6JzFd��˸a�U�W���0iF�!����@��O���E�ԃag�WY�<Y�x5�kL����d:�����L��vcX/��MdZa6�1<S��N�W�:���hB�v����,��@�����[A��蛔KL"��5G�rv���y�ΘD�����>oE������{;7/�i[X4���z�j�����Wu�t�X��n��}��'d1��aTK�G��=0�q�!D�N���6-�A�4���g8bB��c�o�����K�l�$�~X֝��D�E"���)��r��KT��'5���أ?h���5f�	��d9�q��Ĵr1c6pS`\Q�7��#�gP�^��lβ_�Mf,�����C���o>���n�%�����Vۮu��x<�_�
�F��3g�0 >A(��J�[e��R֍��л���r:�/�`g�l/����h��Hh��~�}�.5T+���K@G)�WaW8�_V{϶��{�kƣ�8\������?�:�t�۽;���Ԑޔ�zxd���4����g�d�,�5���Y9�)��� R ~[,������{�ydt"!��:&+� 	�Ov����*�t�ĖIC�`�h߱V���[��Na�B��ެ��E3�y�����њ������g6�6pT5]�rh�����XAl0�t���*1�צ�^��rj�b�l»0��Q�G1N�J�&<�X�,>�[BmaA�����yI���k�=��M`^P�E���H�L�s��!�ً��UC�=�_�}�2�dҤ�����,�CD��y��$]�����+A�����%n�e��/�X����ńФ+��QUB��Q��BgOB>��o9��}�����`�$o瀣}#�E���PѴX-¢����HJ�P�r���Hh�M�����L��͢R��P��8��#�|�[��5Z,}�	���4p7K�����P��x�!)1ow�	�Rz_�ʂ:�ݯ��U��xy⥅r\,�us�0cL&Q���i����t��&���t>NY}�����cR�<��	:i��� j�0��mU#�Gn<[]��CDQ=�2��K��TQ��Q(�N���Y��ç������,�zs�]��P���q��V8���;�\���k�}9!�%~�������Z�ٔr7 S�aH�!9��#�'q���O��V��)cV{�����@�ԙ#ԗ�m�s̳b0)���V�{ݸ
{]h%�Oְ=�5��\�����m��u��K�+Ә�ͯ�,(h�{{��t9�����c��H!|��+��x�H5.������o�x)fD�A�5Ji�Ƅ}><i���vM-��=��_���*W@U�#�$Fq��D�"i�t�Z�2`�E��|M�K�2�b�V�PI'�`�m��v(�Q�~��g�gVyB�z2���� ��搐e8�X�mdo�L_5�����nA7�-(j��1����]��|��>[�v��,�yC�$�X��1��K���Y9-'�G �j��ғ��i{�y�S��$�H�y<����rįl�'
�6���I�\'�{���sF��E]��1%�2�h8ȼ5+٬�;�G^�s���[�5Z���,�Z�&i�sYl��Ҏ�����]�j�sm	��v���}�,�E3u�t��W�C�]��#��ԙ6�U�!%��
�2�}D�+���ޯP�|�f�'tU�l �!:��t��a1�n�����빃�������h�ά�ē8��/Q����K*��DF�1�)ӵn}݌�.���H뇚��A:M��T�}��])�/&-`��*LQ�����{QQ0�\�ɬ ,�P��y�@ρ�È}Y3iq��2�x �*�Lx,�@%r�-�M!��:cd85=U:^�l�4���tH�n�]nؒh�Ld�x"��2��>�۞pca�7O}��b���qI.)F�����L�ȣ=T߰��77(CH�ŀ���u~�J0�ݳg5����q�jj�E���Sq����뭎��L�ߓ�EA%ԾK��Կ��#H��us�;�R��c�Jj}��������&����D�4��)XB��˷�F������]���s(�$�n������^����tX�-QLcg���L]Ǥ+�VӴ�xQd�&�a:})�>[J�^kE:�j��4�[ �O����i��Lx�pJ -�����,/
3��Z��Q.�\�BF����S��w�#f����r��Za�Z`�����8��X�n�*�m�*���;4�\��Td�b�J�J �m���������.��3�B�����`TF�����Z���:�D��bv����FxdYre�m�2�#\��wp�sN��w�F<�$--�Z�R��D�4 �,%�P�5�:�z�BM��Qԩl}~��B��V�]� d�L3�d* S#���v=_<�4�{W�$�Ԑ��S�M+��Y?1_B����P�P#��0�#D�����AqK�w�~�誱U��r�x
A_!�;n]�P�a�F/H��,����T����W:e�'J�uI"RPa�Y�u���;���X�1�a޸/����u�!���|0|���\��7]���>��T�3���j�D|��Kz�6�&TdH��hS�0!k�|P�
�u?����Þ�f�qh/���9-w�Wb���b��4��6��|� o/��>}Y��x��T$���B|q���3��P8P���a�lg�Q'=�/]u8|�8�����`�E��v+���V2��s)��"��F�"Z�T=���e�L�uFF�6�s��Y�+���>�o��* c�FR�Rܰ4�#)"S <�`��:�)���8>!T�ɗAC����,���#gjl�B63]9�FՑs��uV����#��ז��lFܰ��"��o�^'G1��b�{Ap%�ƌ�S�Z_����J��Z�UK�-U%��fY���s�z�Kc9����5�f�m(�U1FШ!AY_�RŘ���MN.�tc#B.I�O�ӭ�`�7̎}���Pj	ul"�^4�I�Q���F"�͑_`�~U}e���gY��Gq�u���V�S�C�]��k�]	*	��~=��e�l�2�룐z`_� hk�W���!�h/����u�:vp��`��p^�]&�\)Y��⌫t��Q������w���9�<�`�."X�Q�L��-G�����ݤ&�筟��	[���O����n�շz�᠎"�u!\�4�
AF���-��1��h��'�f?�7�L��2����Պ�bIӑ�%��5�8�{u�8��u�%�F@_��@<G0j�E/|��iqc���2�ּ�rC��\�8�M�����v���q��kha���1�W3j�p����&��6��|OX��O��C�`����9����w�O��B�kB��Ş)F�����&v��L�V��[���*֨#�8пX/hD4�AC�f5�?�.=�lw>D��;z��Yk��8+B}�xj�p)QG�?~���[�L��;�s��F����c��s_�a+eH~8N[���M���m��߃p�bۻh�%�lo�?��oh����T�\��Z�(2��g��`�b0Q۵�\��$α�mLM�x�u{�����l�f�+�4]�)pK%/���9C}/fIO���N�=��5
�]vW��!����-V�����]#��m�-�/��L9�`EZ��0]u�	��&�\h�q�F�Cd�����Z����9Y�n��)�@tc['YQ�mj%�O� ���i���"�P
.âņ�l�)�m7W�a=�CF1��CY�F��?4;A���S+Cw|o�Ki�^�A�vS�TM�\�d���H��I%�>��P�Û`%uC
z	�IGߞ0��?�R�L�adކc�)INx�W����"Y?EF%y�<�
�D�e���͘X ��5F:�-�� ����ޜ�"1�b�я�`�lyw�>����{i1��F�1%�P�`�W����8�l�_�<����o\9F�(��Hׄ�
'���m���~c�QX��tkʛ�{������� �Bֱ~��b����۠����V�V�������	GS�+�u
ޚlR�N��H�/�vAQnDq�/�O��S���۶��z�<�kl��]�L-�8����/<x���l"����T�X��\`���s�iϹK���$i���F6�w��8ݷ~�CJ����o�43��qD��PZx���,���Ot��R,����;Ր&ۓf��q�|��D�6��F>��JH�4��Y���6��|Zr�Gī|��gE�+z��K6�0R�R�"���i�5�b~$�|P˩��Yh=�ѺK����HE&';j`:@������HK@ܱ�(23��,:�V���n(�����񭻛|9t���+b-C.u�˪��N,{ �~��x����aX*���i+�^�+pMF�~�-�1�������MW�MThn�O%�|{@2v! \�}��3�0z/l�t%M;v:e��ﲓ��L�w/�[I�ս����5\w�o��H�-���$C��Z�m�K$sq�2�/��'Z,��	������խy=�NƦ���A���GI��v�<�A��H��}x����npw��׫�8�5�c�Q�$����&p�)�*����aYB�T?u��N*3���r����LYm��/�˄�>O�������*�_�`����yJ�,�K�b}��x����O�78K*��
:��S��Kv����;4��~�R��s�'�i�������9�8;~�!V_	��=�֔d�~����ք�����Z���O�����a$���L�4���q�(@�TRd�Bj^�Z�R�bgOz�3B;VB0|��2ޭ��Y8:�!nm� ����s���ﴞ�q�PG3���0�Q����]hհ�,�F��
|�a�I��6`�!?��4��J�VY�d�2��<� �̇c-dsi�M�B��~A��ԯˁ
PRk)S6�J�=^�(~q�
�Q����5�is��4�⿵rM;���:(t����J�#����F���^ R�?��%�%�C�<�&���tE?7VLcS���:�8�	��Q�u+6� ��_�Eh+�Ùb8Q�����߽A;����U���b�K��������&�.G�x�W�W�s}�J���[�`�A1�;��ī�$���Һ��:��)��G&I�3�{[�&s�b��N��-��2Q��pM!?j|��z����[�̘}���Q`��J@�)�=�w.p5G�8�>	?p��͍ٙn2Sϔ��R��i�/(��_I��۷���jC�{=s���m��.󖺙Lf����0�a8 �(;.�&@�ݸZνl��(�����u����v��Y�����(ײ��	{�yJ��3���o�45�J�K�a>lf|�MN��MZ��#�Ƀ7T�lrs�;bʠ��;Y���^=����1u�a��DG���%Fhg���4)�ۋ!J��u�cS��3�B����BƤN�BI���ꔟ`Uӳ�'wg�
�ګ7X����/�-�&):�"�c+%jU;i���N�}}u(�1,��s���8X[c8�1���h"�o<�T�02j�K�lZn��dkX�If�F����׿���m�s'�V�!�a��vS4H-ժ�{�-�--7WW�!�,�z����Ǣ���0i���h��K1�}�W�w)�o��=`�~�颒k���}�,L/7����κ�z����\�囒��$cƗ=���>����+��xȉWQ8�P��tUxDc���`���U-{�]�W%�Q���		�KR �*�Xg"�QI-^�چs8�x�룺��\����(z��K.���l�#b�S��k��UH{�[����Ug��~��7&���cȸCCO����y�����tmW�V.F'�q�0LO���(���#�sZ�)gׇF  ���XoqӶ=���S����u�otdp�A���)���9��T+����ф����b2���$��!��[����
qq�t�;��VH����[
����;�G�`iX��LI7|�V�`d�)�4��3�c�3�,�h�λ_i�k�J���,|_c�S�Ǜ;�DgC2�̾BG�xm��p���6��r�7.Ӗc�]�g�q\�n�}gP#����&���J�K��O�9ϔ���-�$u��>�4-��!Z�fv�tT���d�6�u{C�c�����T�z�̺R5h ��#C�X�-��������Wy4E����6<��-�ǀ���n?��В����]+��?�P����ؖ��?�M{�j�d�W��6���i�3rST�F��&X=����A��������
ӧ� ���m���F�+�h�"���)}}[F|��7����l�ٜ��*���Y��<����na��	]"�Q�87�
&M�&�V�&��8�&��F�r[�WA�;w%��>ӝ������@&뢧�gH�6.�I��;�,�բKJ>�������O�� ��q� Yߞ�u�>o�8Ҿ��hrG��P�K���禝��ʆ������ޮ��~L牧��QVZ��ؿ��t������_3����7Z��a@ӡ%)�� �ҵ��*[�ڻ&��;�WnF��ű~���,��O��9���5�ϑ6��C��A������w���2�ޟK9�h 眛m�����5����7j�23�~v� }����4 ���|l%�+Y�����oT���Mb�&e���s���#Q}]�h�˩r��v�;|��˗����g��k
�EW�0�l�{�)l����B5if�/}��s�-�R2�~�A�]2��A�@�^N@3q�w7�e���m�x�u��
�3��RK�z�b�����d ��,j>���v�rE��ޯ�T����ew@~��CD�����i��K�p�HdH�й��ί�$�7;o#F�D�~�n`����h"�����v�.���=���:�h���,�вO���K���<�p��wi� �q�I�*�'�rV[#�������\�w����`��rP%��lMVL�}���K���}c�\ך©�F�������/��c�����ږ��>�2R.���U��q)��?����Iͤ۔����v�V��6�!+G������������s�K|���s���.��2��	��JW"����F�7��m��A͑�"�IR�Fl�d��&�<*ؖ�0���T�n���+DV�&[��yXo%Y���p݄�Cr1��w���L��� +
��-�뷄c��P�5�hSY��
}���+��Z�I}ѿ�_�m�xt��I�N��l���Ea�MWT ��F��fՔ!��d�t�rT��vw:�N0�ID�6V���㟕�+¦�]fڤ�O󿔧GU)�p'0�zu��T�oQ+i�N��������-��>��L/��N�������c%���xځ����8�S��y�)to���Azxo��x��+![�"L��~�A�� g+�{�i�=a���ai�E�WULd�����/��AJ�f��sgց�{���I�8^~��Ş��$G�9�]�r�خ_�a~��k(����t�̱V�<YI��m���B_j��+����ܪc�O;�!
Qb�"@��$��
�g����V�MN���N������4=���}��f=�p\H��Bn���'�,�w!��:�Z�Uي, p�rGfo{,/(������`��$D��$[`�X�G��Ӑ���B�>�/�*�W��[�_�6o��#�L���ٞ/�v6J�Sa�D�!3���r�_��8̛(bF��u'��Gq�TDY����(d1\��=�d,�<o�w̽�/���{�IA��>�Nv��萆k��CcA�`G����dD�����B�D���P}�dp��D�/I������o��'�c���z7OkJ
]�b ��U�&ݽfk?q�<��6;4�SK!���/1��y$�s��4��#@��{�;BT;]�Ǹ�t����s��z��ʥ��j�~��/Y���
7b�H��Z"g�e�%�T%A@E�L��R@���W�˟�l����?�e#/	��%	Oj�J_!E�)�� �T@�/��݁"R�#�A;�k4,��퓥�i7��1�.�u9����i�ل���Q�3�rp����h_���\�Dpk���4�f��!v6+�I:n�A�����G4I��m���h�}����=���5�q$�K>n���!x��Gt�d`�]A��bȲ�e�?������+�����Й����f�.����$�+�$,�שh�Bd|��Ƿ���D�aYc�:�цUdQ�m*���z`���u��mV��3F����=*�0�Ė���ux���4�����Q�4c��%7�ϭ��$RF���`�g�4Q�yq���\���\E^{}�_,�Y\�?jg�-C����N�-8p=B����[���&�k�Ļ��?BU���#�m�~���ƺ��p��<���&znA[Yi�ܲ�e�1�L�~���jD'��`��u#DīP��6�L�ڗ
�����`��.�4V�����ɕl�irI-�u�a���#�.����&:����*�c��_��d���Q����:'���j�W��_ӫ�?�����W����� ���9��^F�i��<u���$E 2��#pǱ���sW�k&GI��Q@�Cd�C�tQڠ�W�o�ň2'�Bh /z��z�2�g�b������mު���BkT��V|VE\ٙ���V�v���Z`g+��N�h�g��]���icLf2��䇞-F��!��󗫂�|��=�V-�K��E;�~{Gy���﹙��L����n*��H~�,�I[�c� ߊ�)��I@�H/�\玅��_���\?��'�,�4e�֝�����ZŵY�
q�]O�$�������x<N��#;?��7�j����-�@i��'G�K�����]���p�K�y`I�S�6�滈���L�G�/DdFbR�c{��
n䕏re[R���Mta���&ET���kˋft��'b[�7o��2�����d�͊8Ǆ��f��%�]<[L鱍�w��
��ZJ�0#B�Jh�gG���N�_�ݪ�a+H����%V<�.B����r���+מ�5������r�y���FM�e&�Hf�Z�"/���L֭P�:�P�,����:k��Kf!�`�	�ΐO	�#@lG[�d˵m�L�C�KR��[S�[X<ͦȾ�?Z�`��������'Xl�u@�[�V#�s�k$"ںb�J�8\���y�����Ո�n���,��Cr���C�$�ƢH3R�����
�X5��� ������6��?��3�ٺfWT�Ia�$�]�{'.���ҏ��1�FeU]��L�8�<��{E�cJt�\oL|0�T�y�w����s[o}�D��$7�n�A��P�'/��	�54�2T�|����|��IDL�q�}yW`���}���0*C���M:Ĝ�������]�,3W��Un�W��봨{1xY�U��	W-�m������QRϼr�r�/����2mƈ����ؠs;��#ۛ���}���9{�pwK������Pw�q���l,�1��6��Z#S����%-4�5���у%d|w߬�pB˓y��ٳ���0-i�!r�a�7�#�<�Z��fo�n�[ȃ�m��������a_T�>(�]�^k��a�2���q-���D�َY��|��.�#�`A����G�;k��4'1Z 1SIPMr�� `��C��M�B !	��˘Y� ��ɂi�*w��t��+�jq<�8m�°meޗuY*�,��22��u�TUQ��,�v�
�D�� �|N�q�#��7��.	�r�����a�S��׳����ϡ�',��m@�ږ���>��@_N2Nu�gǽ��3��C��c��|B����.$���^{��)K!񌜥5`ҿ\�G��P��\W��y��sc#�����
s�)�l
��\,���UL{C%���#���X?&�e.�o���&q��ye�>��q����ٶ��C��y
Nє���]�'!�-���9�u�d�!��my!,��b�6�;�yZ��}�����Y�������� ���[�i�xS�!�VWWϙ�cyL9��%��{;�Ƒ��;'k)l43k\�!II�*lg
�q���� u�<�xh1��lx�A�*�m���S��<��>�Ƚ�'Џ^�����/�[w�$9����K���p?|o��XL�MI̮{���ii���9.�ͅ����g�=�A|�p��T�*�&A��� ���/�8�ӣs�{W��z����6���[x5��9Kb���N�y��A�C���*�<Jz�1����O��hX	"�ui6D�|
,�񯯎�{�j�-��KH���P��QF]����Jbؒy��ִ)�}a��kFv������ZU\��i@���P;/�e۴�Rɘ��'3����������Z^Ƕ�0	Q�r�0����O��b�MF�;�)��F���9���"�}����T�_B�<��}�Uv�	W4\�E��{S�	�0�m�c~�'!�c�%Զ/�G� i/�7a(l�aP�}�sۑ{z����bx�I}l����B�� PZ�Ldc�!�Y����\F�>��f��!�L�	P#7�!/�6ǀ���qsd&Q���Z�G���H��n��a��/Y-����d�|nq\�ѳӹ������g��ظ'�Xcǻ�aƌ`�0kp����m);�*�R�1!�?�-�(��>�.|y�tSgF�R��je�?紥��L�ս�ok��)zܙ�%.�\�R��{���^hO�<MXٞ����A' 	N �0��s�0���b.�ξcH�B�#,���V����@@��[q*恧?/Q|��6ߑ! mq�tK�'F����FZ�Ҩ�Y��+fe�[�Ê�t�NY��Omh@K��������g�u��RW���r�;]柵3��_���i7EOU����Jy��S����5V�I�'�v��R������4e��DZ�,�5�Y�;���Svf�x�Jqs�ʔj����=� R[#X�N3��2'	����>G2���>�;�9^�+&�jш������/����ǯ�
���.�I� �ewqFͽ��r�%��n_taؼ1DL�E?}��q�3*1cP����0��>Ȣ�8ȿa¾!s�4��>��	,�O�+�Wf�ȭ)L�G�|>����'fm��+�0��/���#�fƦ��1��^k�w���&>�ذ}�Zr�j��05G��R�����E2�	�
|���َ�O6��nz��D5p��?����<X񤛥=k5I/3��[7wC:�v���1��:��h�孕��$n�R��B�1��om���f���n̶�u�kb���y��x��x�f�"�ۿ�HN$�J�4�2ػ�<p�㥨b�t�Z�\GF9���.���F@������l�x���ȆS�_=�键���5���I�=�3��vst�8�91�����<ÏN0$[O :�g�'(�!&���=��N�Ѭ�I(�ER��5j~i��.1��>���w�D-W�.�}^������{;ҿ���쇨z,E:O��|����j{�%e�a���/�v�+|�ί/�1�H����N�*�q*��M1����_~$L�:�P�#aaw��ށ��@V-�I.�>y�V�Z�R�N���2(�=�O�	��oj���[��bw;��c ��#��P��6A�L�+�{gM��f��B�#V�o�6(��$M�ˎl����Ȱ�7����od�I�.e�{�ʃ��w*��:��VyH~_��z� ��b5�㜒��*�F/1+Bm=�%�#�3_��*�
���**nh�<�Ķʙ�)���}]`�l�K
4C�	�E�x�����ęp��'l��?�Kk�4l���C<֌��.��@w>��� {K�!��J=�\���&J�|��gT�R	vr�5�M���e3ό��vA�Y .�k�cS�@���0��W�����ߛC H���a����6�G�fD3�u����d9T+�f�.��E�`������eT܆޸jrd_��Q ���OkZ޾%e������$-�p�@ʧ��F3ƣ����>�ҋ��	C�����cJϯ�<�S�?J�T�Y��"���+������Kp��@�H��đѳǱ��G�稫�f�_�մfq�Ǒxb�k!5����X�854�f�f����������;&_���@� B�͙��0�u���ۏǪrv,5f�ˢ�tB$s���'��O.�{ �' d��"/{V���@��t#kʚ��M�9\�0���lV��$V��a��cU����Ax���L[6J#xp�߭�(u1|D�������S�Y�>���@��*,/�������qQY�/�Swݲ�up8PI�A�o���\��^�WB/�g>߆�t����p����o�I��:ܱ�fi�����8n��h�`1Ҕ*�cϘ�e��G1�0�>�vӤ㸤8_�K��кA�﯎`
����;H-�1x��r�U�j�T�͝z�.��O��Q4����J	���`G���IS:ϊ����&<�Q�s�ٕ�&_���ɻ:�i�[!��W)}g��Kh��*��"j��E
�2}��W�(L�U�����bM�whm��Ώ�;p��hX�H�mK�����&=6S�pbTT�W:�䠦�Tidh��`.��)-~w2;=�A#�Sv��?�</9F�{]WC���L���3�R��uK��מ{��G=pt�ӄD��i�}�޸>�����\�>G3�vPv�>Q�$.���B�n&��ůt�&S�a�V����nV�`��k��?ڻd���{[��ӞǑ# �z�.^��j�)�%�|�[��9[p_��8��0Ҵ��ç|jO�Pu�Wz��P���;õ����o��}��=�#<V*�o�+�����@����pQZ'S�#QM�)4�RLs��_Tt�BXҏ�q�X�)\(��j>�'��+���B���)�L�7���A5��yG�I1lEW$I0��U�q�Z=���y�8۷ˆ~�n2�Xej�@;��9&�����z�V�$s���X�[��}�"m�̦9�WQ~ʎZ.~�Æ���Tb<x~gCz�S��/�p~�/��CJ���~g_%	�Ԃ�(�M�9�N��aS�$�\^P���U����`K"����x|���ܚ}^qN|��{,���S�����ب T�}�ƨ�Zwl��<v�9~W�����D=8���&���L�v�1�U�݅XL��5��r�}-@�ђx	TW>�����(�e�gp��_�)ܯ>|U�Nŧ?%a�e�DF�r�m�W��F�i9ZL�<�9c��'[{�ky6�(:A"�G���.��]�L��]�ה�V��" �Kp���K;����R�h��\���#��$�/HuCHθ�@��.���&L�U���;9�/�?8��_Liˆ�f�S�%}�N3�(�%�OGD�?X��3>���./b�Zb�w��q����V��j�����D���8tA�4>9)����y�7�� ���(r�����Y���İ����e�%�Jak�n�ӱ���t�d8�.K���"��4�ŕq*+-&��N� ���EnD��"��5G
����fQ�84�`��f�`;He��}t}�M��]�����)r���d�+R-�&��J�Ab��J'���zs�j�I�&��o�J3�w�d�~ݕ�{��f/��D�۽�U�Z�8�?[���s��}����Y�-b���<��P��k����I�E뛜��/
��N�W����Ns�.�P�f*}��j�9�ݾ����\z �n���a}:'����0�/�L�2��b&��'`X�a�'[�M���쐖�0�Qs��[� �v-��ȓ{o�������*��R���Ė����L5�e��
`���ąx�i�.�@@V,'D�9���&���H!�c��y�ɡ@�|�����PA�4�f����T!� �,�V�:=���L	���>��x������W�� ����_�V�U��)��&��m�ehQ��3�(l���WO~��=���'�q����B�jܚ�F��ԑ�i�A�k�y����W|Hvy	[��'�7_)ˊ/�E�~�C�=�R&��z�2p�2�ۙ!�d�*ٺ4�j�)��t�i�(�S�>�)�ټ#�"	C��U���]���{ߝ��K�uA���H�ӟ57���|�ήV?HG�wOt��bb�=���`�CfF^�bΰd�؂IC&��ďW�wߥ��a�2[)��w����[�m��r�Dq��QJ)^r���v��&e�ছ3��#~�n�Q�0�]i��	��1I��G�m"{޵�7<�7��p]6#�����WMID��$8FN�j�4�N�4�����"p�\ݴK:����t'~<��jv߄�q���#\���_{#���¦�Y�ie�م��T~����o��<>Pq�Mo�LQ�/a��I�] _2P���RX�F��V��?�M�>�{�p�D$(�\�|��&��! ������pu��Kc2؅��0'���DƔ��z��k�+�dEڗ��^k�˲״#��MV��N h|	
������f�����A{<cxi��7��&�ĤcB�Ln�Y���a�͵6����F5�����ݫ�&-j~��~�軦	�����Ȼ"Z^P����R�VF�����=n�I(K-���(��������!�_���j[2��:�6��RR�
��v�0� (!��a�6�n��ԑ��f�-�l���'��6�.v�,����@\3����8�K���xOf/U��`W�����L�+���	f���!,a><֍� =[���
a�����YYl�mE���𸾨�Ύ��lG��#ie?�WPo~�!͂krtT�n@h%���� B; �6�hd�<�����--0o�0[�+B�.�w���-NAd������G$�<랧L�͋2�����֖�ܔ�iCLu��@�9�.�wM��PUn�?�p\o3��,x���d��ͣZjՇ�I4��S�����#�ȟ!��O��U���;�����٨�6��wfd��
/��nH��g�{o�2�$��iŤz��C��[	���Nȷ��Е�+�xE�������)�BS;�o��=3F�u��Y�#�7e�V�g�^�ʙI��-���u=��&=Ym2��Ҏ�8c����:|x��5��T�H<���*�8�i��k�����q?��k��K�19x��^��Nє:�ǉ���M��{[�x�A�fv������hTSv��=���'{I��q�!�����Zp�ϳ$"��)�hw몘�E��7U������13��a�,F�f7|��\��2G���3��v�s7M��ק���u@yg��-��*Xԣň/�*H$��
�z����k紛�4���H�A�[64�ibt��?,��m�v�y���<������4�����yVq����,c
�7ўq;����9���ej�&,<nc�堐a�hVzn����m�I~�H� �I^�p�������'��w��L���=���f�pGP����e*V��Ptq~)�e�E^ SR1��)L�&c�t��9�m�ڪ��>�Et򙎱\2�9�8�Cx���H?G�����n�C�J�r��u0�[(��4�[vO{h>9;�cA�W�[�僿��7`����J���E� F��7D"���$¥��08�E]��0(�\:F��g�����\�w6��f�n��y��V�Ύp�v�U)��7�Tr����3��*�;#|G��h��O�?'�=�]�Nh��b�'U���w�4�l��S\��D�&��(T"���$�|њ{)}T|J9��}�9nJ�1�F�_�����u�jH����|�ۢK֞��?wU��Ȝq�3H���"�c׫����r����`T�l�!&���z���Pv	��4�Դ�C��er<\�����3��{Ae'���ɹ)_��W���	v�+�&�˯T�j˶a�)bBNL��X$�r�Rv+jV�j&��;-��r�;p��~PŴt-㬦����a&qh�M����1��]�?.zn[�:¯�M��-�hx&ᕴ�d��"�ŵ�)lL�&��E]Q0��5�P�� cI��UQ�6��$	`���~����v����o\lwF9���sG.9p��s��MR�4��lLb{�{3G�n]�@�[��@0z��A���37l=�J�x�� �t���PHBEoAX���G4��ci#`�h���,#Ky'�БA���x��/����_�%<.@�a9|���*�|��}�;B���!�~҉��(Hɉ��q�^��cƩ/q�3):`N���w)��4,n寋{�"JP eg�[�c�>��nǫAK�d�ȗ�Ծ��Ta�R��^˪H��� *rܡI��������=�. IS�!���H�KH69j:냗�ۦW��W~r<��e�'��d�V܍M02��h1��{�	�?%������ج��#o�8}�T$rGc
-�Q��w�� ap�?�6�]q�G�&�e�m��I�bJ7��/��~��ݩ$U��=qψB��G��h�m���7"3㗐l�����[KM�0yBy�)�����RV���������!�e9������`$�a�6�'���I���2�>N$�#�����<&�, i�2$�g�2 �I�&�*~¨����,9!������X��o
:5�/�b?a����5��_I��]�1�z�`Z��6�$l�� �e�<l������	�eT6 %�}�m�t^cGREg[��kql��^s�'�P��{�/b���}�����7_#6�QSv��w#���3��o�j6v�����wj-o8W��x�\�i�M���6�2\�g����BD}�.##}����#�o�K6TN�	9Yuݟ"��Pb{	c͋*qB+c���+JA
��i�Z:�3
H.p�P�����J�����Y�u'v��#�����������}���ƚp>׾��㞈�LN1��P����V��sW�7~�aig.��'�ܰu�aO1� f���A����3U���ۥ�z���*��;bSz�&�Jn��O�s���u��ہ0пr�l?������g�TTrƆ�'=�Y,N��o��'��IK���-�y?t[�r.pf�ņ>�@&�$�A.I�����}n�u� ��bdMc4�:%������o�!�Lĉ�ذ"O�-�Z��*��ڟ����H�3<�^�I1���.�d$���=����4I�F.�/���
*�2�=)g�'��(}�^�![td�9��D����:�P�	�Af�bг<��p0'sAX���15Oy�HL.s�o68�]�g0b�_j��D�i[�WR���o����ẁ2I�~��Dhֺ�a�/��%�Е�	�s�ͤ���`_j�DM9Bi�&���L���#P��R
�Zt���C��z'��,�����Q.�[���rW�����:��]j���q�dS�aIW�����4�?_||����iU�5�`��!�`dn�ikC�� ⅘^��x�$�K�6m�0G�%OqG�(ME=������lۨ��O�9F���D�Q��ˠG:>�>��6��b9?8��Lrd�b����Ls W`|A�Z�)��ÈH�b�+�gO�p�G�[d�����'�e��l�y@>3/	#kHq�	@>;(�5�h����n���3w`¤'�΃Ζ~n�� �9�>��w�g�,ĊFc^ %>TXK��;�������'����բ;n����5��3�#q���{�)��R������?��
���:y�T/�ʪ�3�&nS΅�s��?��x9o�?Hm�\�v���d�M/\���=z�+��Β��)fG��*��o/��)�����S<��DI��:��w��¾���L0 y6���r�ڙ@l¦�!�V��=�+�p�V�6M5�ܨU��tg��@�=���l����� s#��b*Z��׽�\0�4)��%:Σ %���B,�^:ޑử	w���i�5.��rlX�U�(�c̀Y!�e�sZ��������b���h��y���C�����D��L��!�Yo\��3������
ݟ��ciZ�M�L
���O�I�ٕ�X!Դ�,Wy���������y�j���jc��j�*��൪c�[#���N�ɐ�u�Ū��g���mv���p��Y�iܜRZ_��<f�Q�}�J�v��9F5�Kj6��;���7>2d�:������3�u!)/���B�Dָ����=���N�����܋kFF_��X)��
@w�w�0m:ݟ/!8ԌR������h$D,�<��J(�AE�1xC��>8r�>:~<�l�=���{~�=�B�m=YN$�{#bc�OlCN�[��@���D%k��
����fdh9
�->��<�m�%D�L����II�^`�W,e�qZb�k�V)
0n�o;^A5��o9��R�
ÇY�vi\�=�V��J��ԒZ4��`�h�FJ���Ϯ/�zb�`����_�s�O�S�9�z\K�����F��'��
fP\��z$�uY��OGo��?�:�p�J�hx��k��?W����H��F%9����j�7�Ӛ�0��ަI����ZD8v�-�������������M���LU��I֩���Ab���]AS y��"k��N�a"���|��ʈ��A�s5?3�K�����@9�X�d���-�t5���>��,6��{�t� t���A��o�{�z*����:Htꥄ�i�@'���O���䧾�x'�ZQ;P�fר��x����h���Ôr\�?/`��E�Z
����j�����]̠��1�˧�����;��\܎�ƻ��A�ל4HJ�T�a����U��E0N9���NG�����Z��%%�c!)��:��Vx;���W�����Y3��w��TP���0^�_5���b���w������%KD1�U�df;OM��ek~ l���l উ7��G���bh L���03(����$ף��B�s�}B�S$N�( ne�\�D{1�%>���T�>�9+��>�ٯd#�����G%����o����'��B�wW�fzbXZ�j��`�C�g>�8`��4v���)�*D`�s.e��'-!��=����sbh��s�/i�V�;D�p{����:9�
�~2��,̣��8�d�̍h\l�{��0�F`��f��ҤJ�-�aXm<��79zң��4�Z��` �w�%M�'������ut�qAf��I��+N�Y.�A���������WW~����� 
�)μE�?H\���M&7柚�U�W޼��C\��$���K��'�6W��1�>~�0��Q�p
��M{qNW'7^�9��CF�=E�(#�+F���A��:��e��iD�VOr˽.��$;����e=L�'S�����с2�⣟!9��o�y�f��n) Y�L���1*q��A�]��p��Z�G�D\wT�>�� #5+<Zdn0�����XU&��5FF��,Q�7dk��A,i7ό��b��s�1�B�/�
�_��8�V��n	W����8�d�3�4�LH�S&�y@��a8\g��6x��M�Pu�0��!S�%�I��Q��/ޖ�7��R;�IW��Na��䟴�"&�r�%���ڎNW��C��u��
��ܛ��ʽ�P���}��!&Z��%���D�y������J�(?T�aln�)b2��x��N�����ӟѰ��<���g]��8W�6��-I?����]զ�H��r�ٴZ(�d�Y�r=A�v�"�A��?ACbt�@�<K���>��>�W9/�_z�Ms�a��}O���ν��,��`
M\c�n�w~ �@J_l�«�,��P�=w�<�����gKk"�����*/:.p���C��#,b}�a	,����?x��� �2�����-ѧ	."L4
�?54��_�p;�NCxDu�y-t��pڝ~бYW�>�*(a��\#x!-/^�$4��2|��v���=����!���e������D�a��Vos�a ����H@Ѣ����N���G���toB���T���7�{r��㤴� ���O|j(�fpG�
���0^L>�H�@�&��P�����'K��r���Ǳi1��E��,����pcEnUe�®^S3C.!�3���#'{��F��B����n\��T5��o	y��y���<�T�y:��i����yG�4B��2-����x4�5�O�Aq+�E��i�^U��4>�c��e�P�%������:�����?�G~��K�왵+X�Lزa,]6����@ -B�u(�.��.�=�-%���p~�-�K_��"�ջ�Lƫcsg(�z^5�M�?�?�ґ�wQE2U�6h���0n�u�t�CA>Q}"��D����XxJ�tm�m��k����ɕ��[_��$A�8d��SQH"���BbA���̒��c���m5rt�93���I�Hpnp��寪�]�5JA��?�0h r��NG(��vUlf�<���~�P�3�\��߽0:�l�l��R�H���5�a0� �O��� (m۟� H��-�a�H?�EkC�-m�fw6Z�1��XP�����@{�'3���}an�e��A�����.B;�RvJF�]-��*DycV%�؜�M��#$�]�
�t$���t\Ⱥ2j�a����#���,D���R��1�W��D~��z�:�?��~pN��'^T�B΂b������>��2�ݕ�.��3+�"a�Q��d�� ���η8��)JD�!�����>q琜��r�%��-��B���'3 �-�]��(��CW����O�Q4��$#O��5��u)l�p�!�+�r%�B3�CpZ���6J�7֓����-��{e����Ʉ�����I�j�G�\b-y��*�O��	Z�y �N�7b�
��7{aR�=�Ӌ��h9[����A8�'?�ŷ�ܜ�q��	�����层�zU��u�
�;�kF<�~��wF9a��'���+��e6A�����>�7��$V3��vo�	���~�/L�.�Ԝ��&7Q�V����Ⱗ)ظ_�b.�����X�H�)�a�-�����8�������xdŢ�m��ެ���LL���h�\�m����_O'Y����,��ڷ 6؈C���(ѱ�.G��:A��ڬ��vU��sͽ��ň���G�QbE�b��ѵ&K 3ayR��� �0=TwbV|��S+�`g�v����w;u;3YQTĝ��E�8;}�R \b��l��${w,��oWP)Z���K��l��E�t�הWh����m\5=������;�2j�������|�!�X]�����E�Q���������u����`rvd���;e�܅9
x�8�`�_r��f�Z1L��d�r;˃����k%A��_\�zO���kwHC�PC�3aĊ�̤��;�4���љc��{���X���ӌ]ϖ��
XfIb�������m�:$�Ur�By����z駏K����D�?.��%�	4n�cYY,��?�H7��	�-��~K/��8<~�-��J�	��\d�����=C-����8��@���|h��H��?�L���Xf�f�"&�I��V����۞)��+Nne�F_̢�;)�����ʕ��g��'4hÁ]ԡ�^�T>�s-=�FjO�<���vAP|���A��cS�r�{K�ە�[G\q�̚eZ���&+��lr�J��V�=БH>g����	�tu<���~jλ?}�E,L�E޹SϷ�s7ު�u⧠�������
&~�a��"�N�?��A7�E���w�;J�&��?����e�Et��f0 3�{i�r�z�\ �E�
��tK.W�
��Fh@��F�ac++�?�fj����4��g�q�����ہ�p��6U�����5e;�Qv���T.rdRޛ��3?���n]�u�,j1	���#�)��;�w������_���8M2��>lI�-"�9q>X%��J��`�}��܈/�z�z�1|�����AW��}����"�d�SI���W����cXjW2Dy�):_��J	S��ɠ�i�?�VPq�؆J;��[��O_����G_nbRL�y�4�=R��w j�jn�l��� ��u��[��l�S^�Xh�A�!���}�z��*P�u��zds������w��T=U:�U(�H�b�$�\5���/F��C�������q�]��(L(rK�@�̱L��8#��R�T/ȶ*M6؃|�K�'��9�{^БʜѰ��_��i�6�jF�E;p<�v4Q��^�q�m'Y�x�`��jlsȨT,�s��/�m!cj޵�04�]U���'9M�@E�I"�US}��K:"���&±�cI���Ӂ`�
��x�Ȯ�1�����9�?�؀�~�(���2s�Xh��9��*��k q�y�U�|4��!��f��l|�'�e&��/���]d%q.H�u�ӊ�W�],<_���m������t�ٓmL�݂M��|3�@.$4�5��ep����M�v���RcMS����:�p�ǃ��O�`��(�\�S�ŎA��}��k�����d�X�CN�Q� ����u�t��S[�l���ێ#Vt}��w((k��VQ9��4]`R'K�8.�sN�K)��Ea��zlbz��ّ�� tM�j_�ʬ���|���_��7�Z\��(.&m�w9+q$��>�6\���G��{�)��)�w�$2�`q*��
��o������Q�1�OjV�zd�L�dR~�	~���L�RG����]p�5R��}rZ�z��F�+C��B��W{a��b�-N=�M͇y+�ϙ���;��x?�YF�z�\��*H9���쌼�j��bP2���()��e�Mâ�f�*��\�a�� Q�f�ɯשA��x|VB��S��d��vFQ��x��v���H�ģ�H���:ڔ���~5⫫{���-'� Yn�E��@	�P��H�|�/u蹇k��S��쐪�w
��q�nbR9�}ZnzbA�n��Eǖ�z�o���{uqr�
}�����@F�K9�]'�ty��F"Q2����u�!��_˫�Ly	a�W$�W���>ӫ9�C�G�U<mB����u�E�##Z�0���؎��-X��q�����]	�����?5��o�����9�@���_��G����]�W��!$J�T)��~�>8�J�Z
1m��ݘ$���m��O�Y�0�G�M^��ծ�0sc���U.��̑l]=V��ָ�C�.�s�Q��(�����N��b�w�g��R��RJ(����lv�в����}�UE�0+'fn�(9��H
���wD��K�;���ZE�]0�3�4�Mg7�xl��Y��`���i�@|	l���vL�$�B��9�����y5�R+�D�a�a����.&59�8Y�x���6i�^�w���$�S�INjk}��#�?z�;0{M�C�[����2����P��0�[�S=,}�y垧[u����������L2w�8�cy{��ؗ����=w`M>��<�IZ\�G�&«K�9����Sо��N�(���W��c��؝Qݍ���0�pa5Ⱦ���j�#����&�RnP�B��/K^�8�*J6_��RSd�3,���՘A˚�ٰ�wv|Q����θ�7�&���\��p-��rgɁ
zb�&���fc�I�P��2�ݽ��.�ε���MN����6��ʅ���ޥ.�d��D�$><m����
 )�u�+<���0�߬�\={̓������R�dy�ƕ�8��dD���ai2���o�e�JAZnಔ,�����Q�I���,(��E�%���g���g*?l0ύq\ �罠;��\cÙ>���vB���B�>v�ʮRA��i�`1��k�"��nh��p��1���[�0P�� o	e�xh}=�~�NsY�
�	��un�k�~�=�P6R�'�H7�oF��2�X"U����i�%���X�;t�	�[Y�	��	��&K�rd��ȳ�k�^��������U�u`Xw�z]w~N��N�{I���9��q�%xZ>���7ZP�������g����F -�A�R��5�/v1�ה��F_-��{q��#�A��O��f���~�8�d]a�AQ]IZ
�,�)Mý�ǖn`�9!�cpWZ!wC>U�ͳv��T�G�E�� �Ӄ�D.ۮ��dwҶ���˕��J��O��o,��.�>b�qﺕ΂�E�!❁�P��l�i�j?���>9c�to�:^��N��r�,2�� �r#*F�ɏ�pp?���Sb3�K|�N�|�8��֙��mVF��^���3�CzX��U!J�!��ua�&HH?�������p��R�r�v?���	�a��O��ⶢ���-�<)x"�M2v:�s��%v�'���bg����堟���\_�(�t��yI��&��`��P?���!a� ���M�*�/\���ĥ���\�|V�)z%M�i؟sD� �0HZ�Q��E5쿁.؛Vc�I��E���ʜ!�U�9
�c��X |l�!�p��9��� ������ԱW�q��`^P_Yɴ�L)e��V��A���5����_�yH4�fj?q"X�a6�
侼�WV�A�I���Yk�VF�s͟j"�����y�^:�hO
elk��r�!/���m6Bi�l��uB�
��r��{�(���� e=�7�G����x��-jѺ,��JoӲˏ���&��ap�e{�2`�V0��<��������0�)�

�/��f&� ��v?�,]����D�5�H��;��|$�l�� U-�ˮ�U,y�x���݄�Nu,J�e��^�?{�э�^K�Ĝ�߯�ًM��{�T�{�h��H��k5S��7��R+�I#9�W�$XLȥ��9�U���S~n90�À�l�@~ӵ=]�&l	�+�
���B֑�\0Î���a�w��� W�r�7Xg%(���0��S=�����|�~*{����&�_�I�Uސ�`X���B��G�N�l�'��[x����s�E�@ڑ�k
7��w r�tNZgM��F1T�+vݱͷ{�W4g� ��^7��6���g$�O5gi��k�|c���T�_T9&u9��w��D(W��"8-����3��x��t/m WJO,l9�u����Q*���%.��8MK��\0gMG5m��^�6�/�����Fk��Ё���nkcc�+/�V�#Um�<���D����pk�����`77�Jw}�u �q�Hx�1�3+���s9��S�̌����I�;��5�d<8^�x��>5�;,W[�q��#�lb#Q�^@岓zLkꍘB2�X{��p�����æ���E8I����r�ӉF�Py��j��5Ν��c�D=��$R�
Cҷ�
[�H0�Y��e���YHm/g�m59n����<�������[�=��k����A��~S�����#�n4�q��5�e �.��V�CRA����C<n�+�l�����*ˀlx%��w:�����m[�!l �}��ڙ��biZ�!�8��~�rڳ�W���@B!xf	9p!��~��BLJ�'����-�w;��4a�����@ҊC$�X���xc�)0�QY�����j. #�0�@�J`q��0p������(0fwچX�K�p�"_��3�at��=�����G"šv�HCT���Q�����Ȫgy�E#��V�o*����wB��/�(�?�pP�Br��zn{�������f���b)�� �75=.;!E:i�}Ş7: YP$j�:Q&. �����O���-��W #@˵�`A���6����O��VI�*A�,�,��C@C/eⱀ�I���ҜМU}�j�V
��u�6�=���n�*��(3�f�X�������k���߬aRr�����X���Y��ֳ,�"@~�)��$(Zd�z�����C�(����~e ��[%P ���<�(,�^�:��K�sV&{s���MU�Rvo�0��'[�
*m�:��5%�|w��ê���1�P��h��軋���~ԝ��.>��ќ����R;r��@)�9�"$R>a�\�P5��6�D ��m�-U���깈�G��J�L���\�	C����!h�A..�����]+��ߕ��S?|C�I%����W,��D��sm�p�����%}٣��#g):n:UU^^Q]]S�>ᴠ;���ұ�燐�D֌�҃OJv��T��	:ݚŜY���VԦL�g���E�W��)z}Ӿ?��Zl��_�dHh��"$Bp�R�8�>��S�?�&3�#�Z*���w�^�SלH;�.�C����͐h�q����6w�끆bd�&E���6N�q =��~��;��g1�j!V:��K0��WS�$1��Œ$���v}�p��q5m�7&���ڑ �~ĲH���7$��-򤗑�d����^��L�
n%���z����R�:��U�b|����ML<��`�k@`��\�1�������`��J%�����������3^���2�F�Q��G>9@�ҥ��.�Zâz��zg&S�*���O������-L��-��;�A�,8��WQ��
�WN�!�t!���������|�c�md��R�Jc�;OwOQ���1�5�ߠ�]4�Rĺ��ʙ�����h9��fD��+�@;�C��y\\�����]˿T�{j�] 5{J����H��������HA!�C^���^�|��f��xG�!_�%��NM�k]G�+����"ي_��2���xr3���9t����QĭIj;t����lhZ�V�i+�X<;��t�Qh���l��}?D���?;V1-k�$&�=^����di���U�OpA"���{�%�0��/���.��7b}��n��t ����A5eSg��ջ����-=V��H�c�=a2��[)����MS>��B���Nr��Y[Xh�$�[���9��x���*�y�}B .�%�-��]��r�/@A?�c�R�$z�X�C�ٳ�D2Hi�k�yV�oe
�|�ۛ6�dGq ���wK���R��5����ޔ�h�x�c\����_�hEKGp�r�s)=��?�f6W\�k����br�ZS��9��"��8�/uT��>9!t���I�&�cl���{�A�Ѹ�x	�n�ۙm�3﯒:c�3�����.��&M@7c~SO�)�ͫE-(:b�����H;�[�h>?��ߋ���,qx>��e�N�3X�U�DkZ��P�?>F�.I���WB���M ���-�fٻ�wݮp��kG������;p��}nڥ��QS8ר~�[�6j��P��g����Qq>n|������ߺ��a������������;D��]�ƠI�V?G������+P
KD,]��$|p8�^_�<L����w���E�T�3
���;FO(F�X_;�2���k��",�in�H(�=vհ@� �@���'l�M�ٔ�-�g�\+�|w��7��j�5-��w�~} *�h�p(��C��wd�
��]C
l�n�FS�UiI���v����J��R����X �������e��+��q��s�/�j�������(�}��d]�L���r�[�*&z����.}j����V���^�:,�ϳ��*�m�+� ���%.��j8�?���PՄ!&���M�����5#Ï�b͜C��hm/���ҥ���-�?��c'�v��#��$�?w.X�x|:�g�&tK߰�k4�,
�Z��^�l�e�kg�[�Eq�{�7�>ù��t�C
6{�9���݀>s�B'h���&�^L!G0�q�S�D�T��֖(��ؒNY^%=���Ktae'�g<p-�t�YoN�;"��H��n2��)ğ��=R$�J^IZ��[q'�P=~J/��q�o:��F,����
j�ÜheJ��
Vp���׸͵B����Z�nȃ�ֹxA�������4�&ſ����2�������u��SA��,�an��� ֔��$<T�r(?��8Dg^�Eb�u���g��W`A�\<I�>K�lȊvw��F� *b�D�o��Y�X�+��肐��m�̲��^�0']���b�q��dAya�'����{a�!�J����VG�?�8���f�����T����_��n�b��l���u ��;�~&
[�Å��/��%8D���/^+�
�z&�JusXV7�Wl{��@]r�0�Ջ��3Ɠ���C�T��}�Թ E�Ƶ=W�G��Y���fdC�Ǭ%�W����� ����7C���n4	Hj��_�i��&z?�P�Oy�����gh!t�??"̸;�6u�r-{���fv�
2FiP�92Τ,-;B�:m����Ѹ'�_m���~��J�P���	�O�(ޢ�6���{�B�qc/�47W������Fw��&�I�)��W�|���Ṱ)������zSZ�A���׼��d-�,�g2�a�Q$>0�f�ZP����8�ǋ��ǃǪcʚO��:$�����
~����JOD���yZ���\�vT:F#VQU|���_��X�t2�A�R�|�w_Lĳ?�ѡh�W�Fth���qZ�x�x������MJ��1��\�D�w�{�f5��hKO8��K�2g�%�O��c݇ܨ��=�n��XS�&��p���;��k���ثC;g�f��H�\$G���`&������L)(w�J�;�#��f�V��aSAJ���!�T��DF)4�<��UHn�z<װ�0���RȐsp9��(�Մut:�$DW���O�1G��7�]t���_��O��v��wȒ��p��z��8t�:"�����8�:�K6�v�-���8!H`�H���
X=NS����Zxo*�fY 9M���(9���6�[�ցt�Rs�������j��u`2bw�)l&�g�I�1����Wv�����bM���Q+E ����+�ˊ�1Gnw�rOYX�@���P�ۇ�4�>����˥�u�� �Ng��;�l�^�ը�vy(v.���=��S�R���Q��R��N�n�pZ��}6qo��<�_i������[���0� �|�]P��rY���dF�S�7V���~�G�4�*���Є
�$=WV���\�����t�~آ3{ �������d��{��bҧ���0U�ػ5����r�������Y��q�Z��E����N�G���:Fޮ�lib`��@%AHUD�q�����(����ɍ"'q�q��D��w���cd�K>��z�� 7�
��'{X�O�=���b�W�u>��s��y��ֻ�(��Q�$�w������ϻ���:�\����\��5U@��C�dXu�N*EtW�k��`����)el۵�+Bg2�2��b@K�j�ΖZB`+'��&��^�W�F=Xp'��9��t��>?*[�h�ˁ��b�%R�X���<���;�1���l�h��O��g���Ȗe��ş~��	OĬ;H��z��o_P_���$%L�(��i'�0+�t����#w�9DeH��X w¯�5����b�0Gd�5I�W�H��P]'oޙ��S�zP��quAV?T�#!SjW�d5�i�)�qQ/ԋk[��ܽ�Om�$g��	,'D+a36��8[��[�|D�����*�Z��N�.��}ps��z|V�`%���1��,l]�eJե�4��ܡ>��_��*���7���{+i�y� k�p5PP����c{>�Bz���o;�f���p�~�P.`u�&U%_@�n�D�=w�|�]1�[�>/\�=�_��h�C���!}����]�+il�6�n"�xj�����9 ˣ��{^����'G��*o�Ab��y�h�_�8��H)���FD���,�'{L+�j(뙝��3Yh̖�"���o`�ҭ�i�܋
�N8�mw�'U�E��?�+�ƕ~�+�94�kF燕�f���	����	c0N;5��:���$I]�P��x&�{��h�z=씅�x�=W  f"~���\�X�/'���`���t	FbP>	J5��\\�� �Ͽnгx����x��B��}�o�P�Ի���B�]0�s=Ţs�Y֬�:�|ۇ�7�J��!�z����'15��7V�2���w����K;FcX{��c�ė�wM�Q7>ۓ$���m\h�A�d���J�������f�#����2}����l���V6��.��<�{2վ��.4������$���r�?)y����&Ŏ�_���.����L��!߰][j�U\m�A��>���N`	���,7�1�:F�/����#����}ǟ��(���C[Jc�5)��K��d��'r�ٍ�
�(l|-�����J��E�AX��(�&�F�{�����ÒB�.l,5+��r��=��\�M�X��N�˺�-@������&=!�
�9�Q�_<ti5�O*��+���ĕ�@��tg��{�cl�	IG�e��{�����iĢYأ�i��  ��_��ER5;�_���(�q!^���J�����j��:��X�}�A�<q<���&�� 6��r��l
Cs��5��P��Jw�8C,UQ��� tA���ǌ���x]�p�����}�z���!ٰ�t�#<9L`.hk��F��ܛ�7�?�)��pQ{R�v��i���b|_�x�	t����{��m��R=�A��H�S�;�hxg$ȥ[1�x��\�5�����䲐Ԅ��d�K'`\2�R�A!Z�W�a�,��F��ha��%�긏����T������ޣ���*T 	26Y�j��7��Ae�ģ��K�t;�.�)W�k�UU15����u����T�=I.���ٟ��2�)L���O#;����ҡ�������@U<c�<d����z���ը(�{��<��4���^ ��Xw��oana=m�R��-�OU��y'�8K�8��s��}�h(N)f�&J�����Ѹ�͡�}Gf3D�jM�ܵ�!�n�
f�Q���^[LC�ڤ����v2j���Eɇ�y��3!� ҵ ���ݝ�Áy�Q��	�*�y9�8Ъ�����ꇋC��j�):��R�X��&O�o��B���h�@'��	�K_L� ]�4�Ϟ5֟q��{9=#�/�G�q� 	%0��`�K(�W�����Q�5=�g��O�f�,�:>ܰ���c�d)62� V7����#8f��PA�w�!0|;�fC�2.��t32�Po6���KwИ�:JrE�R�aRZ��.�N�����4 ��҂�y�?��3Bc;H���y�X5���V�zJ޺ }څ#�ť���Qp!�%�{Y��R�n���SzN�@��%U�F��+9���������4�W��ԓ�?���4h�<S�=�1����EF����'h^g��]�Y�)�e���E�(���ז��%ԫh�@"��?�)����h���;i]`�էs��û�Z��Y�_��X,���Q/��E{�ʥ}gkQ��p�K�Y�+aׇ��BcB��O�m$|������4�?LI�_�u�ur�8�+z�ٕ�2�GK4�ą]��7ٱ���C�;����S
�B�
���,�,L(m�2{��K��h�_z����+��
�~�H��=�֠'m٦��d@9�
T}�P{�:
�kq#� �Sd睔�b��J�s 8I��RL���]��#do���d�jI)�L��|�}q	A!�͂�����`<���&>�-���R�`��I�<�>i�Q��}��?5����˅0����>)f��A�!�2~�ըKn�v]�`�²�u���<-���J���\�>1\u��ʷ�g`��-�2�Kp����ɡ��/�1(m�u�*�y�Q��ɥ��#0K8J��(7zpU�.;�ʅ���^�,��Pj(G7�G<ĭ9$4'o��q]�/�6j�;��P/�z�c�%�Η�q�;6��JDg�?o̿Z)�>ȡ��H"�y6�eP�r&�H���f��y����0�n'���8��܁�}FA)6{ye1=v�i\������n�u3���n,�39�ɰ��}2��IDwǲ�,|�{'�$�.� o-XQ?�L��[��y{@E���{��y�Yx	M��4+g�Uq���,��1�����?P��RX�}�MY~����}=����">`��z�z�/G�g.ytп����><���}�-ف	�7w����������~鍊�_�Ʀ�*��g��#��@�
b�F�a���D��j�]�LR�|uY%�H.�,Q�����z��߀�ǺA�mRΙ�8����ރ�,"��ei�2��n�����0L�gT�dP]�
���4�\�$H��g��L`s
1s@"�;
�B����iY���s�K��j��K�b`CyP�?��yv(����`�i������M��U���Ve9L�F�.0�
i3�]T$��%��t:���B6x��G��+uhޗ���E��K��x�6�w����.5H�e�/��{��!p!w!��",c	Z|B��6��5�uB�#�Åz�Ec+=j������6߻i+�u�����*�b��t��u�Nņ{�>wm��sx̇F�yU;'�G9��>����T�թ��$����q�H3/ʧ������?�8r�c�o���C-% 	����m�߼ΘD �aE���Q�- �?'H���%+]��H�ݙ˛|Adϳ��$y�E�KU%i'u�Jm�O`��j�(���x�Y�}�P`|�?�~�Z����z#� tW�A��[[�E~���g)��4�w��*[���,�� ?�6P*���)���Q~�|��ӇH>�D����V�*Ou0�@!�5��F p��/_���䯥5���F��M�X4��piY�,�����8�����\Z��n��TI��@+�ʃ�Y��@�_�G��L3����k�s__��(�a�z��~	�`��7V������j�����)���Ѕ�����V�r�0����8,6��At��+���-@�d��u���DO
�������hP����?fP�i���g�֙ۉ-���J	�υh�\q*�Kw����y= k{H�7��ɚt[Y!��pc0h|@@�_ݛ��G@���'�;�q�K��L@m��/�/Pv?T';ݹ�tǢ�{����G�`."kN�Ӂ��V+7�ڑ�6�Z��O{mUNyVjP�3�ߔfJf�B���F�^ ��W;A��0g�wk��x�}���0fsv���C�\�Q�����1=lW��>�U��(Rv:u��ݘB���Xڏ>&�0���DZy��7;ɾ�)����r&mDŭ�G��M��Wt��F��I@�鵁������� �����E�O2L�C�P�m`�D��/%�p&u��a�	W���P]�Pr3 �9�	rTG��ug:�q�hF�f�E~�~� и+�ڙX�h��ޔ?�ْ����r񉎧�IY��TaD���/�9& ���䩟�AZ�����B��VG����cKF�xp�顁;B� kjn�
a�
[ޠ�� @z��>t.�V�;Pף`�79_�.�JB��`PGQ�<(�������O�|����,3d���5�/��N6�X�VD����s���˽y���<[�?9�,5��U%�bt$�L󋮋�F�A���������D���W�9o�<��ŝ���R��,ߐ`fq^MztK L�H�Jݛd�S�]�)Ft�����������;Z���~z ��oq��|~7�ъ�����?��1��$���̏:�����Eԫ�|]�yW� |r
7�َ[x6C��vyVF���{�t�%��s��<F��C��aZ҇�h���P�OGGW&A	��w.�S��X�4�I��J,H�8 �`��2���á��_�	O�b�e|Qk��)q�CYQ�_t�����X(>��U��6Z��ސ{�ŉPF[�����`pݩi��ϟ�r�m�?���p�Z{Z.!�C��6�ė��sK�Jq`D$��z_�I��ݰ2�]|�T#r]ρ8U��� ��=����\.L����"�.��t��˃~�WigT�A�����P*��Tt�p�U�-@Q��rp{�_@�d�򄾟"�a7���*�7k@�dy�*��i&�kS��FؓN�aΏg �
��g��+��M,�9Etq���I<��Ӊޘ[ьi�O�to�|K��{�N����+��aeEk����j��yQ�#�?$�(Dhy)�*���:%<1*�r;�����h-Q�����Fv����v�����N��A�Na�{ԕ��AJ��B�HGN�}��4T�k=TZ<����7�z��it��S=1�N� lh�ݖ�.��S������!ƑPS@F��l�6��G�#��G�����R��G�E�� ��$a����Z%*P���o�G�6N�����0`�۶�O֏>������7|1�œO��{ӝP,�}#Տ̶�f5i�9������7~�]
��Ӯs,l�/#PE�'Й{h��JW�3�=+�l�%���4��^ݰ�_\�rxx+��s���k�)��B��jq�{9!q`���ۨ? �p��ɴq��o�I`+f��l�5���ҨU]qn̉��;�4����s��n#�d#y�yh�%h?�S[������B*
:�xjAZ�u�Ӻ
7%k�9S-��Ғ_ ����GO6NP,*S�������\���KCcͱ�Ih+
 ;��X�3�ߤp���C�n�Lj�X+d��ݫ]��L��_���&���2�P�H��3���4
/]�������D�I��:�����ҳ=_�O��*��yB��7�FW.��b�J�M���B`n.�B�o/��cF���L��9�3<6'�$@��h�'���lZR�z������0B�aFR���l��1>�*I��:gy-��o����ODj"$�1��)�=1�Jq��m�^n Sq���'���ґ�N�&	%f(�[b�|0F��5�*yt�uJB�n�����u�K�r�6:\� �`(��c����l}h0g�����5iU_�g'�g����/~��nʕ� �a�
(�GRˡ*@�ڜ����t�s2�d�'��[
Juuv�Yi0T;>y-F��8�L�'
��W���X��̻�����%tv�N%��?B����F��:nP�ы˲�~�+
).��H\�]A8`:�7Xˊ�eԣO�OdՏ�i��T�����z�HF���J[���`����'�q�O��X'�Fc�
E2ɽ�-�q�B���j�`���s�cj�p�̴�I�)g{��X�����x'f�ۗ���"2H�9A�Զ�������O�h�{F�Q�a�@;�ysoz��[���.�b���'�>�G��:5<9�ۮ���S/���Kj��T��T��m _\�b;�VW?F�Oy\A�M���F��#2Z��J8�o��[x�(����^{�����I��J�xmM��c����W�xDz��=氺-6����mq\����]���G��9Y�͢ # �M-jc�K�)�6F���F���昲ͼDs*�ٚ/�p`_�� �������*P��i�x��R7�	���sxUPr�H�U���)�����rx�H̊\���^�D�Z�'�ȉ@���۬�z��l�/i�
w�蚞j9y�v����u�|��������fL��	R�D���(�TKP!F�`��u^�O�a�*T/���yجNA�v*Ǌ����%,�ϒ�?垗��J&v�b1x�6��l��]q(P;�P)'�����Z�����̧�c��~6�e=��/���
k���!���,�N�M<VB3�⒩r�V��C�l,�C����*�/fέ�b���ªr�j	y���,OF[�s%�J|�3��^�4A�*FS��&��h����2� �E;<�;���c�nQv�З��u����)��Ǭz<�����
�Eƀ��v�,l����z��&��?�=��R#�A�g��4?jh|` 36<i6fh?]TlQU���ʠ0�B*I��5A����;G��?��L�c2%��Y8��ps�6�� B.s��ku��4(�1�T��tHb[:�|������d�c4U�U�juo� W��,h@[�f'�zz1vZRTr�E�"7�%�vw�{���9F��/W��d	Z���`ծ>�E)5n�F����N�âv�p�1Əb�/�GB�&c�#ـv�t�Ȑ|AF[v�3��յf�ӟ���5 �� �E�h�e��&�h���}����zqg���H�N�H g�������������]f3å���;��B���e��"�������qr8Ʌ�aS�h�|��³&Q�oB8u0��h���Iվ��?�K���UTg�  ���� ?�w�}����ӏ/ ��m0/@t�`<c�H��h�3%H�}L�8�3�%qѩ�N`�eM<��0 �Ec,������T���hgm.l����� �V��ATO�x�I��rJD�%O�zQ=���2� ъ8M�Ƌ��`�Є���A�P��UH�(��;p/��n�x�-e'	J�Hg�c�5M���,X�1#kģ�(��%ش�|���6D����,�}���������a�~�L�җ��h��u�>����Ew�1_>�i�,}���`�nE�[��AU���x�젨k|���W�G���;���8���*;��|F_���bv/g����2_e�߆q����Y0�`���St��R�u�'����?5&:oL;12�������q�Jł���@�����}�@�6"�D^��p=��� ��Jd��A���
Ϡ%���h�祉*%�y��t�[4ɻ����	�Gtε��j`��sň,DI �o3#m����[�N9�o��c��LE�)C�*Kp~�#�/����D�X/�!S��Dԃ���:�ð����^*%�p���;O|tN�K`� /�|]cpS�z��s��O�����n f�7 Z�t�o�ӄ
�@̈́��!#�d��0f�2�$0 7Od>O_�&��������i�D���v�#&W�8������Sʭ?P��*�mY�9�e�ۓ������w��%f���h�����m����3O)}�#y��k�$}��ɮmk�[��y�h����N���׽[m��)EUf��F�#'�ȊIg����󁓴�b/�����|^��Ma�
+�t����6�ϼ}�W� +�C�8^ŀ+~��O�TSsȨ����m��R�^G5Ŭ�@�=�;eܱ�&W!�}���"������K��҅��Vt)��D�x������(,��G�t:#���5K���0�\DS�D�5�M���C=ʌ�v-ws�8��d���w�QN:2�Ҥ>B�����:�������?Y,B��W�fEp:G�}<��z��+h/�"@��u#���8 Ɣ�&t0mmrݴ~�K���q��W!7q9�I�K=���U�c��%'�p=k�!F*��TKI�e��_;��ճ�W.�
?�;ΐ�c�i@�$��W�AȐ�;Q�|9��ٲ��'�X�)5��~�����w
�7�y���V1�n�H+�4�~�[3�T���҈p�А���cU>P~��حP���3��E�҇,�s���[�*B�1
q1F���K/�i�bu	�7���qP(/��E���!\���dΞ�e���1�����1����W#0�v��y"�C�s|_��n-,x���aR��QT�q��z�u��K|K�8���HOԆ-�����^�[p��X���p�t"|�Dɵ�X��`���ҭ�^jg��8</���.�d��c�f�Q��=B�2_ھ��8��d���G�%Z��S�W�6�:�4�Z��H�lѠ��I�Jg���)���-(��5x��ۧ~�A:�U�a��H��8r���y����5w#
aȁt���x���I�qߒ��[�Ѭ(	����[��*
k誊Ro���Dz׋$�;�LA�ۧd�qJ��m|\�f�ܧXI��h^p�%�ە�Rlb�����ېafl����������dU_iU�2Y,l�4=b5��	�P����|��\s(���l5�3a.%�>:q�s�8o� �ɩ~�M��N���l���Z�!�#���zQ@Λlν�m�v�֣� ���i�<�&G`MQM�!u���"H+�x�6~sV�rv�Sz�7�dq����5q��K�:} Ɠ�`��o��5�>࿜�}�I l�<z��d�Ev��~
�P�7a��H6���$8o{V����mA�hB��C��Y@B)�ml^�Z�Rp�����V),�Є�;����=��}<	=���n�8�E���q�3R�#k6�J�Ö+P$2MU�"��X��c��6vD�J�*3JD�ô��4SkΕ^k
^�
_�ǡtm� �L�寉ے�b�K�����$�>�@E�~]��:�$� r�Vũ��$E->�h���㠆v:��=��{�ݤ��,�����1�_5��3i��մG �W�{�Cy�/F$0�$ 7��	Z�C �zK�$|��e��`�L>f�i_��~��z�t�Ky):;b�)}��T���<-��]Ŋ�j�ds6�`��]0�<v�I�E�e�&D���� ':���L\��AWXHT���Y�*�ͮ�+�!�&_.SQ�W�l<nA1��XB�p,�����'�����V��.��BͲl���Ӫ�q�{RJ�W�`
_�Y�O�UyQ���u�oe�
��L��nu��������3��'.?n��]�z��|�v� .釲�'LڄF?j���Q����B|���Yಖg��_I�do[tV^���p����'͈x�}0 gl��a�s�� �d�����	s�I~?�U�:��>��J^"0�Gs�-B���t�ˎ�̬[azT����̜����B*��L��S�t�4�����M����xʡ2��R��Ay��k-�E:n�U��s��$ʜ�����8ѓ��kL�j�6� h���v9ם]��=%i�z5̴�b�>����Gt�$B���<f;v(��P��zdg��J"��ޠN�N~�.��M�R0��z�����|m�1�Ui���%����1�,����V�"�<���h��u��w��p٠�P�.uA�;O����;���UT^u�i١$����ly}CXVL��<n�����F"��邀��$���q�)X D�j�z��@�h�g��A�~���1�̀���&l1h�ÁK���}R_4��.�W�>N�6sp.�d�nĢ¯_��9d�Ͻ0�d��e�pC*���P�dO���i)^�4�A��>s�&�o����;*�<��ˇ>�'�� 
�;��+��̓�ԓ��⤖���)��Um	 ��K�E}�C
����� E����!��z�>!ʭ��9k�-֍f�(;u�F�6N�җ��A� �6�����7�N�(I����E��ð��q`��lx��^��+Y��L i���f\Q��R�ܫ'}�O�ˤ�NJ�t�.�l'�@	��Փ�ˤ�� �2�h��2t��l��"80qu�'`����2J�,�$����e�V��j嚿��zU�R� o���M5Aj}I�\�Q�<;���6@��r�t���s9~rm��NR�l���J�r�x`��r�p�d�	�۸~�pl��Z�� z�Y ���*[U'cl(z�q�_��5��9~����w�b���_��+��Ӈ���B��M��B�ƉYhL1�c]��Ԇ��0G���=N�#c-[���P���d5���ϵN�1Q��kN����	oK���t|�
�e���́��&�Q8��}����=̶:u��|�^ajF��w��E׿?�v���	�|��ְ����:�Y�ɲ����r.�>趄M�χ��b؅��E�u�t�4�&�I�����}����Z���w�wj
YD$�z4'C��^s���,�#���h75f��a�p���E򷽻�g�c;v�q��<��Ѵ��5���lZ�r5�$L�O��-��z""w�2����r_���L��Dn���_�$��<�p���;�ТOډ�C��~.�P��щU����
E~��9n@��~��έр�,�+�H�&��V�|
r��@�?U�l�]�n4o�P�V_}�B�̛]��_�^ݫ�ۡ?�k�m]6�@ߜ������ě��yv�?g�T�(z��e�y�DWQ���H^I	l�[�k����j�&�{5}c�\N�k�R�2��&Tl5�� TҀĢ�j��
O@��f�P;���c�S��6��y�e:!���9Q��t��>KDܙ�0O��.��1���_�㭣���gza�=�ϣpÍ?�=��b���Zp��n�E.���$_r*���?j���|�F̫�h��S쑧k��|u���y�~J|�ד�d�&HM��bg� �L��&�-�2ڪT�� o�֢���n��U�1�[�İ3���C`�y��%��sX��D`�w�F���lJ��~b�l
��
V�>��E��|'��d7�CB��L��Ln)`�s�l'�Zo����Z'P�Bh�Ǘ:S�@��W+�@N��6��	�H���}R��u��ݘ�H�{��H���\1B�,��x(�c���8
%��h��v�'���+-+�r�e�����2��9oN�����9�"��,R7��sZ�������7��{'��ja1��X�e�4�M�ι;�2��T �������n��S�	F�1��{��}%�h+�ؐ�@���E�B��0l$5�J��{.�w[р�����u��.���z�o�ǆ!������>�a`��z%m��0�~;1䄓���
���s��K�
�E�^։|����1�˛�y�,�� ��"��\�v�i�������ϭ��9<^� xS�#���/��p���^�	�8�_���x�[�����t��/�D���+r>��Q�Y!��V����	Ni"�A!b�.�2PѨ�L?�k+�����Y��?\��_4�P�+Q���e�H�k*b�M,�[ZW����`�/C/�7[�Cؾkd�<�Z��s��C����Pi��.�i"c:Ds{~���kg4[	��_
����t�V��j2lu�a0�I3g��Ѭ�c��I8�`��3룟�@���/�/[WT��`@�2b
S$�
��?��O����O�FɅ�~�6-%�n �Б������ʴ��{�$џJUm�i#�-��nX���(R�~��`Nј����A���%��%�jR:؃��9#]��t�0:��e���䄢�Gք�bWAi"�I����Ms�0�D�q|��c���%�҅��ïQv9�v�:�d���C��*'��o�Rp�FVU��^�<<�m���P�E��6�t]�x��{��C׹]-�
����s�E��s�����Ks�z���n����Z�)m����(� ^�:�}d:B u�|@S�r�#حAeҤ|��� ���e�����`���U���$�:���ގ����{~����U��N���,�����
�./ `�M-�(4O�$Ő���p�|Kz�U �����&�е����Q�72.Kqo���������o3���C��QԀ��VO�Q��G�����̙�7�}���6r�����Z��\Y1ubrs"�V�`�/#��	�;����y�g��*PM����Ut��4PyB�@.
f�^�$�/2gc��}��H{^�w�����~���m�<� 9����?�'(\����F�В�643�'X��XP��w�EY��{�;m�K}S҂�!���*�I���NW�Q�?^���5%z-���R[����c��$�"�D~���z����g&�]H}��!O�je>u=c�Y���u/]�W�!���%t
�R:�ٜm�lW�n}������h�7����c��������Ѩ������s]!�EP��qY���^m��p�.]�o�ZŖD�ԼOǩ@'$�UyS�I��Uk���H}A�%�$�޳7 L�o
�
�Q���n�5U�q>�������_
��������I3���oC�S�a��[pv��Ҥ=Sak����:tّ�Ô#p���0�}�bC�����.|g��M�5ߐ����j�^%ܡќ#�H~Y<*�Z�K�Dp(�Ac���Ϗ2��ͤpu�֚�l��������ai	������<m��h/����;��4>���n/U[}��'D(B�<�9����6>�t�^@�=d����-����hg (���!��7��o��K�����m|����ޔ/A��%0��Y �
�uT���~R8A�C �w�և+M�ת����]9�F8�=Ҙ�����夵�{���6?��3�l��-:{�S�
���3Ն�ih���dϧC}�<��MH9N�Άc�`c�&�>����T}l*Z(+xhr4h��P��w�G��&q�Kҏ��@o9���=�o(�͵hy	�ߒ���8Q�?2��)RK@�ePp�Ľ��>�S~��%�=C��*q�	�k���!JU&A���h2�MZ�%EY��w�ə�Ķ�����s�2�À����D6��b�y�t�I���� �;s�d�^�'�k�Q=/ɧ�P��1��%��&���ۜ��S��v/�=g[�9�A�~�w�r�EY�0}68mJ�/цnf��Y��ػ�1G�3so��@��1�D�'�G���~Z8��!��m?�c�N��-PH�E�kg��e��n~��<���Xv�akmWޭ[P	��@l������6!bQ�n���|�T�@>=��^�ʅ��v��B�O�A�b��Dj�CV�P��o�qOI �|�c�m�๹l���au�^8O�n��&��$DRB��P+%���Tv�{	��D���Aj�:�G��m~8ϥ�5��������_+�s�wn1=��i;,%}�u����-�/��@H�dA%�t3����qv�-�7��*-Y���j�F*6a|���EfD���Z�ƧdӕD
�b����Ġ��!����Jr
Q�J���PS#QM�~~�궂��S�s01��<�R��D'1Z�+"<֯Or'�W�U]����K ��S�(h-nW�[4b�}
N5[0u��!y��ٴ�!eyqN$R9��oE"���}�@f�j��<�iI�d�1�ײ��F����O۰�&-oV,��u+��x�frfω�At(�K������1���L�p�����)?�����(�RdqPDU<�e�&����]0���kC,�ľ�z��R,�t�K�������d�D� [��Z��d���;�m��%1�i���GK�=��ڪ �}��d�*?E��ȵQ�
����K���)���B���<�����'��������|����Y�T�Ìn�Rc�C��u��y���4�^��y��X���D�̕T-�%���%��6�.6��1���6_���1@l͐N��i@���>,�:ե�42�[7�Udm��J�3����t�hz���̞;�8��s�.W�jF^Q-�+O�KQ
(�w"��\i�B���U�3Š7yn
,B�(�T��x���`n��j�M@��ߞ�
��|G%E� dT��m�q(>i���.����a1��D��:Nq�Z��T}�ͳ익�r,��]���_�dn��gM�����E���[|߶p���~�A�Pc���U�y�r�eRR���{s���ҽ�M�B�H��cW)RV.�|9��[����.�7,�:�q����ܰ���]d�8���� ������[������D8Pw��.��p\O�E�#L��S�[�K�<\�QڦZR�"9>v��7	���ED��n��%�����;���2<?�[�����ml�+^G@���m'����R�,��-�W��'��17\�=����.o�b+vc����L�Bܚ(b�b���}��gkY)��g��W�pH�4���-�
�%ҕQI/����f&�wQ0���>��t�C$A���r�9x��Q�۬Íe=������U2���3�B�U��[�g�l��:٠�`�5s_�[�s�8���Fe�ֽ�ܛ����l7��Ӫ%S��
��-������/�~�:ig��*��k���qtF��1wGۧ��� F�M���ፈ�b�+E|�ِ�Tl	ȧ7��h��ŉ��0�?����Z��o����
�삨�gQ�Gfo�+{ǭx� ��.�Ǫ�wL�8E�,�1�D�B�*���)�p�JY�g�=�rGD�t�6a�_���>J�����&�q6Ey�2gk�� ?)��
y�����b%$�"�y�i�	��N-l�����H�!L��2� b���37z����V��M?�ኞJ�m����]�9lr@KS�皗ҥ��% ��r�&w
�,��
ۚ��'&٘�%��k�m;.�ĿQnt��(��~����^-Q�@��r�5'S^ײH��&c��d�^�y�6T
��4|��ڵLx¡mI%�+k�A#dg R!��k�Lz0K���� �Ѣvi���F-x�S`L�⚆��F�)�!5�SQ�X��[̘�mm% �<��*^q����4��c;�HHh[/�����f�����.�t�A�.̲�T�=�HDI}���Օ)�|�-ua,����j�X{�L�5���5�/�u2��i���o�´��X����v����iq�@�xvβ���j�<>�A�|��y�T��� 4y�Gv��CE��q=�"��~�s��Km�[U
���բ- B1��.+p	Z=�Z|�ǕZ�hx�^y�/���F�L!�w��JW�����3���fvN����
[n:�u���Oz�-��P%��+�m�o�"Z�2���z�����sl���j�yuik�km�ٝ!-xۙ�>��_5�t\�p�o�ƎT�f��+��Go��G��T��Ƒ��'�~7@N'W��p�b��8t���� �ݒ
��_2�1��`Y��k�O�G1Fq*P��V��D5Jb�����V�.�"�Vħ|�\��l �>�U`�{e�c�@Zc�H���Q-��ڗ��0X��="-�I��عP�XEㅍ7���aZP]SV��)	^�)��'Ѱ��7�8l�,:�RO'�򷳙-�w��/�P�=�p�£�@xi����� ����?��I����CN��l�V�� �RKX�W�/�B���MW��������RE177�o9?�Q�$��f$t^�����C}*0����I�U�gNzw�Z�GZP./�rc�;�#[w�9e]�� �gc�J����u�q�Dl�$�~��4g�����$����$o�EO.:
��yD"Q�i�ň�[l����WA� Rhs��*٢���Q����X�#�8��z�g�~7�k��d8u�9�}�W�>�Τ�,p�������rX舱�[����B��@�>vY-m�|�r8��b���{!ѓKTAK�R�G��`-�5�e������>�v�V'�c!W�cHPz,���B���7�_oBϽTA>�IM)tcm����K��ơ�M���)�	�밨�g��@m^����2┼��߇�[����i���xM�sUg�j%������JmD�E�,��V�3����~
��ڷ`=V���}`3<���B�ݜ���xLZ1d}�R��|�
�۹��j�͉��[�d[��S�̊#FA�Q ,W7��.֙��z�ȥ��B'��^i���R�T
7~e&q�{\��Y�y�_<�_a��Jr�V}��V�Yr���5P�Ou����7���
ٯ7mJ�l�@&Sk!����h:�!�����{���z�b�ci���X����.�}�b��B/����
��qX��ޘ��@���T0�) �A��M � J����Nr�ARr]T*f���/qZ��`E2���g�Y�Y��dX8�gN35�N����R���F�)�|39�{)��y��L�1������E>�^p5�%'=>��0&m]��͖��״�Ny'.:����/A<� :�x��ݓ����
����P���ٷ���5�Q�ݛ�X�c�a�c�ϟ���k��jH���b 4�]&�^dB�Ƕ�*��/��.���k��궻�� ��˗n���ԂH�f�.	�?��z}��KN����7NGxg�>]�"^�8�~t]�>s� 3�4E(�[�D�$m��������(l���˚��!�w�1�Q�/�2��]C��=o{y$87�-�Ro�����ˆ�ԉ`�T	��j��4m��P��o\�y4�ۭ:]pk�nE�!FX�c��}(ךe�P4�˰�N�	DD��/�V'�N#��5�A�Z�?f�҇|=��3;^�����*����Je�m�בɸR̺HX]
%�1�EM&��Ųm�\&�t�l�(֩�u��K	��.L��Y&��TG��˩6�ɭ�p[���[��Gmr�����Y�`��D�x;�66��54q#�F����1
-?rA�i�V��V��v�@�+h����qs�,
"�;�ha�Ur��_&:���g�r���A�g?E4D3�{��iN�B�'�!0��<�����{<˪?���Ac����V�7[�o͊���7w���#S�'�����[�P\Pi���t��� O}a����*Q���&P����Y:�����!�{����Ve�x��	T�l�N�/�#jK�^�0~�ÈM�]�N
���[�XQIžJ4\�z����B�PքK>��Wl�M���'6�����Wk](�v+������0O��ʓ׼�؁(<�X�#h��al�?��Ʌ��1��^s�m��蜫"W�*�
g�Pj��D˒�j��Bd] 44���>��K.<F���F�3�n��=�����T&*��j��$�x�����j|�
���g���z�$T ��+e�`k�"k���͟k/�Ɲ���m��u�9n叞��7�9y���i���ۛ"�6'���J��H��f�)o��3)ݮ�OL:���i���k|��>&&�J��rᄼ�g�>#��3 �T�O�E�)Cڟ�{o[g4p��H7�`�?�X:��"5)��Y"ԯ��(���?Kp�{_�� �~���<x'�L�F�,�V6n�ԏI�ӱ���M8
%�o�,\��v"© ��	f��N������0�������� Ġ�C�E�)�$���7l6]3[4�L�e�-�Q�!�����7���57!����������|��ė�����V�*Y���&Z��7����&|��~Jl:r�st)��5D��X�S��
=�UڽF�0H�m^p���&�Mf�^`��d܂�1�v��WeO�z�D
�Y��X����[��\��ׇ�o�:
�Y�yQ3ۡ��{"5�U^%\+��߇ ��dH��B�|�Q�g�v�'�ey�D̹)^��|x{Y�m��w\�5GD݄��kQ�U?K���&��wk���v/����1�h}xE�Qd' ����o�En�����7�]�I�}N�ь�)�X(�Yv�B�p���.
*��5;4�{nZm�,�d�������JG�c�3�<�9�A�-��c6(��j�������ʪc�8���w��4��Xu)ǻ�P��NG�;�Y�Y~�t���tV�6�����0�in�p�o���ъ$�BR�?�~F�@V�r�«��O*��Gn�;�<�\!W��v�	̛�9�7���6� ��0����Uuq��A|8p�H�u�.�3̡]��P ➭v��sIBo��hZ
3�4C��DߔYPj	y|\�ӱ���x������1_�`�M�����Oϓ)SEa���)	En�O4L_���=����,E�I�~�y�}�;�I�1�d�$�qI@����o쵀X/�?eq�@Y�Xk�@S��¢��$������ ��Z��03��h����Q��,R�.z2Hv����}|�^Dk���~ܰ/�r�;/�� ��hB�Ǒ%����5W��$�5<<�|^?�I�[Re)�����h�Pi��(82	��u	I[4�'��f��xl/�&z�v��ߟ[�c�V���;A�)5���d@�%�4���ȗ�� "�賿�'�g��\R�Yq�8�#�#�Ǳ��������C)*�5��<ʀ7�㛖�/h�tuE�Si��j�޹]kj�(8��BH�	��G�eE���i{<��)!,���Q��@$��xr��
��(>u� �����r}�*�z��#��ow��9��s��ڭ[�/x�667k�լq@ˏDG���ï^�9��I8?�\#	e�CU���O�"�AC� ��'���������e�GҐmtOqTa�R�x��0dpw��/>�>�k��lx�y(�Jc�YX�9@	|a�8)���1YA%�P�J[�ޒ�Y֠鸠@�J�=]�d#�Gd>�9`��DH�{�7-��r��7;Z�7xr�3S�܌U�q:��3O���A(ŵ:���h��p|'��@�0�q��"���1�h���S�A�8��"tpVz{z�Q Z�ӻ��`�f�#��!�J1ʃ������ȔOIH����o���W��֥F�xaQ�s��n������3����s�p�ȰV���7_|���I��t7ӯyt;&f} �����u	L[	�6�`j����/�Ȝ�ī��K��+��rDa�ͻ��W�x�"ru#}���L�p�Ѵ 9*k���6��e�@����Vo|�³[�1�Oͺ����L@���r� �9���U@7����S{��j�6<��`���[7}�ީU8
�>f�H��ҿ"b�y�vUOUhO
�������6fm�P`Jԕ�n�d�L���'L�N���&d��kh�P�6(OGݏF�5��;Y��g�-Gݶc��{q�1����.,��2�×g�Ķ�C{��d�d�O��V���A�4��Ͷ������i��;"��c��샇���Jj�=���qF�%5��Pb.���P?�m�X�k�n��Z�A�h�)��!p8��wPsv\`Ma���B_c�ݳ|�Y��7*Jf��'�ܹ�h츩������ 
�`�//b^!S���\֌j�+��E���-_ƩM؊(��n�i�J*6Փ���w�0��#�Eo���'�:�f40MbOkv�`{X��:)������Q+�D-\����!��K�(s�ʗh���e;yBZ~5ި�o?�E�u�|��3��b��`��鹜�J�t�z
hH�M!�(L�}�,-�|.�d٧���*C�U��S>k/�8�5-*��y���D��b{[���[te��%\G�0	IC�V����cl<�;�Ƒ[Jɕ�Xw߃�Ig�XUǎg�t�i v��l�U�q2�)�|j#{��;�י��O�'�(��\2%8A� Z�_�NsZ�t�n'�#�5�f�U�L�sz�"֤a\q8�L(H $����#���S�ƽ�6�e�z���9�YE��hme�ɝ�+��3�5��3	���}'[7�8�<� ��*ad3��X�S*���`��j����.m�Jb�B薚t&��WI�E{IgK��.�q�H�m��$fg�bG�<�����FY,";��x_b�P�ܠd�"Aw�d3$�.��4�xI;M�9-`3>�A)�
�0 ˑXS�qQ /�x�"+Ck�,G��,�j멜Tړ\�+"�<<D��6�4�ǩ�|k����ӊ2O-��wR���(�P����hz����W[��tXp�Kv�G�;�r9�Q�A�g6Ji�B<>���tU�փ���.�#=j������rx��{��jY�n��CDA�r��O����W�|�V�y֢m���q���`�T܅��;�ک�3��=�O�>�xM᝻�P�HS��i5�0'��ט��Ќ$����I��~���=�[0�G>���[��r%A��nao�0,8���ӌ����m�)�{�<xY~Qk��CX���0�o�ۜ.��Z� |%<��2)��os1W��Q��O�q�{zr���ф��(C%߬��ì v�t��������`a�2c��K�gl��S_�����ުK�.oIdq'aFi���oJf,�m���e��̏�7A�b�}����t��WEW�oo�	ؚI�g����@DǕ�T���'�����k�L� �I=����%`�$�3�W�*����.�ς�붿���	8��$Iߩ,�5V�aىD�[�ż~���h_�7ޔ.�Ht���g���J6�9��oO%��иx,��r>
��5�����>�G�y�s�
t&�(#�Yv��h닊r�㨟1�1i�Z3-]cš�iA������aB���=%��F8��VK�Ϡ�W�1�g�(c񄈁�3�;�+��{�ɎH�ܩ,a�X(HN�p���4߁P�Q�$zAյ?�KF8�B�����b��ؗ�I�E�x%wC|���[�a#��RQ'jI���YZ#]~z�@N&�%5^�z��!�%~,�0�lpJ��u��xɣ;glF�pc�5����Ae���u�"D<� ���FN�i�R|��W3<�a�*!�/t��HĪl,�<�.���S8�Q�f5�=	�
k��	���\*�� C��zvQ�f��z�غ:V0�AL��X�BF}�g ]�n"e��ѡv�kB��XeJ��2�{�;;���m�U��Gd�^t��l�K�hZ���U� ��P�lD
bd�	���P���J��WX)������a�z�$�Jdݕ]>�butl��J��7K��u:��\DV�P�w�j�[-y.��S>�u�l�I��b%��K>��+l{�V����od�Ҩ���gW�
�w'�bcS�<�蘮�w��.|L�$'��U񄚶�2������ HD?�~��k�̻����t��g+G��rly�.�`;�A�i���������8Dx�S#+�ܙ>k�M���s/��te����e�-���/<겟7���2�����v"���tse!L�D�מ�T��J��t��{�$"hf�W}_�8�ן��j�d&�铦|E|UF(��)� ��k��DHV������`�7j�u63��2Gqr6}��[%��!�:	���	�%�r�.�a���@�%���'fV�x;�6�֘�2� ,J`���5��ܯ-�J˼���Ƅ��z&X��W����ڹ#��t|��]v}DAᆈ�!`����l�`|bv�3ݖ](ZE�B�dY7ػ���^M�&���fL��H9��YϞ�t�J�n ���_�\'�+2��ŗ�l��6�� u�Fu�T���)��ð8p_���8���?{zw)��-��V����'/�ds�Z@1p�̇�%���1&����~�NE$����+@M�� ����s��cAǙ$���i�$Q�JO�s7���ИM���;g�Xw��SO�Pmb��#y0X{p �A,�=?��$��;�I��U��M�b��-=3��w�Ҵ��F����=�t��)�{ިo��cf�ٽBx�U����:��B[�ľ�J5w��.�˳��5\Se	m'eǪ~��?�(L�f�5{y��+jSd�8Ɇ�����K7�����|��R�y��*?W��`p�>�*�������{�u�ڪg�"OΧ5�����ۈx�v��8\�������%x�=� +Ah{��f"�X��`�(�"l��+)I�@# �d3�ŘGR�54���O����NH��98�1�>��֥X ����p�O0@�?Ϫ����gu^lȡ�������8�v�"[����<w-T�� -�C��d>��+�K ������c8+�}zb����jβBc���,�|�Н[��3����g�`o�&�o�f?����@Fp���ۙQ��Pff3l��p�P���U8���<���/�0�����Ca��~i
�_b�����JZ��;q�'�?��N�+���w6�=�Z���^������eM�9L�<3 y�ۄ���K�5������PoW��p����<ju�+�0p�ΰա'���:�j_x�bh7�
93�-�,6���<�{ot	{��U����6bf�ȏX!M��ꋫcశI�#u߬���K�!^�9�o��iƞ^�f��ˀD.J+	+Z8"O�<k��Q�[y6R�_c|�[�	�҉�@�j:�&��נ�=�@���cz�|J �΂�+3�2�7������r%R�Np){6v\�+ =�<M}��:Hy��d���w��qm��Ǣ�Fҥ�(>;>�[�lhs$<�����L>�����tp>�-�o>=����y�H[�rPJ���H�����I��KL2[�-&a��B���ї�Ϊ�K�����&WDX�S'*�H��0�&������fJ�d�09Р� p�m�Di��7��KNJ�=c5R�%\�$}=w��k���>;P,���8�����,g�)	"{)*#%->��>E�����(�_y���"=�&�*������yz`���!��I�&ީ���(5(�Ɵ�P�Gl�*W��jF�+E�	�7	�=�χ�Έ��*w�!(=�ȶ�}�h���c$���ǔA��A�X�Q"�x!ҧ}d�[U�)���E�#+ܹ|��O�=ͩ��C�%qǀz�Ҝ�e�nm%�˟wꙍaKl��kw1���hH7_A�ƚ��8���q��U� �ߨ*P��r3���7<�}��o]���L�����&�K"�N	Fm�/���5���/�a�`H�v�X�Fn�,ǆ�����o�
���C����x�7�_�*���Ɨ���.B]�Z�QR�ܤ�#�ҧ��&	CC��.�,#�Ĝ���̀?W*�Ѡ�������B�$h�9��[Sf����H~��V�p��dt6�9�\�ޜ%^�q��)m� ���&���=�S�Ӓ�&�}����^���1 ����ϼ`���m �6@'�F�P����S�S�R��Q" �LC6��*�t�A9�=09��7���!ȕ��5Z�����n��d[R�.�L��kDğRG0~l	�FO .�K ��I�W3|��v���_���0�
��k���Y�uZ+�L����W�4Vm���)]K1qe&!#��~&/	��8F;�ߍ���ot�uy�S������S���(4=��}k�IYX(����-�*:޶�뭸6�,~&��"���Υ[����]�3:��\��\ׯ�9|��3���� ���b����z�l�S�l9���7�H���:������Y<�p1.���hP�ݪd6Xh�E�_x��1ܥ��e���.�fH�޺|͖��*{X'��T���A*�6s�h��^���f��4ê��N=G�����M�C_b���o��qF$`����K�?�������U2��*lpӳ.;a�{;�q��.D����/3�X卆��1Y+�Z�]�}����/t1�21�a���J4���&����%�{���k��K)�,c��_͘��9��Ye�ߑ1Wybͮ퉌F �,=sE1�JL�<ª�6�(p��D�wQ�%�&�F�?���xa�)F�6��/�����F\�d�b�Y�H���lã����x�t�Y�� C��IԌB�<�Tʋ#��Ӓg�Qy�{��;Ľ+��2%�έ=c���c��
��f~9nFL��_ef��Z:�;���BX��=f���[x�&�n{����
�+ H�f�zm�������)*��:A�6d��!¥�:��V�P�.+��u�|T�ź�ܕ�;�f�)U�A���l:�u[��c26"��ԭ.l4�~��mݺ�x��'�}���.JwEl`� 1�xPc��1�jlnDBP��O���7nT?���<tm�"����a��zX����@��E�U"J�)k���y8[�m�<��?�$
��\B���2H�~iXb��'��Ԓ ��4�"��R	��J�K��G/X�u�]ɾZ��	b����)n�|wD�K�`'�q�d?�*m_zA.�áb�
��I�hӖ'F6֚�NCP1H;*cH�oR��g8�����-s�<�a�OQ�5����phJ�1�r��L/�G�^�I�����,�2���^�����?�`{^���t*�$�����;�����ajq�}ˋ�8�;���+�|�6 ���M�x&}>%�φ�F`,�N�����s�mWds@�t�l��?����
�0Xh�WX�&}�����^o����ɟ����e���}���ή���5K�����b: y����h��m}=�XS�jR��;��2X��_�	�5	���P�j�ɻcS4B����������\`���ў�Aۂ�l�TY3y�,aP\JCv��0��	�����G�1�2��a�[HGy�α� )�jm8�p+
if|čMc�m��{G��mm]t�[`dr� \����I���&p��?f%{d��!oA}��ۆ�b�]%�Ak��e&����%��.G����j���rc{��s�7�TѦ�/g#�e\�Ke����/��h��I����2�Ok��b�D�����f���b?lv�To���J�{�	H'@�vږ�O���p{��n��H��U6��.����t��j<�&�	gZ(Pt��F�j�:�z34��=�*G}J��|���5�t/��1\ʨ.a9�a���{f�YUǥ��Wy����
u�)��7Uw�2׎G|[�4�Ȋu�@nS,�'�f��(���?�G޴k�;;���#X�A-x��gmx����>�!%�H<)R�퀣Nݼf�����rW ��KLK�K1�s#�=�� ���
J�W��;��YЁ�@�G�xКj�B>lK�o�=�6d%l���	����NY�c���~-�ƚ���15�ܐYd�ӛ��s�����\s�$��� @���$�>
L�ѝ�#0֙����G����[�F���<ڑ˪��5w��}�1�0.�$��U�Ǖ��h�:[M9�>`�>�sK����r���<DN����$^8U�"��N`��pM��z���]�SROeK�֪K�62��0ɭy~���}/�4��ne�Ƕ�_t�=���x۴s}��[���F��)����4Q}W��98�)���6p���g׽��],(L��E�F������j��cs*�%Jf�Vz���C����nk�� ���e������C)�� ��x����n&Y'ewq*�yZ���7�TjS����d�L�8Zo"���R0�U�P���?�w�]{�m�{�;㥐��Cf���-u�j2��y`5��[a��
q�����)ω+��S��χ<K��U��-}�����z�:ſ��D�"]�Q�Xd��F��A�	���|�K�l$��,DP_�v���]jx�(��Cֳ����I΀9��w�!����_���ȫ��<�4�6X4��ڟ����-��9Z�A[���g܆�	s2���;��:"
����%�0�'�-��oМL(4[�0��.P��C�"h�s�za���W�i[�"��YA-����!s7���h�������"�w8������-��n��D�7}$?ZÖ���LL�S����t�ڝ�6���I|
4��[��PUC�5 �ѫ�L�J���7�f�!�h�C�h���m��7ڢ=�+�u�#Գ���֋��j��oF��@��`���	����C�K��Y��w4)����6}�P�}�}~y8�]��9��?BszU�_���\d��	K��$�ÅGz٧������b3�|�CdY�B��b�0� IP�Kƺ����t@?ܸUH�!��6>��kٹ)~�p~��8 
싵}��L*xY}R�_�w"l������˘Ӥ
�,��-d��T2��2Uw?�����/"*.uޝ�d��� E�u5�#���4p���M�8���iXpW�-�JA0��Y��fz�{�o���⸼yt�ܐ���_Χ��?,jV���*L�C��B���D������p�g����+��Z^ҷᨮ;=l�ڲ��^5����q-����Ɏ��y������J��M�d���Hh��TC�W��(��c#Α4�����s�g�2
��`�	�g��@�uD�5�K<U�z.���8�ؠ�m3���ż�e�M<����7�L�Y��!�i�26q{T��^������&̔�7�2�z��Y��n�a雤ʖ�]U�(A�bf��p��9^�Ю����O��N:6ZB�D�YʸO�D�
*;8�O�@k͍���5X�܋�sf`04�� �n��}b)�SsA�����.���k��fH�{���訤?D��z�G�t��I���r�!�f\�)ɔ��B�Z��p��I��dܮ�����&F�c��3�\�9�&�����,����0���)J�{ͥ���*���j�k�a+�J��W�?c�7i��l���n�?R��'�C��d<1�0p�<�_�v�7ż�&�&nR����V�f-�zb&�&�Ļ�����ھk��o�{f�j��PP���`pae��D�|˼���>2� ��n��,��O]K��e�*�-�M홦����Vh[�!l�G��{��������xh��RCr�m=e ;n�~�`��I���V?�Ɓ�D4�Щ�4��z�e�H(��|xP��^��&��i�������c���Tklq��KtF�ު�a�7����=�m��@��˄5�*�V঍d20���� �(�ED4�zi�>��>���0؝��xR%��w{����I�������z�mrA��3�Om������ܡGq`}���6��~��+m�ܜ�4�3�E��6�E+I��zGKT�0��*��{���_AΛ�U^s㮣W��k�Ū�u ���xx�3�b����6�:��w���Ab�n���׹��k��Ӓ}M�+c�0*��e��~h��������*��R�6(pb�ޭ���᷒�>^���8]'}�X���:o�C��S��NzU(��mx�"�.l+�#�i���%5�����w. �^�	{>��B���BO%��.a��e��k��Ȳ)r�#�0��%�(�6n�j��	���|��9�������~pOO�G���a�7u3�[p#����\|��,{����Z��f��c�;6��%J��\�P�a��q��z�9��j���t��F�֘O�.��cp֩�=�� 0cS�ݍ�Q���t'P�'æ�ǯ��2�te�������P7�1:v��nU�W�E�Go��,�=l:�Ӣ����V�[3n��ᨈx�s���z���I�JQI�I}1��R�d�^�:a�\Ҙ҃��G}F_�/��/�>�I���+S��:�vҲS��V�`�K����M����X��&��?�nC!2�{�ǻlrDG2����?e?	g/��ۥ�>zY�)���#+uUu�ԙ���3F�}�f��>�1��8'0��6hU��/`�ד^� .Z���8�� ���(𩘧�8�9��or�{�},P�Mс�<��-�B�k�5�q5z� Е���� S�d��T���Jh�Q[�0y6���|#�u:��<(�㛚y%�.�טŞ^�<��h1%�p�%�<?�P!�%E�O̰�6�k#/R��,�j ��'��n�����L�<���hs�m\WD�E���)�ߦ���V���L-����9U*�*ID���p-�Cv�rGN^���������S֝(~�}�e����$�n�R�I­�a�험��	�`"N���nZ��)�̤���g!�!Emj�C�r�5�E[�ţ�Z�����R�b�����&�-�����TT��A8��e�5�@��0��q��о�6]��oN>�#	rF38-�=n2�* ~��j*:hY�Ϩo ��N!�m���~$,�s7�"��/S"�M�.�f��%%��>�n��>���j&�~\%r	��Ȃ�[��؂y����;��~E�xi~�|������Pz&���a.��Y9��<N�m��C�=�i5��;�I��#����IfG�ao�暷����oPYh��2_��b&���o��ۜd'�F�-?�>�`=�j����{g{��g���פ�f1i�"�1��>�h�x	]]����*�|p���e�$���z��eC�߉y���J��̴/�$6�|�����en�j��ڏ��M�ٲ,rR���؎��~IN	���=��~f���-i WW����&X��'���8t	־���>��"��#ON�x撕�2�i�]����F�lk_ z�NS����� �T	ca{ �pvYC�k�_j��c�M�~�U�J;���� )U%�:���~L���O�pnk`��u�[�����.�á��V*a��.i�Wֿ�c�E:E(����/4�;���%1翃�~��i�� ��Dz}��\�,1xD���YxPI�.���&���+�3��9�{-mH��n����� ��-�āj=�y���[e��qH�تc�.�î���yP����4�|b.r�"1e�r��$��>��Nd4��u�WH���mHo'>n�F&zE@���P��N�to�[�ǊB�D�%�/<�\�Z�P��ג���L�=��\#���wL�ƙ���Q]�$���W�3%�]�� ��8���Z�����W�UZ|�@O�:�$��{汍�
�b�R�EW�L&���Ы^CP���.
�N؄��i֍v�4a%f���G'�f[����n�^�j+ִ��������G_�)w�GЛ�������>��y���/�}�_O�+�*�>�6����"|�J�C����=zp�\1^�����\��n�m^�&�f���%��c� V"[Y�8���`���^��/�y#H%d�*cEkݕUj���Ky���;��Ʉ!S�'{n���7��.���
|�
�&�7�c��(��Kx��h�#��	k��~mz
�l�[�ռ3h��[��43�)/#N�FX:շ�QE�ʍWS�yT�3�����-����6���;Rϴ��J%q�JQ,�bI�J��5+Z��9\l���%�� #r�|z�!J�j�_p���T��6+5'ͱ�V�����B�,#��V(�~�d��������R��\�{��
���$ͩ8M�d|=p�����d���ġlޏG�8
V|�jLɲ�����S�Хt}�h���%�L���=(U�#�"��������>
_-Hx���N
��k���'m�..���}���(N�\H�f����T � ��9(W�dq "4b�`LMdB��~�p��L�0�V	Gr�y����H	��3�C�����\�ӛ�E�5�����V+���Ge��"!�}�p�A�5���s���f�Z�eW׫�X���e�����E-�����	�k�b�pG+�k���Hӧjj��aJTh������a�#(_�@�n�l��q�4�e@�/���H�h�);���N�+�S�0����W>
����XSB�A���ɭL��,[��]C`yKT|*�:��Y�XY��2�����L��#�9?i>V:f� G|�?bՠj�f�2ҹP܅x|�N^�K�MK��_֭c���h�&f^Y$�9�K�;�w	�f�
�v�0�6�ur�[��A�Ґ6%��_���6g�Dϩf�6��1	k$˜(�ת�.��̑��Y���N�;�1!����&���J�=����:X�Ʊ7��`�j*��R�� ��D��̣��{n_̛��=�5.H��Ӣ�a�4 ��|	�xE~i��d��$k�k��=�7�iF�5f�96�+#5eO�7���~U��
4a��Mg��Jn�U/P]��'�f�E�vMZ-�� +:�����r�!~ڇ�F 9�â�X���Ex��t��~�.�����L2{CG�[��u���!%i��L�:0�K!4�YE�jA�I���yюF����wN3�ԇ�TS��H�71z��9���7J�����4���=����Ł�Z�K�e��(�M��鏤�咥�3�T�(�/��'���.}r8�!�SY�e�c4��;���3�t�>�!&�ۯ#:e=�6'_�G�<;0�nฺ�J���x�?pim6�QG���[k���ԋ8Mc��K�O��.x%�-"�h��!&ӝh�= �"6)]����~���dB���s�L����h���-�|>��f1�H�+}��a�� R7�d�Yq�kب�r���S��U3�S��A���&S�ә8^�0^��� ��j�8;�(=D?Ϗ�V�E���T>w��G�V���l <."y%����6耄��h5k�$�	������y�o��i����\qQ7��Z�6{�gl�Z,m��H�2bs[��)틀��{ltG��#�ᙖ�0��!8��{4hƠGH*W]��(s��Ԛ�K;8yс<���Vj�?�����휭��9�",D��������}-Y�V#-⻖P�	�j�y�E\��a֘����֋巌��$�
���˙���9��3��!&Rڀ&߳|�d}>��F�Q���o��p%�u�5��Tn�>�F�ӷ`����͒bw��c�(@~�d��<YAQ��<^;X�Hx˺�%4�����=��ᛍ�m�w+P�Fld�/��
lM�(N3�"���$�O��K�d#����p>eГ�mO�X ��Y�b.IB�t�K�ЏnP��M/ǘ�}���|���9�e<��t�#�j���~���9��S`��Q�n�����ݽ5S���T|��֣��?=JW��>.�c�H��Op�ޅ|�q��p�����N�9�&I�2��ڰ0�c��R�+Vr;�1���ho���U;���g��?�:��o��~N�y��@�I�2<e��䇭QG�:��z��d��Xzf�=��� ��N��q(��o���ba���\b|�
K�D�"��0�4H>8Г����̻oD�=�c:^ԃ�9�r�=���0��l�O���1#�y�)zⱿ�\���,xc�'�:K�v}����R�fԩ�����oWC�'���1K��E� 1�u�bX �!ȕ� M���Lh��5RT��2ˤ�>�i�̇5�
l���2���=΋lƛX�,1��,�]֙2u�-#�y��U�3�O_�i9C�g��y�|����Vֲ�CV�>�t+�LtJ��)�*h�U��u컻�6���5��!&٨8rԽ=zIbӣ��e�K��EhS]�fw��>���T�[w��#/�����@hBp'���C�h�F�d�ɺ�W� �J���\���9l�?3��,��������Eh˾��C� ��xuF�!���n�d�WI깯��m>2�\�H{n��9�&B�#H|��kgI�- ��PA�aZ2Gu>0��}t��"�G4�l9��F��SRe�JH��|��U4�<��g��~.|i4�@`��U�U�!�$�9�Q�~0Z��1�՝�a"�`gV��ev�?�" �.�Q4�x
��*e	\��RCAs�2�6����\]nKȥ��RV+���C`��D��UE�8B��Zt�yõ���P���)\�]����cP��T�|d�mJX�*p�}B�L, *Jڒx~�<�Ss;�c��3@����'����+d���S�mĔf�,��v�=�� u��]*���V���_�������P����zOf�R\��z�4�+�Τk�Ĉ�ƢSA��������W�w/���\�b�9���Ԏ�{���T]$5���
�-Lt{K�ѪXa����z��ـa[����������/��f~����3/ҁ5�4�D����g��H�1��\��޸����wJ�&�@"��:�G�E��>�=�@��������:(j�}��S}�~LZ��k�?�p޽��'��#�mL⁼;�@>J��93�Xb������5��9�,蘲��R�n��N�44R����i/�au�y�����Z�c�D���j�逦qdj�޴
:K)"k��hЭc`��g��yB+\�ff|�m���"����7 ,�4��Ki�e�7k~����α���6���jjDm�_R��W�Df���T��+�6�J,p\�Z���X��c�i���L�(y���'}�i���P�e����8���[)V<��R���p�A���}��1Q0%n��z�P�'+�����@P��+K��L�L��>P���M��#Smd�֙��E�Q��/C�$#e��?ɠzaq�cn
�\�@�Rg]/\*�#�gi���\�+2�w�*�"�e��XWmrW��bKƃ"��&y���6���E�l��m���x>(i���������"��T�.f;̀�T��#B�s!�<������S���5�3? `�p�UKWA�>uK����g�]�V�wXVx�'��b�XF}!��C!l\F>�;P\�r�~�9Ft�_��*�
�D��轺ʦ)Fps
2��J��V�8����_��o�/
S3a%�,�Up	N�ӑ�o�꼘f%n��ҥ�z���wM7/�I��2@q��/���Zh{ϩ]ߟ��v�I?�
7Eh��R߇=��̞�d�*2���MCQ���B��asRѾ �"Y��b9������+ڎ��A��he�ɣ��@���ӽ8O^E#��TS�J����ZF��pCk��,B�Ȇ����m�J�Tw�pʈ��������&.&z����%�rKV���t�e(f��w������	X�f�����(� ��糒 ��L�?�$�qT����S�%�H�v�N��^����kJ)���$pI��>%8U��'zu��J[�O��C���n�ѧ�#�T�Ug�jS3�%�|��b��e�A?��lH�Wp�o��ٝ��w�h��	�F1�	:ĶQ�t&��m�/
3]�~Hb`뒟��RR�+K[��p��ɶ��x�xn<c�}!(\��$�\ꓮ�@,�T8˲�6���~R"�5�.���$C���x9������E��v�������F3���U�!$ E��-�B�Qaa�?W�\^�e�֬�A#���Z�+�?ZW���y�{2��(�/[u���M���{���^eCX��O�r��y}�U|�
�Xw�����R&�c�vW���L���Q#<������9���	L���_@�K�ϊݑ���.��v摝v�*�D��hJ��R�=�@Ü}�C��;�ᳵ��X3|���Py|��<b¸X|�'�,�,�e�e�y!h"����GJ��D�L���Z۷�c2jl�EƩ���78���2��C��3M����%�)��1iޭ5�M��K���j.����Vǎ�
L���)�nbג�џ�d|)Aʁ�ǯ��՟H��L�"��fV�W��v����,��b����%n-dؕ�72��aI�!�!h���S���!T�՘��S(a����P�\`s�>V=4W�m,���*���H�Y�WҮ���Q�Q��;Q�xa�Z&"�{�N��(u��_����bO�Uݿ�(*\T�3 �`��{��q�gc����?���a�ϖM��m������_�sZ��y�W��b�YEAXF��f ^��e\�_���c�>q�uKާk���a��*Qw�� ����Y�`�G~�&3��í�*�͟�)n	rC�Lq��z���3���SBbVw�y\� ��R!i��1p�#�Rn�G��M`ԹL� �#�?~ыF�e܁�v[D-
$S9��t$�ǵ���Li&T*���8S�d<���M�E�H>R+�߳D[bO��ʃ:=�M�&A+N��S��C��~q0��Z�狫��ӿ$zRC�7)�lQl��Rgf�:~V=lZWm�1� �,�f��cG�(R�P6�^�s;ߤ%�|}R��3d���k�҅a|9�
�S��)5J�h�\�}q� �홲�+R+8��a�/z� �������\�H�/�Y��F3�l��.AN"���)K����������R[�9�׮�y��&<%-��/�^�N7e�Q�@~��������+d���"w2��,�ȭ�A������[@Ex�,�s���r�F��p"λK��gK&	j"kQ�;i��6�Lb�m�j~mZ��ۀ�T�k�W�?�Q���P��%a���tu��5�^�B��ჶ5�?��Q��!��?֗w�|}T<{둈,�nz7�ly#e���e98vi9a�� C$oP]C���W�V]���P�!�� 5!@MFNi���(������uE&����*#��t�|\��00�|u����N�)�^I3#�1���t��񡩔Tw�E�N@R�*��5;H#k h��nWk�E�տ�S@�S�HV����Rq��y7��)���t9���������.�F�f�����X�EK�)�v�εК�O��T�/*�v��r�hj ���EK�X|GhƦ�'�_:�U�=��!��ޯ[�#�"u�{��$��Z�������i��w���H�ff�v��D�i�i`�7��q���^�����o-:m#�/�N�z�,a���l�G��4p���ӭ�aTޒ�N�S.V- ���oqKҢ�{:�R�H�����YMj2&�6������Mb�kaY��b�@"]Ux�*UZ���k�	�P��ϒEm@>j���B`
m��eȮ(�N9���FvPb
J�/An,��aA+!
�}�M��u���>�/��?�]o��_)��uֿ�V���Tm��lg+w��7ʷ{XZj2��Lֳ���������㬹RR�Ju�ٽn 㤑leHJ�=;�<8�����r!��Ѐ���p�>D�0rJ�{���I�J�X��*#���`�~0ہ����S0���,�����'��'lY(<3�@T<��;vn�Ƴ�$�lG�i�]Ê�k\�Y��-��l��Z���Y�,����LMq������OPp����6��3M��!J�[�����-���Fc@6}/g�d�eQ������QȌ[2,����` ��(㫼'.~��8�[1����b�7Tˆ�򝴤7��.�1�rVI�ǧ#J���g����E�Oڏ��w-0@)�p���8��F5��'{�e]E�B`��]��PY셨������dR�3'��Y�k�Fy��}�m�',�����N��a��0�M��V� �X��r��Mw��?�_�[Kf�UQ�
tt�9�������^��ٔ%�\���?���k����9]�X�Z:���!�u����24hV�kۗ>��i hu"�mC�{ �x�"���i���4&CK
�C4�L�=Iʽn�bB"���:������Bi7�3yL�	?�-����`�X[�m��;m��ܛ�Q���Ŝ�(ү�\d?ko1��"=U�l͝�(2�e^6���\���jjAi�H(��Bʏ��T�c_�������W��.�|� 1cʡK)��K�5��K8�cNFzxg��@!X��Z/r�sy�����W4&�yۈ�DI� ��Z�����C�Ji����H*w�K d�|��+�6C��<P�t�_�s�$���=� %K�Ɣ�>��U� `o`ie?N;v�ch����$�j�1�-eŨ�[�s��$���:_�a*�)3��%A�Q��P.e^�q
�1��8=b��`P4�2��dRȥ�=����ne��E��4���,X5'`��j��S���|dX�^�F$v��Z�����.�-G���%I�����bXe�l��dIJTQ�#�"���������a��-O?
�%���:�b� �$LM��J۰��5�<Xr��������L���D��Nv�=d�<kр�Z]m _8[LV��b�`�U���Ϧ�5�?V Tiy�lm�Y�4���(-��Y���kO�A�� ����� ��-T�=
�U$`���L˫�WB��'|�OE����d���=�K^����I�i�2�:����|��k���`��������(����<v���E7�������Y�1^HH5�	����Z��"3����;Hf�֤@��u����u��E����p<���u�z�������ª;�`��� e�>[��&�V�L��5a����MEJ�3a�Gl������*d�3i���Q��N>
-E�N,�]Iu:�)׷�~vQEt����n%�*��p�R���xT״5�#p ߊ�[#;��5�l��c{!|G``��:X�fW冄�>�ׁ#S �̪���Ӭڛ�X��ۻ�?|p�R}���J��F�(>��]��_B�Y�BX���d��݌��8���Q���i�l��ɂd{YA�@���QUE���`S��v��x5�02ҮTB����B=]�5,<�+�@�"��	�Ën:��WwQ$RP���?���Y��~É�5�J�ޫ�N�e̳˪��_G�����v8u&��G3�A>��f4}��;����]��A�P��mfQ�L��\;�i'[�ޭ �Q|�䂬��h�M�&��� q�I�$�wX�x�է?ֻYmCĢO�pC�>x{�&�D��JړoM(S�d֞���f�ݚj�A;]��VV���>c�ނل�ÃAUt�~�s!ٲ��� ؼ��5�A�a�����\�(�x�P�<�����,�]�-Bzz^ߊ]!ﱆ�T ��iKI�����U���:�~j���+�{7�u�GO�̬�������F��?��5�_K���D���WE��y��.Ø��=��;��_&5D��(����q�{N^`q�q���ȵ�1�5=la���Ǩ|�B<9���G�	�]�Xf`��8t��O��!37b��u%�¦���Y�sX��&��eL��X�ஸ$��Ug�m��Qu����'�*�}i���-�C'���$f��\)��q|��������j�I@N5�?�@r���1��\K9�Z��dg>�,�H� � �y^��|��nmTE�E����
4h��T��"ݚxs��������`�-��Y�K<G�� ��[�h��tOsR�F�:G=�g�p$㹨���1c�h�')kv�M �j{cd-]cH�>>�Ɉ�%��g�ӂ�@)�n�������s���c*Ja�8�Fb@^��L0�އ�<���hU@�ͫ��͟E)TLM�Om	�q���t��	���*���lA�b�)���,��ע<^c����+M�n�~>h�@�:�~?Ҹ��iL�y��"nTJK�Xl�R�W��
�2��
���,o�C
�倏��&���r�o~nT�o�X]�=bt����#��В���3e�l�%��B��\�R@��ba^3:�G�Y�p]Z�k�����a��?��x���!�T֦��/hļE.��;�a���5M
JB��|G��5��IU"��@�pѩ3��K5��#Ixf!�͵֕\��H~�7��C���c={�0L��84�.�����/��ՄvR��,H��m	�Y4��׳�t/
��٬�	o��U0��Yӷ$q�$g�����}�PV �^՜���W7X+^u��{� ����:Q ~i��>ZtFz�b��_]T)�ʻ�<�>o�ˍ��řى& t��j�B�ܑ���P�8��D�{�r������!A��2�3r��.��Xx�g+r�~�7bVɳ�j����7U� ���2�mbE��&0�֬uhC��f'Xm(�k�DζA��&sUI�F�t��*s�e��s/j��	��8���I`^j�$[�B�X� Z5nr��@Np'�L�x�m�nޠ]���~ě��)�GH
�k���n�~��N��D�Ќ���S=䂗�Z���X�k�e�����i7&%�fo�OR�c�ć5x�W�;�2�%�>�6N�k [Z�2B�1�sȼG�B�V��(�^79���A� -o(s��[��	 P���i�<ִK��R��Ly}*�t,��4z8Q{�xw��06�Gu2�w���p��/ˊTi�L��hR?�_�걽UD�9J�+��}Lx5��~ұ�3U����!)�n����?�\E���ctȴ����g[��Î"e]�p�\|S���pȓ'':s��G�v�]C��`GxP��n��FTSR@q䆠6���Wj��FO�K�*�H�'.�H��G%���7��%$�M�4��f	U�#�Qa�Xq��n�uLh&S�>� !��0:���������{��z���+1�U%��HU�~0�����邠���=B êvb��x�N0�>e�u_�����+��HMe���]��l��+��w�)����IS)̬Ei��L����N���	ٔ�7�([�F�� bFOm�]O�S��>��?$�؇f69��Y7TE#ϡ*�>"2H֘p��ф��n��3�(����/��k(R��5�1�k��4��v<x5��'�����C��V�i��y�d����D��B'�������!���l���D��0b8*�P9Y�}�)�B7)����|xi�q���f���D�ײ%���ߙ$
�1eg��עSˁ}�z��`a�0O/:v/��*d�d����Li��ܸ�MVu���AY�9N�D dsp- ���T��6��p_�HV�N�b�:j�K�|�N�x7-j���3�jS\���B�������c�������V�s3~�����>Z���F��'�ſ�r#����p��me�(Ny�_����|_�|�`�H��)#'r��)C���߾�������h�z
f$��L~�D�HG�ƿ��"!������+��|�Q�Y2��L+����0�D_�KA���р؝��>|tG6�ۆh��e_]�.T3S�����+	p_�p�Or�˧uM[]Ё�U�~�iJ+�5ʑ�� �! d�,SCǷ�g���!瘱V%W�jh&jEq��"&����#���H�K1o�����UJLn�V�'����-&�}b���W���c�;�3�	z� �`oy`�J���\u��s�j�~:��"�Euǘˇ]a¡5����+�d��{"s��^���a�˨�#���as}}ޖ.M/�=Q4m�B9R��Z�i3���B$��S*l#���
���,7^!�Xv����r5u�s�t&yk_����~�t�jnnʪ��+Z��o;������>Yz��hE�I�q�8ٗ��O�"!:oI��!!��F�8�d��4T�9�<r��Jg��%:5
��p5u��D�r
3�3��X+d���5����j�4�3f譠UhcV%���̻)�n?%�;'�p1}uuĬv��A����6E��Q:���H�ZB�!�=�l/@1�>ȱ�����Oj~�́L?K�U��Qa
�
�"^��d���|�3'��{�4� 8��H��t?��7>��!��:��$�㰄1��5�s�cQ��^o(ߝ��D��ԧ:�ޖ���E ��M��2~�9��rvdc�f
\�z��m�_M�ah�ͤ*�F}�y�m�M?��_/���=�k�i������G����� �ZQL����L	e-,"������0�к�b<�g"�sD�@�J��ɝ[�{@hfZ�a<z�����	����چ"�:�޼�Y񱰁=d��$�U�T%-U(���,�����@x�t	U�ݐ)ub��m�C�%/��/���m6n�G&t��<��@��ɣ������w��̱;�06�Ҟ���Cp���ҙ�4D-�W[�F��I��V;�<��)y�"::�	m���
;4~`3���@��Ox���∭�r�o�/�BBC@�e�o��Z{�bHK���"�[���mz�c��DC~C3��t�`
��Č	���Ce��� ��l�M&�N8�<C�}���=��N�Ϯ�x\��+"�EZ����\������ak��F	��G�6��R��J�t��k�"���ʭ���\��̸�'�\9ȋ�jS����| ��x�h,<m��u�?΄q�r%�B�:�9��!c�xZz���*T��!�6���N��,��Z5���Ww�`�ľR�`���gm�g��R�N��(E�\ש��h)�m��n�I�H�x��)1/^�+� '����Щl+����ISS��Cix6�oڿ	-NH�(��G���1�Y(�����M��G"�Z�`!�E~{6��JO��n�Aޒ�n��w��uQ�R%���1|�����v�'��a���sgE��ρBا1�@y����]�d	fOZ��ܗ��|���G�)�WAX?Y+�L�l�h	�����G�W�<����n0��+�SO�V<��И��KP�lK��l6of����ƽh:�+�q�0 bw@���U�q��cI��
b��t�awpH� Ï�x>�p�K� D������EM�ӏ�N�)�J�_k���GT����w��;x�⥙���ǬTzb��վ�X����R�ŅP�Ձ�7���"!)=�fm�X�(�����#��<v��(ot�R�%.�R��ΐ�T���c�ZL�7���	zM���f-i�A��H4��'�K}6�0nn��j�R�M
(���ƾ�p
3�m���/bV��om���� W߻K1�f�o/2����V����������8e��Bd�^��n�w�)���(�����Kj��亀'E#�Dr��o�WG�1�IE���h��.�����^UA`���u�����䋃��`�,�tTU'�8B����	Ļ�8�k��gWQ��!�S.�2(����vl�Z�,�`�2��������<��VV��A� b�:�S������2p�z�4�#�:UgZ@\8֬��"D�E��0T~P�B>��L����}�I�|�����:}����ߢ���]ު2�����n��p��-�I�@� �
Q��&KX�#dDI`,���?�Ǆ�kz����e�,��S�\xxk��du�2&�V�-`�ImN��82tH-L�o��</IYƍ�_dS�	:�[���mP�g��GP5�<>�_�-Ս���@�$�ya�%��M��.���be�Z��pҙE�ڍ���
�l����)���GC�q�$K>N���X����H�K� �S��=��X�'(,���$�û�����ONL����O�{�<��ec��;��߶ޣ��m+S@6����V���e�����Z�(WA���|�j��v��"kP��qp&!�`]h��<���M�
0C'/�L��8�ѻ�V��ɍ��S�t[���~uZ�2��\�{K֞��8���uGq_�@v�̌n�#�x]��^�f��3ȕ ��h�5b�jih��s�y�U�X��j�L�����w�LP�`k��cI��R�����+x�K��dYگ�HK,y�-�s��&l�������N�ӄM׬� �z�]��������/dũ[�����[װ��؍��ːot�i��N��`�*h+4J�m
����� dy`kޕ2���T�5�� ���)��c�Y��ͱ�\���ɜ�#��oz��Dm��
�N�)Q�n������Ke�И	��z�r[���U�k� +�R�9z���l-���O��?��d?�,���8[~и���Lĳ���;�.���.l؄�v�5�	�Z�M��0�i|K�a�+u���#]I:#=��6���[�)nYUdWp�1Wă�V��w�|Z�>̰��O&���#WA1��@8Z�4l`-���'�壛��y�Dܘ��sm1V	l�d��ǣ��;Y��aJ�U)ʀ�{zY�'��Y�#'��3�����̬��nO�Zj�~�c� $��`�K�и~��}��鉃:���g��~5�&�( ���m�m$�PӨ۞�������L^ �SbG|�4g���R>4{E( EKe��X'�W��5ɀ�е�m�Mt��?IX��'��� X�m:ڈ~�����5X�yֵ!P�WP�G�x���Q)�OhϦ���1�%t�fڵ�=�*1Glw��x!V�`'Wn�p~Γ�L#��$pv���8�!.`��}��^�4��n�S�GC(�0���2���ld�)oF�q>|5އՍ�0��4����tv%���E_��q>1ST�w�; �����=O_�x�"S� �V��aw
l�ȇ�?ugx(�)��'��oFM"�PE��H��ر��c�Q��@�T��X���2��9V�P����p!%(�PX��RX����h�-�'�6#p*iu/�G��੮D��' S�-h�	�P�	;|yx�~�r�:����+�>��T!�q�\a��~�����i�����U���� ��.-�J'������_�:�!�H+��2��� 0zbMy�!)��7*�a�h�
m�.r(����7	��-�J��Z�+Vz]_���g���p]#}u@$m<��%�;�[H�vc˯L�#�E�D��9�h�p��m����-��Jd��^����P6��N���zQ{U�k�Z�$�V��%�R6��,��p16;#p���7?d�Yr��2�<���z�K�������d��j;rZ�occ�=%2�)�����[��@��b|ʁ2 vR��E�XbE��ߺ�>�>-T���_����հ_��kk>����H0�y���{��{���a�\cd+F~�����;Hr��߮���ZF�U,R��tp_���Fu�'S�����-�n�DlK�]k��?�{�¤ vƯ�v�%�@6���}T{u�w��]|u�ʫ��<d�V[7Xݵ��0��6������,x<�2=��s�H�G�����	g~eS�!������,5zp	vH.M%C"�����OM�c�	9\��BKi6�!u^,;��(^P��	�ka�j�!�����Eƥ 技D�1�I	#zW���՘��,���-گ��{ldkls��`-��݃h���9/J�BS��yb	Ϲ܃L(�(8����S�Łt�����<�M��IF��[��!㖚qT��5�;C:2h�����́�Jt���H�<eW�H����9�"R�M�
���F�t�I�(�@�o�]��#��5��4w�X��Q�V�����������S1
v;���T�- ���p�|�A3-�֐M�F�J�n�YUx¨q��ZG���z�_�cY��!�y�^J��x��u�£�-��W� ��ľ�ƺm�����}�)�t~~ʵV�R��yD��跔򼕧H=�=K�:���8��-�g�|L��i
�8e?F^��Zm��T�u������E#�@�{����w���׸���Ϩ
D�Y�,��Z!T!���b����DNY*KT
`͝����]� ݡ7Q�N ��dF����<���s��l�+f꠼�3z��>q���O�ߨ"�r����觴w����V�|Co�󭥹nP)v����T�"����T�eCMWs��W��	�Ӈ�	&�j��i?E��9<���F}ɠb�7s��dݕ��6H:^���Ѥ^���r	lg��G_�-ؿ����^��G���z�Q�j3��!����3���l&�,�A�H�՗J�7�� ����������L1�N��v` ��g�(�D(����6�����#}�����X��Gj�~E�	a���A�0d�Y�]�{��4>4f+��N��G�5�r�.ǈ6z�r���/j��pU3W��=o�MRO���������R�ӊ�L:���F�	�e�5�߱YNRՁ)�N������C{�;�	���[���e����1fe��<#�Ʃe/�AS벓\���R���%��*)���A�:�����/�TQ��~���B	�e�J��7��w,
^�)��^؉r�/U,_(�'b��iUĳ�K�]ML��RiR�`�*���[�SI)�,�F;$35[}�V_�I�?�UIA]��Hl1ќE���.���?>]2����VD�`e/zuִ��:�"�B7����o�)�I|�2Da���������@Kb����5L8)O��ɾB,G���aIJ�B���)�%�0�-��,A̎��o"#���Z��/?����6{�F��`^8ϣ��?��T�%W"f�y�<�r�m�*ꐜb��Rs��|m����Z{��G����qf�*�R�V��/�H�e�H�h�y)��x.�!UD��ǿli��`&/����C/3��Yzn�]5XK��w�~�:�����@/4���`/Ŋ�V3&�U����>�*>ç!��l�v��K��c���S*l?|(&H�p� Ir?��hȵ.�CW�W�1U���qRZDm|���_H�$��S3�N>.��0G&gGL�(E��ߎϯw�Q��i�K��k��D�L��|���5]"�4�\�Mh�\��U�/�_$M}�G�5�$������?����g�:1tl�,�B�@����-9�� ��99�PW���Pd�����	�������mRɰl�BxmI��)�ڨ�"�lo]����r����E��DN��֒q)�-;x�A����H�BJ>�ް2�
�rb�zՈk`c��ԯ��d�g	Pzz
u�k�1�+����}�[�]��T(�!�u�{Q t�h�+ҞRSh�������gs�\oơ��_���i��b��cN��!���p���Y�0$)[��O"�i����7A����%Ĵ��&��尲�j�any�yW��{�[���(�w��Z �!�]Y]���"���%-K�~I��#�ȇ]�K��d�-Z����o�yes�M;,D8lT\w� �M�����_���6��K��-�8t��M�T(��G��!��,�C��
"}7l��DE��sk�0[c�c�S��@��8�X��h^f�#��T�,�qj-���-��uj�� ;}\����C��1��.�"8���FX �l��[�ř��.�~">��alţ��d>̠��ec��V��up�֦.#��3�r�T��q�J��tJ� Y!$V���x�T���/+���ߚ��Q1��k� p�4���C��Q�V6)b�����cf��r|�
�9�����`�t<����@0�X�P�ȇ�X�( U��/��=muS�/��D���#�A��B���O��J�#�p�FF�ǚ &�(�r����5?t���ф��T���(�������a�(�'�K?�$��"���Z�!�O�,͛E��m����!z��=2�)�B?�C42P�δf�{yq0O�q���a^c����\"�s�ŝ���%X�脀|����!9�[��R�����3�4�����b�A���{��35��w��>����\��g���lR�ߘ�1yQ�W��LhN	�mM^�^Ncê]]���nխ�?���y*�Q��B��g��M��Z���J�LŻ/�	p�[E{Ct�w�pMy��@"�����%(	ҽ����D�W�ڔ	w�*��+j?�5�� ��Zxz�*oƄ���`��Qb�����@^.�Qg�M���~�D�tlXez��f����O�_Z�����̔o�M�^������!�>�Y6��"ٍ����l+����z3��>���q?X��{��*�̵���i;�gWɾ������U�n,���e^�)�߁62�-�M� -����i��j({E��AS[֔��)���lilIG� ;�z���+9�1hw��pl��V;Ed��]P&��4���K[%5Yr�B���z���/^>�y��/������x��y`�5�E����@�&�����Ĳ�$3�CI;j�k#��B��u;�XTW�ZWҦ�Xx�� wRu	&�c�Ā_�)�؟Џ!��`;;�J�)�B�KY���5�r�y.+��ԇ5�	1��h烽x$�oׅp*2����j��g�$���0D�U��=8�����l@Q��B*������ �;���`�L�'�������P�0���ݴ�Y"� ��QS����ډ4z�!��>�q6��Uʪ�S�h:w��K��[Dn�q�7�>tIȥ���5��[MJ���B��ت(��'&;��2���\����W��]ZB���5��_,��U��d���/Bl�FQ����]I|�龻BB}˵�)��5NT�n�s�"Y,��v��2
FG�y��vE���Ii�̲��LzN���H˫J﷘��r蠰���-���%���֮������#1~m��1@��hX#�U�	�7�dxn���a;\�3FH�D�*��l��v��zD��,$�9�ou��E4�n���F��HoYһ�s:�äޜ?������Ѫ��/B�R� A�*�WL�զ�Wޣq�b�v��]�Gň��:�RL�H��©rŔ�x[\������ִ)d�NL�C!*����P��Mw��3�٘��=���n�{�AK���1`�x��`�܈�,���YD�|�%8�� ��i�݊D�cs����j<胘y�됶d�Dh���X,^���&C���X�u�%�w[AB؜��г��7�=3A@h�X��N��Ie�]c(uk�Y�M���r�L�	y�B����&`cЀ'��"�D��P�*��8�� ��ѓ���8?�{��O�K$Ukŉ��
"gP��BeJE.��\q_̄��\��6�u�T��P?���C��o�H�Y_���|��7P����kb�k�A(sc;����M�hB���ApQwȪl��&Ӹ�c�{���s��ԭp�t^�੓�H����|�rH��g��{
����Y?�֧r��[�r,�#��2=N���ʥ_��&Һ��r�� [�'�S&�4j�*���P�s>(if:m��Ą#�F�j�݊}&g�����cAݫ�5�<^�^B��U�� G���"^A�q��ħ��{s};�g��qz��#�R��Q.��x�r�A���N�O�L�=�c!�?f*���^ay�V^A#87_Ģ,$�⪫@q3�����ڿ?��pF`~��o}�J����	�|<[J�̻�ߌ	b�.�៯۠|�	)=D;�JoWk2lv&\.^i�x/��:V?Z��4��ޚ�ӝo�k^"���i�"��S��A�9�oK�N����Ҩ.�ވ��A��=��_�0�{*m���P8Nj7�z��l��GW72�z��2o ��,��_i�t/�K8������r��h0SLAGG+wj�5��w-�e�:8��{i� ����s�ߡ.Y���+Z��2����%L�!��g�+	wό��w�OPu�D_�6�F��W���R"T<D䡇�t4ޡa�B)]�9�~�(�l_W4)Z�K��S�_U���P��(@��h�l4�:_��O\s+�q� ȕK�X��$�IP�(v��=4ye��NY����N��}��,V��~�t�tӒjr~;��G��h���Z;'����ZƲ0��bi����i.q��	"�<nв�|M�3�|���0Fw�Z�uI��b����z1���L?��gY��P9Ҭc���k�4x_ف�Tg���P��*/K�tg{?���5���A5�ڈ�S�>zGٌ̕����u��yq�3U��x�~�,L���4�r"��xh��!��h��ū�3�b�(\h1'�G�'�BY�Y
$�GѦoJ��V�;�*�����%�A�X-@\k�<��&���R�����Օ.r�$�C"�8�����dR0�-�!B�&I{�jj0���L���0�k�U{O05�	���R&�<��\�"ZB��}��C�VZ.\_uU˂�?����Y �����ҀB���y�����^�՝�,9Ձ�j@���wrezt�W��{�����uI�@k��ځ����u������\�=S'>��V/Yl2O:R�:�s`Q ��&�gd��56���|��10fhM?-_�)
.]=4Ip+߀g�,��� �0���;_��!��#����� ��25ó\���Q�jCKTy���_��fj��Hƨطv�
�cŎ���:�Z1�������Fp5n%NXHO�ŋJ�����QE��●g	�����
��W=�e��A��-K���7���=I���%l9������Xa�F�a@n�{��HA	Y����
`[6�>G����s�8�?��f[���15$�&�η�t�܍[��� �X�b_K9?�5��km��|LX�\=`�� �zv6.C�T�#��L�U�0ӹ��~<��M9�k)�P/�����i�~���������&E%1����	2Ra�-��-�^�wI9�pn��߁�Ы39jW�_�!Nv�o���{��c��6}wR@*8ٽgu���ݵ��6��j�_��ģ|/³a�(z���C]z+
@�zi_�ԡ�8�k�Os������25wx���9�ոt|L���p�����!�N���̓����e�h�v�����}V���-���}s%���VL���v��.!�L�(�g�����	��?�U��X�X�z*r����w�ä��2(MA��VY�����N1D�@s� �Q	R��5����2C�Qy�3�d�`+p{G]���w=���PK�k[ �O�u�0��@BXV@��9��RĨ�AL���;�o2��&N�$'���$����^uF�GصV�Q��S�I$���� �7uc�Q�J��6G����h�Ԅ����sH`�-�Og��"��`��y�M��gΓ��z+t���m����7�P2�p�8_����X��?B
�{ [r$�������F �-ӿ��!ۡl��m�_J�.���"�mPu��ZuyaTϧ[M6�+����!x+QE13�~u�1���,��D	�����g�}���zp.�����g��@�+�P8�#�)X޶4��/IR�
{�Җ�z��"�EyŘ\,u����h<�� ����(�o��v�l2$�^�@HMA@׻ ح�m�MP�m�@+mĖ��7fK����0<�J>�K�@P.`̄�H9���Ħ�y��b�"����
�.o��|9"����W⮠��<�M� سg(mJ&���MD��qn����;yR��I۶)�>��ib�[�.�.���r����m7ߘ5���y�YN��De>�=V�I}�o�I�5���v��Mg��f�W' r��<����ϺG
E
�4L�*ŕ-�2>I�RE�6rh�`��8�(�+�R.����n�|�y\X1������x����<��ԣ�@3W%����F��{{�؀8�,�(�{"~!�ǏC3�=(�?
���x����6�r8=��pߑ[�K�*|���Y�ǒ�ih�|8}��M?�R���n�sp%����l�7Y�h��Tc��e�6y\CP��W�2��� �n�ku�c�.�.F?��"�������B�����qM���QS2�%"Q��J����c�#��d`��A-�-[���0�B�6t����s�� �Q�'��hsp�%��"�*�w���?pTh���Ľ�˕b�x�ħ�(����f�+�ա����1�K�q0PN)�dփLSH����ZڅDL��cDxo��|~� --=e���p�r2C�ߞ4A'(]{���w�( DM�,8{{�f_��r)�bB��F�l�_�5�l?�\ۦ�A�EG
��� ��d��3}	v��L��P�$�]d��=Zl� ���:����-��NRA�bb�yAj���1���q�}�^x��W8�4}d�d�ߊ�%;ѵ�����WR�}4��i�W*���ȕr'O/v������^I����N�&,�cr�Fr����6����,EZ!��w��ႜ���\��*T�!�В�eq��|R�K�h{�_��x���gU_nA˯].�{�/��UV�Gl�^>S�����9��4}������A�ĉ�.& 1��hYfݢA �������ꜝ9��hM(a�+ �K�7�nE�����#�&�a-4P��+�!_j45�[6w��劁���OJ�١9�g����2����(�n����\䗱���{��ζn�Ӳ����c���ea뗏�?�~�?��fa;�R���|'\>��CҶ�x�\�k�H�[�@$�0x���(ߓtG��������:z{�չ��yF���{�wC_���y��5h����		�2�׫?}�[���z,歊�r�f�H��μ��"�h��Ng���GdX��T'������l&Xk�SB��J��z�Q���"PZ �rt˓w���g<��QJ�����2@^6b22_�*��-�Uǀa�M���4��"�ю�j'ͱ�\�+&흫�)�U��c�|�rɔV|����*������e�ǹ}oP�z���<�i�5k�)l�'��E�)�rc�1��ZMqZ!�gK�p�Hu[<R?[[�į}.a?q��o���r�)��g,*2Q}�a���`c����}�#>�_j��9D��Bz!�Js )�b�T�<u�=̆[����(}.6_��WN,�|740�s£r��g[</|)���)�ꗠ�# �?�6�c�A��2�TU�Ԋh��aܭītL=@m2�Hn�D'�;�` KB���߷[�����{�V�𿬩(�N$N��Ü�T�O�oP^�4(��WW���? �2��T����g�W��d(����Tj�4X<J���'��#As7��ℤ�qu���,4Z�{_>�JB��YH��ԲS�͒'�_�EG�ZF*�u�%}���d��P�J D��ݑ�''"�6i���p����6��X�	M�B�3=A�
�	Z>���]��5���Y��ǝUzv�\g��~���f��0��\X ~c���D�?�A�4�W���@C�j �勂^��M�����
"\�]��b�L��7g۴9}J:m�vpE��I��:��g=6 �H�?x�сv2c#6�R4�m��7^5��ȟ�(0#:�r�`����ga�;�����_h_̂�q���3<F)Y��F׺)?E�͏O*���*#|1bp .W�j���Ք�F<c��䋸�Z��q{�l:�����~� $&o8%�i3J�!���6�/1v����qy/�3�S��h���#�}��1����oE	��`�"��7DK"� ���L���B~�B�H����t�e�A.�,��Jg'���ڊ�y����]��ie���i���_�Ǽ�2�̩t��������/�v\�yr�bM%�3Yֽ�=bw$���g����qSO���X�b�y$�@j����u��l�>ª����L3趚�������9��U�<C��1�\+|�S�e��e��D�b����ZI��ݧ�W�c'Ϩ��WBQ����Pwb��EW�LZc9����N'�C����8�#mH��.��&<f���%����a���6��%����b�֜[��%w^�,U��dg�nFB��=��+��g��L~�4��@M(0'���Ϣdi@?P����� �\xi��3(L�{�����ȗ
p�}��J��U߶'�xn��L�!�q�n�<�#t���!=���x�;f�8åS����&}�@A69��*�貘�U@�V��ĥ�4�y	ߨ�~%�7�VZѵ��gUZ����U�J��y} ��O�Ht�9��''��t������ �Tʴ�,�A���&lin���.�<m��E�)d�7��_��
U�S��4�,�e|w�g��S:���T(�j�Ο��K3T(��F~��W�CB���ąr�Zy��~^'�ؙ.)�8VC3���oY+�?�uj`���J7%Y��_A��d�C���GJV�����_�v�v��_hu��[w #��ў)}��6E�Ќ���^{�A9�����'/?#��1��˛G� ��:Ɛ-g�w���[�1��M᪬�d4ÄDx>��-Kc�G6��:��]�:>E���zH#v������C���ѡ'J�,�Vm1��޾�QY z�{f��/э�	16o��w�2��)�S߸t݈�ӧOQe��г�T/T')K\��9ȏ:;˅����6���P6ѷW���"H�����a��n	�7��2)�Յ:�X
o�����.FG���fMP��Db�o0����p�Y��	/ �[�L��d����n`9T���ȨZ�O�)��E��À����u0�Uc�J����al�9ݛ�*���g͍�^LG>
�׊N�D����C�X�ˏ������0'��I��n�B�欨�M��!��~J�]��3�ה�3�x</ik���/
elj�-LWW�9���R̈́:]��v0i�R*7ݜ��>F��&,!���x��蝼���.ξ��,�J����~�l��q(T_�h�����L�q�MQ������c�n_ߨJ~�>����l_�m����B�VF;�\D� &�^���`��n9�G��Vse���(*I��eJx��xȘ5��0��q3�����QA#�ȡ�!a��30!�:��2�E�5���Q���
���J�L@���p�T��ZO����/)��V=�b�|C`!=i���J�TjJ�9��wo��C4^�]�pX���as�����N�h2����&�-6��ڏ
]�:U�ѺYz��4�/���ם��iL�F|�E0��x�o�����AǷ��߉��t�Ek��������_�nz�����<٠�n/��jH�p�h7O>����s|����:���U�Gg��@VU�$2++q޵��8�����*��9Y�lo^��`R �V��W$Çw8T�maj�׈�O�ę��cś숤��+�F)���/yУ��U��B=Ї�'nNm�O*�mr) ��-�I�h���Wٞd�)�t<^)�����D=��6޵�e���M}V|[v�s̃�9XB1��3��/:��#��@h<���;���u,��W&z�9��Me����7�O���5�a�B�^�).Vd�>;�,�G�B��m噿CZ�P.퇩�L.�~�$",�i㎇��$�y�Є����Ԥ��1��r���S�b��zYO������?��S�xK�T�	�&��_9݆�2���=Y�tem7n2��W�Z@�p,g��q?I��,kNn��j%Ml�����f$W�xGje������(S�Y��Ѥ�<�=i����&�H&���_�(ux���_b�P���R���at���2lGb���-���q,���$4Z����7�!�u�h{�b�����c�$^�=�k���/�����qXN�;N�F Q�PrV(�ԁ�\��fT��]�����X���[�l	K�Hk��W�g,���M����\����nz�`}��B�oq\�|y}�	
�9ì�D�q�|�j^����Jn�QV���!��C�FTy���T���n��rmSi9_�K��EX4��6Q_3l���H�i/�#�9Ok�O�o<���� $BzT>���je�#1l�D��w�TE�7�����B`�c��f��i���}�9�[Y��%�>zs�$�Y��"}u*u�(���2l�5kR��RT��:��n%iw������r`Y�W��~��D����帴=&��wO�3!a�@g)�+n�.����)�%X��)c:{�@��F	
u�m�8֞��I^��zki��E��Gʢ)"�%}�=@��0�g�ɾV�P����,���Ț
O�(Ի��_8�{��\���a����vS�x�
�(_��-N3�)��A�|��ҽ���E�������K�r��$u��>L��Mo�^Î��_��cg̺�V�76'������m�"7�Tm&'�X���؎��^����ґa����}�*�1�戙�.����x�g���
�Š�d
6�����DF���$����Kcj��jS񠢱y<�4�����_(M���PG�(u�& x<��p�����n�w��|z$���u��[T�9i��^��&�y�Ȁ7Ri��;��mw��e63V�2��g#��� >V팛�RE�OkC�o��ȳcȪ��2ڹ����>X��[R�U!'Wɬ���;2��Հ~2
<��*c�g�r��R�L��� ���� �����@�<CA�ZƮt_Bn�DSOu��(�)��Jy��-_�\=�W�~B2��� j<-�')��z��9����yt�O�Q=D�D~�պ�ب
h�ϧ�o�SX=�-�uk*����@��o��p���<��UЪ�Ʀ4�fZ��G\�3�I� �1Ǻ{�����7,�Ҷ��L��=����G��N�5�
.˒�i�u���b�31���%��'��=�ɥ�k�S��J���N�y�rnPN��>��%cM{g�m������	H���3�"��<�,<�e��Et��]�0c����<n�"�_�4[�(�p�HTl�Q�*߃.�M���̲����̼�����4�O���QCt�*�Z���k�
2i�z����0��q�0��:|���g-v�8��+M�׮�l�`��^���?�f3i�LYRqL%�*��"�9���JMăJҦ�|���t���K����+W~��9��>�����b���G>I�&���T��ݚ_!c������ӆ��ew��=\{8I���jl[���E=;��\3f�W�?����[n�@/ l��D�YC�� ��A��H���D�P{�"��	4�����;t�ݟ�j&a���A�D��Y�x9U$�QQ��D?阱A1᡹�VkO&��#-|�O�D%2|b��L�?��Y��%�'�J���h�_�,�[���� _�ɡ0i$�7$�������^�DO/��J�;0�����T�h*���ߙٳ'��
G����%�
{�~��l�K�r�_�ezܳ8��J�<�S����J`[bݪQ�m���1����>Ն����*�5Dk.�%�i�f1�i(������ ���G#��]����c[`�*�U����[Ea�?:`��5Ate��'>�%S�y��Š.�;�I1-1�x�!���`��9O=;�[���:t4�#��NLŠ�s�������||���7|p��)�>۱�n��J�
�H&�1�+�������b Aw1E|����m@�����$^�2�hjK�ež��3�,!�(�)ҽ��/�ޛգ,����f�n�M_���[oG�)D��'"�r�{c�z9!�Dh�V��+�L�P���f"��|p3a���I1�i?�z�r%�B�0?>q���0Z�-�Jq�
��zi�vY�JÎ0F�¹�J:
݂ξ4I�f��9ҫ�VlX���h����p29t��3�S�>��MJ-�K��+�?x���N�=�rY�l�8�򖚖~V��^���(�5�����`]�,�6�r��c��Q��w����6J���L���k��H�<UǔiDk��+u��7AV�ru�$��,O@#$�FxrCu_W1����Lj�4�3�e��X�r���=2�c���/$S�c!������LkC��5f���a�ˤWi�Cg�>�)Ȍ/X���	���v� ��M�љ�9a{ET=ڴ�TS��uK*8B�/�`F���z��k3��"ZFf��6/��Ԗ��`>� ��$-J��
��H�5�L��9�QG���8��riU��=�T��Hq1)��_��8@)Q���S�Ks��
�Zk-.���v������ܴ���^?Tj���ԑ��b��R�D����,9(?j�&K�f�Y�],�7��5W��~��$�xL1Ў�<���]<j�9h�kE�]��{ηŔ��ʺ,8AT�eUW�˘����!�@`'8�pV�W��V�8w�9�p�]1�z
�v�+a.��>?	���I�v[�x���j���p�:ќñ�V́����89Z �q���N���HAzl�&�V5���V76���<D6�ۧ�AVu�Vx�}�����0Q���,}�R�iE#���k�������P^�o{�QS��I�aF%�k`w1+�w ��1��w�?�9��}���<���L�|�#�I_�kP�%�/�,X�ZI��AF�uX�}4�ؑ�����$Ǩ3�%�8����E�P�@�:�r�)n�0#4�QEM0!i��r�!6x���VHv�?!�����V{4�2������-�3����Z?��4��,n�K����a\UG򌎫\�7^��Ǵ
��\��jg]	�̿�ޖ�a��j�kT�D
�YtDR[y�L� `׻���ˬ���:g=��<�t#n�f�n,6��!ZU<l��?A����	M�yg��1��XV�������W@�?I��w���O�6!�g��g����2 ��}�V�?����S;b�����=�#7�`��%��@Z ���&�H3 ��b�~`��Y�l^ L%���)�e��8>+~Xtė��?��K���X�ܦ8�s���iћ������$��չ]��K�����甤R�W�YoJ9��QR2w��Vë ��]����
)}�-r^5�A��Z��-<�3�wIg4�ӏ��*���PKŉܗP���G,{7c���r0�PO���-���<��{x�T���N9\��XQ��XA�4{�;X>L8`�c��(��-`�_�A�]y���]]d�z��ܓ)�Q@-�9��7����8�v���b�j�v��Z]l��r�5c���h��s����`�{)t*��\����Qk���Dh��H81{b}��p����Q�ظ�b��3�^2�����+�=�
y4�y:UX���3|��&�*�-�6����T	��έAhP�4|�l�<f|D��y�pjq7bE���o��OW#2��$! �]�B"��r�h/v�!O���V��e(�7����%[{��#�Zƴ�:z�D%VM�t!�_�k?h�K��.+��G,$D��u���T�PeOi3�6RuG�������ė�
Nb��f;���,�g����>X$�w�`�f�)��+Wx �y��1�~��8	�Q �@ڗ\�c�z��d~Fr�4��塄������]��~� ��`�B�ղ���YpE�6��0�tgܠ�b7�'f0�8(	V��)֡?F��7��,h���d�!��:6�~�����ϊV��vl}3 �xO����4$t�)�}�^�k�w[VRv� �	�]z�kt\�P!h��??�p ?�k���K:�A
�:��;�cƄ��+�;Y�MME�*��-C��+�jX�?.j����W� 3���9��:%���g
��21`7���({ڒ^��1��.�����\7�-+�p@5�lY����-�E�p�� �L�ψ9N%�?�����L}�+��� 5��a+���ӧ<$���_KQ�m�SR�-����Ty����ϮĒ� ��+���#��4g+�t��c0�7��w��ո����C)�P/#���O� &)������(m���H·B�r�+g(�W�Z���Ī�H0�`�f�@W�ͭ��Y�w��~�%�}�.ĝX?��g�a�vNQ�X��T�i�'o���"H�G��!�(2r��3��p%�^����}q$l���YX㢰��T1�@���������%�#�2*�c��s��p���|R�H�Q�< mR���0s���I���D@!?���R.`;�n�c�v�ƞ���1"讲8E�r=��{���n8���s��5Fݨ��PK!���K��X�v�fъ�S�K�]-�����f��ʋ��^�.�i��屣�-��.+�i�橑�fT^��&��m��#�L��@�+h�=	m��_��2��p>cZ���x��8Qc��:��5i��#�V����v��%c�n)e\hpC'5?Rx��;��)�n�(>Y���k�����E}�A�i��<�h�#�&��kQ����9\@�`ac�Wq����r�f�y���H�R�J�n��`YK+2�3o���F�xH~�(����R7�/"җ�׿�v+��liC���2C"d^����x��Ȕe�0��(�T
 �\(2�(�"�ȶ����'O�@J̳��.�ǝ.#�vZ���=�!;-��9	�n�Ը�@?��p���wy�A�6���h�iґ��-��_w8\~��X���\G�vL%���1��孽 �yQł��VP�9���B�/z5�ʒ�ԉ�����;�/	�IT�YR�9E��Y�c�h�R��(�9uH�qJ�]�1� R5F6�A����^���V�T{dCT=k���D��#���~�Eq!�&���17��W�\��ғ���I#ίZ�����ǎ-=����WGѕ�G�,�0|)MIA9�닁at��� �K^9��<}�[�������T��&�0���ʆ���]"��g����0�_gM�����Ho�4o}I+2����R��Y�n��ji�8AR��-E�����nn��x����u�'��9�n+�X�̵636��j��A��E\�0�11�(��S�@f��{����|�_��&���F�YQf�O�(A��GѲ��-�=6`�Iq�:$�z�,c)\�<N)-�L���s���?�`o��>�K���%�g����Z�ՙ�1�$uۯS�J�&4�you֩��`R]갘�87�F��"+����L+5�Q㴤��(��I==��j�8l� }�+�;�p�;����i�16
��'�q�&��a���M����C4��<Xh�96��ځw��L�5�>ʒ�t1���{)��BuM`��Zsޅ<N
��yg>B��L�'H��$J����AA��r�~��g�ϔ�,��r���F�5�s�V<o!X�>`�$��`�~a�k��3BO�
����JE�X`���1����4���^�s]U�W\~e%!ZFqڐ�dLb�ŰJ���H������ek��jL�	�	,�N׮���K}�������Y�/Z�k����0ܲk�!���D���<�-֪3`���_86�^��Ɓ�Ɂ>����)������4�l0{�Q�����+�ۃ�?�-Zg��fV9_�2��w��� E�G2\(��3\�C���)=��t��	 ��&�[JD��w�X�o��`UVL�4��24j�=
Sށ{6rx��p�:����zo�{�J�[��Ĝ��Ҩ�.z�Z��j�I�v�j��s�0��G4xUz%��3��RUT2�cJ��e%c,��B�>Cֱ� e��r�MXh��#*;�at >�F���ݣZ�$��U�3��<��&h�g� ��`S�j ؟c�m$����,�wh������Q^P�����Ԃ�d�^��9��ʮ������Zda�Y�&�"rn�<rE�G=Adi?�@|�����_��#gY�p�9x�ݏR_y�p�[���j�>��ߗwJ�Y+���u�2��Mj�̥�(/��8*�{iC����M:�d�׃�Y�;���*?�������xo7�2�J��Na���p} `m��Ld	�O��GP�����N@i�����b�W�}�������/\̭%�%l!y�LltNDj,e׿xSYjUsx�~��g�ےc��t�'��%��z��v|�m�.I�Z�wL��w<��%���o��fH&�s�ъEh�͈�ʑ�z7�w�7M8{(��OQ%�a�+�ƶjv����
)[��>1�"[oF�3y|cFj�6Gm�+��q�[�P��4��&�2�@�E�b2M9�����81��tL�8W��:s��؋ĩ���,�����]b�����Z���f%�]B�j��}&���i�r�'��[\����om���١u�^����Y�4n�ϝ�4z��Q�k7]����;wAʛ�,�խ�u!�[��mH������#�`[��D�Hfy�Ic�+��.p�Ȍ+M�A;%�I.�Od-�:=\��H�>sY�w
Vu���B��)�YQ��6���<9�P:cxP�B��sx��?����ꔞ2�d6���,�������6��Vp�������<�)F3�o�Ub�*�k���D&�7#*��/��7ͤ�������������ؐ���u�����5-JF�{,߻�/1��0e��Ȭ�^ޚ�|�1U{���:n��i�R��۔:�#�+������`�Kl�����ˀ��>��"��͊ǫ��&�l8��͉��2�RK�/7~��,:I��"\>�c����G�I����D{��ʋ{�(FYg���>�^�ހNϕ(}�?�X
�w����@���zՓ����`(p�Ɨjgm�2Y����Y&+b/J|�GOhm��Z��O����Q�y��.y�(_qa�@aF��Y���0J�	�Cĩa���w� ��>F�4�l4d6�V�\E\�J��j؉DH ��~�^�2�Ef���,�(\:�r���|���%��;p��L>������e�h������S6�b�Af������wu�RJ�Lm�6n�@�����u:66�%Ը�Wf������iW�ޑF�����й�Ƃo���X�Fո�EF#��
a�T����!�o�~����E���2��T�
j�=�?�֘�'�OvƛcK�&B��(P�U���N��� ���$��\M��$b*Cy��m)�8���qD������kV��&��rZ�4!����0��7}�r��@��8�+j5n�wL��]�Kɫ`C���M�����7�J