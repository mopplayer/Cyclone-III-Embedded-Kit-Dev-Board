��/  S����3�c�ub��_NЀP���t�,ï�!U;�P{�g��Oj*�x �*�'|�N�Q]/]���8�APvq'xrE(�v3q���_�~(5����p�V���ه�7)�A�c���>S���.j1?�u�ƌ .�W��Gb�6M�[�B��#I`rV�qY�W��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��W�Q��L�Uт�X"��ؖ��1�O[�B���:��B�X]U%�n�g��5����͉�׃PuO�]��p�>6BD�d����MNM�è�%���*Mw��s?v5��P���]�]�$������[�>.��a��B,�g��Lð�p���f[����R��ix�b��B�?�o�r�hV��L^GR��zҀ�C揻r�K�\�>����q)u͞����m&�(��G�FY=�����ߝ�@�b`�*�{`�3�n ��K�31���G�g�r�1�Gvd{�t+C�X�J��\P뙏�lBO��9�����s`���e��q�h��c�?*y˨���HI��h�>��R?e�YExgU!�Z�C�>!�S����R�Vȼ��K�V�=<��A��%��[8ʔe���k��*H��ej�h���X�R�n�DY�%�zp]\�:]7����D5��K�2�nWl���zf�����*�9�K�� �Jv����`�A8,�ڂN"�E�� q��<�ɭ��"a�Wx�/�~��h��V��<Մ&֊*���/ w����c�
����p�C���37~�DvQ��vh��(Y,1M:b��8��t(�E�C1K��a���?tb�ܭ>ݿ�s9��\m��ڴ�s\����K��榟�um��9�4���X������u}�I�0�Х���c����g�/]wZ�g2�)�6N��Mywf@�'���G��T0�&�|�������&J	�k��v7���RYS����WY|��#��M�Ͱ�w�s�N�mP7l4\$��T��ս�g?b�j���1�c�>�u��\)q�(^׊F��_^�V�c���ئpJ��	��q��|��'���Ϸ}|L>�5B2;ӑ�"O�	���,`�d_��ͽ܋ߟ/��m��$�?
9��W.�'b��~]���:�hS��w�G�Ä���(ܣj�U۱l�ع���i\��d*��L�$�0�&vװ�\: I�_�I�'i(�*���k�Ls/��?���ޢ{��7����u��:`w��܋<V�`��b���/�/P�N"����켷@b�(�ߓa_Œ��d�PE����W����9��U3����T����|����y�u�B*�~ҋB����#n��3��}��j�����O��
�z*�w8�C�� u��2tG��NvEI9,����H-��p��@P�n,��ܞ*��ؤqj-ߖ(b6`5T�/-�~*h���9aJ��к����t�\
Z��<!�}��X/�2�]�B~¸��r�N��/��_e�{IgLO�Ռl�kH�@%?>�%A�L$�<=��_Y��)���]\4�!�����;�m���.�d��h7S���Fyo#C�*�oaO����d��+�e{NжM�,���3Ґhcl�8;z
=tl�|6��r�8����C����X�g`��;���,~�Y�D��ﲇ �������Fކ�	�"��TR�#Q^�Ҵ܋|Є)��\	ȣy&�Σ4�<c͛�ch��	�}��{)j����*a�,!��И�����k�G��������
p�d
h�����Z�Sb��U�Ń��{s��h�B~��Q�@Y����N҇i��(ۙ`T��4>Ɣ!X�ʬ�'�틍�^&��`�Y��ȡ���kP4��-ϰǟ��`�w�6:������T.3���8�s�q��P~Eж�Cp�� ��%wg�pn�@��4P�:��X���Xs̞���O�U8C|=S�ri���� �6�%��� �nڷ�v{���9D%A!@a�i#��\P�V�w[Y�UF�ݘ����'��-��MEm�����Mށ��Z�OT���}j6'�^��Du�j-�qQ�\�}$h�X�wdf\�)�:�Ժ�c_�5̹FƦ��y�:����/���G���Ff�Lp��q��~@e(gB�ʒMЙ���y�F��|�͟M��AQ@���I�U8����4�7�Ȓs�5��A[h�[P(h
vQ���:rVC������թ���ദ�$��`��id�	�!��}�X��ն�'~�TB�8�Uꡡ%������}	�;����<o����A���%����9�J�x��8��0ɰgy<�:j^�2���K"B�U�y��s���0��5Y�J��Y݋n��Հ}*(xׄS���cc9�SFv2��ډ�����?���;�ל���A��o���+JM����)#�L�5x'DA����i�_�gŐ�8m4� �X|ZrM��a�#ݼ�����Җ�C}v�P��،��H�B���Y�Sʄ�����8�T� �=�Z�����&.�!�H�N֌�E�����x�<O�����}�H�=L���@�"�K~��-,p�HO��*l��L}*�;H��9��m��d�c���ƪ��	pT�th�:�;���3+��#l�bjr�^gI��>��f��O|�tgW��R��ma4�$c���x�=�Nw�A01�O�E7�z*�F�N^�"81�����=�[�L0FTa&���눻d\z��.Yu��U��^B߲q�(0v��U)��Yj	U�ך�œ�Z;S�����q���=����u�l�҅��O�'j�Ԯ�4�M����K�OΨ�	���8�'��2�#��' "�y������F�֑Z��-���l9�kT%ߢ�SĈ�!j{�1�ZQ&���!~�s%|�������	b&�������b�DB֑]2��1��E�pO�#�g��A���"Bfȿ������=�o�S�V�Օ��@"�M�<��F�vߍk��}�w9𗽓X]���	[� S�fЦfn���k %L�F���&S��s���~�����I�p0��<���
��S�(7����9�H�Dע��~V��$)y�?�N,n��N^��u���B��j�!u�F'8�*�.�YMfJf0��ɕP?����@(���¾n#72WL·��l?A=.^�GJ>���yv���ú����~*���XF"�0�;	 ޝʆ��ގ �;�%=	&�����ۋV�����d>2��<z��P��ngʏ��iж�M�7*F7!J�.�Gӗ�m��%�&E{?ۻ�QGV��G���A�!7Ȣk��1�<�U�� E<�?����&ξr�b�P4.�t$���׻,�ɧ�*sS��b���O��:?��W�K��@`�_2��@�#>���n>hĲ����|�=�c!�X�/�[�γ�t|Z�հD�=��d͒?i�d�4�����N����N6�Ph���J��iv�`�Z~���{�\=[�-zؓ���^��I
����Q�#��fA����u�?��A �"��崍G���M�6D� �Qq����X|՘�+���A5��oI���jW���U�0�a��Px���2���y"��(�W+Sf��ތ78\9V��V:���f��s�o�T���`�����<�IZ��{`-W��о�� 8�"4�z�O6��17(g�	�����m2Z�̞b��eR/V���R���f����uNqPm؉�i-����[=�DPV	+�#
0
 H'�p��@yɂ�6��c�.�]P]����{�(�,t�4\���q ���e��x"�6B�������!����Qj�;?�iX�I���L�~���L�1� �|��q򹅃�}���jO�� ����c����
>uJ�t���`�3������;f��JRq}'#l��;BF���ˢ>s8���-Qq�B���vdB���y��L��􆄻�G{%�Ipـnse�����\XJI���m/2@�(Q?Oȣ0�K�<F�-{�D�=�'�4�?�R_�N/R큢��FFH2�I�R�E)u����j�BbK�_"���X ���ҡ�s��L��u�W��°k �i�ù%�Vv[�E&a�L{�\�<�rp��F
�AF�T��P�cq���.��*���_�L�DR�ʀ+���*'��m��4���B���qF����]H`}��@#��/h�H��l)��:�:�f��5��ҫg~�_A �oe:� �QyЮ�I�����zv��OlM5��*}%�Ll�(�ѵZŮ61r3"R����Q�F��`�����P�o�����k}4���nn�9^����\�?���-S��6�����(�-�g�$3���]G�x0��S��@Ğ �5m�l�<�p�=�VH�q�ޡ��m���>���zB�*C�0ņ���>�7��4-΃g���H'�,�}q��Q?t�;�Y7��bT��X��g�0����?���M�j�I�ꍂYp&="W^.�@9i���>tO���T��_�}�Z	A�D:����j^{�Rtb���	:Ƀl���2߮��	)����W-�7�CC{Z�󯑻�tvCM��L^�gJ�ۚS���G	DƺtGԧv,_l��Ycx���� ���.�Wu�Ie�6�ڱb���0����[��_5ga%�B�~�^��
��_ء�u�%vU,��EځQ��5/��g[��9���2�W���S %
���w� �C朦��2�m)m��OL�,�����-�Љ,G5y�nRx7gܳ�%~f׵̲�>�,�t������jIS>�4&���K��)�E�j�|��iy�Ga�[UL�d~� �K(n=���|�t���������p��Y�>������N9 ���>1:�k�{�:�����
�zC=:4� �OiUs�81�6� a�	�����d-���#LW�s"���qeW�i�1܏ft�[�������eCi\�s��\I(f�qM�Y���|�� {%BF��@|�:o�^wul�0���y�!V�
�����a@@a�g�'����1 �1Z��2�z�'�KM�kJj���">�3���NM�+��jO��è�g?�] �!�+g�Sw�K?�~��2�[+>e0����	h� �f�B �A���E��0��$����m!Uf�x���q��`���5�؋+j��^S�@�I�;��	�o�U�b$�.��zN�6&j$�h2*��ӿ��r�á��&�@�_T24��B7C/�^�)���0OAߥ�W 0�T�Fן�R�X5�R�a�����u�"���w����p��`���!�%�jD��L(e����H�ˠ_5.%������V3�q
�E�ʲ��2��R,�7��_H� .��X������Dh��K�	ZF2>����/p�&�Cf�z{5�T����`25[�����y:4	 ����,�������C�]��@��AE��=�(ed���c�.��ݼ0 ZM�'.#�_ h'�dN�7�W�������5�;���W�~f69C=͊��bJ��W�,�7���'��7?s@�EMG2��T��e�ϝT�3�I����c�=���[�,G�Zʆ䆮���>@̛�O���E�$���^y�v�e�"����Ѳ5+�(��7��Z�E��\��^x���܁,`'�Xb`����-�M3�A?�f���[֟����53�b7��|�t�<:ǁ+Oj6����B��;E���%.��vn �ˑ<���y����y��rfKR�AC������ e�F���DPn-4����=���N��RQ�W�⯗%�z�QPx����?�l}��A��Xq;X��ĜU���o�l��ͨ$� �ْ;�(�g5of��%:pI��}C]F���"[�8�j>�R��#3J�'�Qd\��^x��F��XP�0�ɭ�:�}�t	@��ԫ:@ͷP�9����[�!��2� 5�5�\�7��\����[4�C5�ֶm���O]sTÞ�%�5d"
�l��9��t_��M��`�'Z���^�Y�U����}�q?]���LA�� �f��6������3�<�A�"����oFb܎T��h��W���Ms/��X.��t��,�IꟖZ*�˼��R� XP^�i���όb�vk��Q�
հ�ҶcM���������%U����Đ,Żt(��(����K���0dJ��a�T����MC�oi:�ho��k����%�Z��;�mv
����Po�W{o!T&&Ar�I/�S�����;²C���$�F��ƪ��[!��`��]��]c�Z�GRYb�z�MO�sv�|S�w��uK6c�1�-���)���5��M�A����1e`���`���q����Pj]�5��q��w�����ߗ�ӿ5�rb�q)O�g��)��u���q��t�y��k/g��q�׀|ϒ�ԹSG�E צ��F�SO|�Ќ��N�li��!�Q��iR���k�� }�G@��=�	z5�9��MN����-NY�[����S�A�������R�	�ݪ{��c�7���8��N�9�[�P�0xE�BrL���YQ��^��؀b͕�<�襇e�[�PZ%�h��fӾ�{����O&
���A���f��jMĨl1NB�h�n�����L�֙�//�#N�!��#�g�V�f�!���dY�]��'�{��[~��;.~u�(έ�D��1�4�ǁ��y���V1�i&��h�zLQ�� WW�Ǧ"v�6M�(¯+%�D6�ϖ�8�├���)�󉰴� ��C���%���k�!��eD����@c��]�-�2K���+Y�̭}���C�p�꿗'��Uq~
əz���I����-^~	Ó�tɋ�"qJ���ʁ�Jp=E�R5Ϻ�ڀm+ӝ�_��My,�5�x� ���@)��s��ؔ��W�"B��͉����Ӥ�c��[rݛ�*��.���9O���[�	��t�`�����3�>m����j�r��&~�8�;��{���F�Wר|��9�?�UV>����wr�ԅ
-�T��Z����i����m|��*<H&�Y�U߭��i#9�ek�8��Y��x���B�v��d�`:�'�����rZ(P1fd�Z�N�����z��ٰç8Α~���S�Ŗ�c��uS�wU��������{�_^�A<y��2�mBIc���q ��Jx�	M���?Vy���윋t -�iՑ���ss�NhU�����o��r*l� (��1����j�XZT�⋐�+�����u�@1[���!�{�8����N}��x�3���pd�G�N�;����B�7��4t9.���	e�a-�=�z��ϋ����k?�^�v�䃑�̕i�-��p7(�F_]F���V��p񲋼ڶ���Fa�1O���ZN�uL13�4��������yd^��g��	~J3��D�U�6�'"�|ҏc�Эo�b�<����l��i`�1EC�B!WO��� � ���_B�Ι�n�:l�3[�R[��Ӫ�?Wd�5�����4]���%p��r��r�WY7�n���ŀ]qY[ǋ;�~r��{�Ic�1�.���cH�P+�`��(_��w�%�����$��/��c�Et7����c��V��rS_ZS��]|��7���̕S��7"�$,�S��LS����:LC���$�0��}M����y7S��b�^}T���@%�Q�T�]�u·e��$��e����]Ģ�}I�6�15� �i�c�I��q�d�Ѥ����I��ut˖����&�^�� u��k�z����� �5A���pM��\���?/�H��V$��RI���u�{�XV��i��L�-o�e<�V�HU,c���:D�Xe�Y�|�'��c��-���K�TA wV���Y�E��b롚���&��p�".)&I(��?y)K�J.�yQ�vq��tg�%��3w��TwF�`��{�ε\���C�41ʺ��q���UID�!����2Ju@����f%ؙ| �Ѵ���ە��ʬMC�x`�������������\��K�����b��~N��O	ܨ�g��=�km�oh�6�Zx!��*�ب��`2e��h�UKy='��[���Y��2�ɞ��;�|<����C闊���]�����+�Z!3pЂ#Q\��\�jX��a/�JL��W�q9l*�2Tn�KJ�%\����'�)ɒ�늨��ه]��0p����srN��F���4�^H��C�]f+��$a�xb��D���G~ot)������|k�6-��vZ4R~z�NS�SZ��ɪvd��]_���{���#�E�x~�~�}�����.h�c �
����nO0�E�HvB�6�Ͷ���
Z�g�7#6/�5���[��6�n�[)�~ɝ,�M-����/>�YC�'|��K�����Ix:n
L�f�
|��e�$w&��}�p��$zBj����$��æ6=���=��<Ds76-q~�M�ɠMI��v��c�}�L�y}�1���skYM�#�ǐ���#���,R�T�Ƣ��I3c[7'��q�S�����m&�J� 0�8��$�:@H ĺ��>�,k��������ʴ��Ӆg�yS�t�m6�B�V�� A�����^P^��(h����>�x����Z�հ��y�n�>��E�ka��C�~`36�@5��g�����txoq��{�~�q�K���)�P��r�;|r��|�[�`0^��-�����N.Ga��§�
�5�����s:}-7I�.%g��#��/N�,I��G�: s�r��A��Z*l,�+�8w0Zh�ԏu磜��oeW�����xw9z�����5*V��3������3c��OOzQ	|ɔ���(K�x'��ϳ�[�J�����mt�B�Q?i�2:�L�ez}CA�H
��X.|��b:m(W�!v������􍹴̖�.�mu�ױW �,"�3�A����qN��^���� +���	����q5P���_�~^4k!�<x�ҠmNu/�J��?W���18y��<��_h�:i+ >��t0��>]��;S7B?4��}hO����vb�2��6y~!a������a9r#Dϑ�H�"��q@P�>���7Y?R�BF�_]w�iB���/M(�t�LF�,�%���[Ei��&�]9ȫ����.f��w��b����ױ-ڎ����?!3)dk�|��	3î�3J�s��O�P�|�9�!3Ⱦ���ي�����oe���������hR�����cq9Y�QD
Q�^K'�d�He�I�w��/1W��6� �׽-%�IϹ�A����T��;Ff�aLR��JD��B�8�ܝ�!U��E��K~��c.�s��}��nmR1���bϰ�����!���Yb�ôے_�PoB��K{FM��Ds��Ƞ���vy��c�㠂���p�c��y�����!䞿�g�=+E>�e�H����qj��w���v�d!pI'E�P/~ٍ�,Ļ�z����-� )�Ce΍�Y��,b�:U]u���d�'��8�7,����	��G��w������5W�`��O��ۊ�"���(��l��U��^�ͥ�?C���H���.B{ῥp��as�L�9���>|���9�ժßޞ��|��:vtb/��@��;����d(;�/&���,��iU��� UK<}�c@ac� �7^��Ҝ��̕KR���7�;�3�3\3������Vʺv?��r�!B>�������&l��U�N3�����a'Io���.�&n�$@,")bG���ˊ@,��=,�?�.)�;����$�}	q��% f%t���r�U��}I��ʿK]:��V}z�����J<*� �L_�x;q���I����$<N� ����,{�EB��U�?c`��T8i�^����P+�mB��#6	 �6q1��~���h^\����|�\�	%��G�@H�]��X��UAG0��1N�O�����[y�X�ؗ�v	�p?�.��5�(,���-��.-�F3�����t���"΋����?��W8t��\�K���"1�Ո�9`,?�h��*h�eEn�F��N|����I�B�*%P�b2� 4�<ؖ_h��վxẌ�!�ͱ�E�k���� ֖o�!��\�6��ke��rJ�l�:��/���l���::�lC0܋F$�F�s@��7aߩ�xMQnfZ��]E��AʏC��კ�L�`'��r�6;,G�P����\�e˺e�Z�#��vkzxD�D�\�wz�I�OJzn���A�~HnxXY��@�+Zp��7W�?ŝ��<�TfcgTզ�W���Pw� J��-|;���DW�b�?n������0 NUKɍ�G�]:�ՇTm1y���%۷�y��Txa�����Uc���.��5�:Ȳ.�OP�� ���k7�I51�c̑i�)ȟ�[�d��M�Bz���<E3��D�'5A|B̌��y���σ���<��e��S�T+����v.��ɿ����B�}����ث����	��5(��hlglZ�/(���_��� )��2t�0����)̹V�\��'�* 8�f�be`}��������ER~����Z乱�^�S������F�M�����n">��а��{���W���O���&�8,���#��sw0���s�7��#+n�
]W>��n�����lě!P� �_���G�r�����������e#�s���H龅�u �.��:Fvt,���㯠����-�=a����R�	�G�W������U���<��k���@/VB�ɠ/d?^���h�̈́��ۯ��ɦ<�I4�02l��y�Fޣ�����ֵwi@7�D�w�T��Vq�u�.ø�{"�L�qM[�ł:�_�RĒ�@3�$j�!��ƾ��ΤM��<}�E���������ϖ��P��I9nMS%-�uv����ȫQ�&���4�$҆�4�d�c���ӹH� π��9�.�VΙ������A.w�Ijta~d	$7=1����>T3R��\[Y`���5>���L�M+¤\]T��t��k��?��u^a,L9q�����'�����5�VO�v�'J/�i��{m)�N�x�� ���p�4f�Ϙ�@���pk-�-����y�5̒>A�0�	����Ɩ��VuH��������VI�E�6O�s5Ay�0��铊Z��#\љ'h���W�j;F�\;nx׉-�l�?�	���J*.T�X�4������g�<T�M���E߇�Y��(�Nl������9/��u�t�ݲU	��ې�s�-6gEhb��A
?�^�1�Pt|&w/T��ә��vB0^ݧneP!/���� ^�z�Z!�����I*J����Ҋ���uN�ƀ9i-�:m�3���X��~���QYI�Z
�cP!}��"?��y�N$�)]���Fe{�7���B������'F�����Ŕ�(L����L���H��1G-�e�z��+j��@%���U��������.�Ce$�p�7�0�U��co?HYm�|��-<� #��=��kr[�n`�F�,��J���p`!V��-n���{(%�Uz
�-���\^�EP&p�ƽ���+p��RZQG7Ԫ�&�!�~'ڄ4���e�K�O)iG|�fI;�b5�f#��Ň7�^�1��k���ԁ)�a���8��A�b��;��s�Dֆ��Dy�Xօ��ĺ=��	2�z��r�D�E>�a����נ�Ns<"��۫�2�o��{�Mȫ6v���ן%������8ǿ����M�}'�x�rC��`�&��;����
��ӂ�&�V��Rj	"���dD�����4��s+�\Vkh��%/U	����VB�N�_4��uV/Ԗ�M$�ߵ��q�8XDK�A>�}2*��͂�֦5)J��$�'��52�:x7��X5u=�e��Թ!�ԧ�����m,��FH�Vt�|M�+�����Au��2�'b�.�~o�H��ܡ�����N�E������Gv��^��}0�uT3�wM��sIQ�,&=�U�jd�&�o3���R��=�T��Ɛ��f��{[0E&_24��'>��|�u��Ȇ^�q�0�A�g�:�eKJ ���p�9�+bv�)gV���T
�8ە��Q ��.7�p
�Ya�OWa6���m+�O��� ���{	�����-���,�rZ��f���ϸC�.6�r��u�����_��@mO� 7x&R�6yS��Hr�?̥z������uyv
�ֲ 9�d��;6�������|�,#q"��2���H�({�����PQ{�������9��5KD�p��	�Ȼޛ� �H�H`,��X�8����rPx� �ʧB33hY�W=?�Cj������m��h���7Ā�fv�������߯R�>f��S�[�u����4�_0Ƹ�M|8l�������~3���,�qص�/d�E#���V%�����g�7`�=����ڴ�좁��t^�ѹ��4��L�tcu��6;����ɒ�L��<�N'����U]�ސ��j��p�U���Vݧ�Ke���d�]��D8��h���+�B���~	 �G���$�����!�mgV{�298m�6�����I���x�Üh���E|��soy�]83�}hac���~#ʪ�������v������ˆ�k�nF���_�!7�~I�hG�6��_���wU���X^�D_ڙ��]�#�gh����n�hv۵�9������2���gul��!��$���j'
dad�s�z}�V���Lr�U��f��̗wx=�ϐ���a��K�W ��D߁W�.X�e���%��q@�K�R�&�5�+x�З�eԺ~��j�`1�F\ʉ��	a�&\	�dÉ�_6��I�{b��4b��3w���0k/���7),AY j��������/���2s��_�֎�2r�`=�?���-:U���I]SBd���6�AqT��[<��o�.��W!���I���V���-�]3�(@JKU�KȟW/Z��� @�V$?p-%f��6Qf�4_��Kl?v-����Q�L�q�'�e������T�Y���.(�.�opY���t%�U�I�z��c���Eի��u[�a\�R�8���^T9�u~"8炱�&S���W/���QK{r�"��E\H������ "�f$Gn�B�!D�T�6�͋~�#����H����L}Gũ�'%I��&p;L��
䀏�e^o�]��M�#A?e	s �Q�����WzفUn�l5��]00���� �h�_b�7y�S�x]E�#h��ݡٵ� 
}��
�Ԭx��&���� ']�C7e��3C���.�x��_
�R��[ �M���#k����A�����S~\W���j_E����x�J͘K���a�V5������%/b�"���L�vaJ��:�*��Yqy�����H8�ڍ�FU5o*��{����C[��@n�k��1���ل����v�Oފ���*�'y>U:Sz���#�*�2������������0�.sA�3��*>4�2L,�7���ҋ	ɰ?�TʹU�h�����ȍv@]�5ʣ��-� ����� 	#�n[?�Q���"�t2~�Zǿ$�g%�d��/ ��w&V
�&�B~�O�ik_O/�ڄ�Ʌe{�`�f������:���-���a)��<yL�x/EN~����r��lG�F��g��0��TA2NK|ckn�/4�\�쨖�}��@����7i��F�Z#�-�ῤxVŕ]��,'��Ǿ�o7��Nѱ$��H�Ü����<�"�2|��.)~>����k�ڼ]�_�RU<O�����$���!�U����k�k� �:�t���]�#H�qd=�jY������>����E���O@D�A6�<he�������y�-��=ơ�h�~�ۢ�c��w����>vC[pS깍��ly�my������W2�R��L�;�+��Y�(W����j",UZ�<>d�O�Z�}�~4��yT�`�v��)��xQ��I	]�x�_�?��vA6����]%:l�i�P9��4n�3�8U�'?8�?�ܰ:�WD�_l�T��S�a?� ��Fn�%<�66������=�m:��,2�Y�H�����چ���~��'Wp�L h'�"v%��nn2��s�؝
�
�fJ%7●I�wY��OcC'�l��1Ʋ�L�c�0Ng��f��5:�~����H��1x�,h6�jp�	]0���w0g�B����|@�����@�=򪡵{�����QWSzn��ᙪ��)R��uݚ��[�)�U�|q��nTl4[��ǂo��4��8/+�OŐL�jtR�%{�ɜ�Iˁ!��)�k8+�Q�e�2���?�v���i,��p�x�BuF3�9���6�-���{�uО�o�IZ�V��V^��߄�y
��W�]�m��Nq�
ġ����uA��24�pԾG�ɴL&-^�T���ӯ�D�#{�ǈ��H-;ʸE����S� ��$Q���b�CA�[��U>�,M�>W�zd�y�[N'�g� �4"	0P��b8%�ִU!���E)W�CL�O>��L��9ꉦ�wh���})�ɛ�D��sY��\��C��=�U��N�<;��y$�x8nY�XJ%�EYp�֞y�Y���/ɜ�^��_�
��4��C�$��^F�3���U3���~�+/l^��)��[�q�&vXlV�v������/b�5p�ѕ�U�����i�H��Hr�3]�:b[J(�d��;v����_���P�t��焺s���9���q�������r`V}��$g�]j��K��i:0혚r���rh��oN�k���r~Ṟ�!�V���3�bQc(�R �=�Tʌ�}Eo����$��mnfЦy��	�Q�9,��N$���*��Ya�0���m�:\�����/3�Q�. �t�<����M85^6�ה��Նpf�����z�����#dA$$�����h�	p˩��N���V^qrъN�v��a��C/f�/�d���{��W�S��a�!��sm7�E�&�F�S �h����`	���ZZaoj^���K��t\[ 	G�]�p���� sS!�������JO�X�[9ZC����`Hprɓ��IR��cd�����yC�c����#��U��-�ƻ-I4AdB�oS�Q1F���eE�[����忝%vG�-^ʗ�����kg�ނܥ�3��F�-�g�ޮKd��F���{�|����a��-���hLO4�sB�o��d�t���_E�~2 X48!�� φl�o��֋9C���:�$��V�	ц�<�E�8���`�lmB[��.(̊����9���Qo({���^�ü��w�,H_��5c��2���r:��������j�
@�ޮ�1�^��$����U+�k�N�`�ٳ��g�18{yb@���]|���"�D��P���u7X��H���8S�a�r����a(R�S&���g�E|T��|���H�?�6ח���9M��������7pD�*�W�� �p���S��G5��+�xԝG��m�Ϥ(?5+y{_0�Q�
#�m�d��OK%����v�}s.g[~Q(��n�,�@�:q���j�)Z����q�X<����FQ�X�a̫iZj�D6�jWf�� �m���r�?"��K��"b���uW��&ߺ-Y�CrJC�T0��A�%܍��¼�~�5��j_��`m� �`���O�m�� Q��]]��r�4�����e��K�A��Lp�$�rp;d2�hG/B���L�����}"�U��*�;�1��#M��1W�Mΰ��+����+��x(�2	5r�B��.��qs_�7���R�86��7�%�;C�V0�h���|	d'9r�I�Ϧ����΅��l6:�p�r��)��?��/���M�%nO�T�rWJılAd�xE4�K����Y+��%EQ]-���m�(	8?�ł� -�lP6�+ˈ�5�JD=�!<���}D.���(w�N���@��=��J�-��s+��Vd��qOb�Cʒ��-R�����<Ɨ�����50�3�g�J����9�YX$?��?��vc�w���Ҝ?��u�۲`=���'u[s���ο���`Vjw�\Ye8�(UB!��Ij���Q�^ ˳������K��>��$��ěPq8�I�B+�j�*�X~�4iH�ʔ���	=�1)��CF �#Fc8
u2��%%��H?y	��]�v�H�z$���f����!#����>����3����/�`Wo�;x_��o���q2YH�������<���W�
��_�NϷ�ڂԣ/��%����Oka���n�BV�BC�ԉ�����z�q��gD.��^�U^�E}*�=�K� �8n$Hǫ�j���c�}��&20������֙gY�k~ m������E� |@P�*�n\!�-*��)�4�9�	�ek�����l�|��V;�v�]`� ����g��R�=:�S�	�Wˇ���a1��<�5af�ĝ<X�s"��TO�Q qB�0_mf�T���~=�ag�$�h�S��
8�0R�Gw�х�=a���j���AAY��S��I{���x����� �Bq�P�ȯ��TG������P�tâ��I�;?*LF����o\]a�$zaPm��v@0a ��v_TfҪz��k�\ �c�J@�&Э�j���|b�J�L�G�}^a��PE	x�V��.��á�W�����h
k�즥�sh,�,�<xY4iE���Ǭ�6�Z'�_ms�w(aZ�t��5�I�jܨ�>���O��Ԗ9Ta���� q%�����<B�)�� mZǃ�u����r�W�kU��EQ1��Ia����xo�I�E��!�vb좼nQDZX�)e�{ޯ]��3\����%c��$iKP��]��k�Wˇ|��7��:t��č��#�X	ܼj*�Y`�_��i�\#��Hɩ#�e��^H5j�I�_�}V�����m�\s��񃱝E�y���c�á��PՔH0��f��TF�kjY�
&w� ��`�Z�(�����L<�]!��o�E��̝K����*�Bt�	�bT���Ŝ�=�kl���s^Gh޻�Q��pT���R�M�!jdF(�pם	Jޡ?�V]s?[i)tz�$�q@�|�s4�q�s�Nw봋`��j��^Z(f��pSQ�y�A�C�|�<�����ETڢ"V�rD�Փa,��ڤpB3<�Q�u��HŨ�N�n��{!^��t��9͠y�y5��:�	��K%���l#��Q��f�nI�A:*,D_N��Wa�
�h���9���
��#�&�\)
tr��0�m֕�`kw&K�a�a^ U��p-�2,�������Y359��PM��v��a�<S�k�;DΏ�eh�T{P$�hjw�i���!��T��Q�k)����x��������7%ť�"��2����!�O]H�6�^���F4�i�(��8�W��=�L�r���V�P��_��_L���R��Yeح��P�s��� ގT�I��Z���>R��9e)���߼IL*#c��f�O֗��*?_�e��:�� 6nȕ��yB~�ޅ]p���D�xt�܍Q�9�1�L�Z��2����ǅ.�#���"�ˮ��x�&�]MTY�:'� ���"̿��X�(Y���4���/���x��y^��K.7P�vN'�l.Q{P�0�$~�s㏴!w���ݴ9���uX����p��A�D-^yV���L��/�ߙ\N$��v�F��Gn���H��[��I���I�$#�����6�b��a��q �B������-��-sCQ�=�gz�0��e�I2o_( f�2	1��-���Ҿ�}M2�;���j��43�B�b�����5O_0ʙ�����Em!dp����r}�󞱎t�r^� $�3yA2���'��ۑ#ږ��C9�'��&���\��Л7/��6�=�=O;)��*A�cF/p����;E,]�].�	��}�����"4�ʖR���Js1o��j�^��I(��8�PY�	�n^[�`����x���Nҿȹ�Ĳ�8��y�_�&%|��Q�}
��f�I����/t`�|=�Cw]��e3�Z׫x�N��;�kvclH)n n�|ڙ�#���2κ9y����T�e������m��HΰW���&�����:���8 �#ҳA@������X=��jE�x�S%;,:#_w�'d���(�5LS�瑩����Z�<�H�d�8&h�M�D��ͬ1�}yR��/Q6�U��~j�{p�$�O�-i�fS�j�&��9�k׊|�ɓ��Z8�7��a[6y-�dL�^��wֈ\�Ԗ�;_�9�O�2g2ך>x���@��-#��8�n����0|_-�C!�XH!/�{!���Jm�(k��l��kR�XTG�}9���ˋ�����A;�/۰�9�ܱ��� yŽ�IY���]:ת�=�&pa�a�1B(Ks�+�jJ�Dur��������hw��Z�-�ֹ̐X�2����Y���.wP7}���Qꊀl]�N����:��\	I:����|���*Wl���<�-�⶙���$����j�ٸQN�j�����:�XP2$���aR��<�� na��T-MNd,-P�c���6"�z��6ϊ%�a٦��5�����ǕU�A{�U�T��Ľk���1OaL��r!�M�vnُ�=i� ���%�k<r���2�o�n7�>��)ȷ��N�;��؝���|Ҫ�Y�A'\�0�	7W�H:vC�1X���ThX�j�ҡ�y�����v�E��֛�n��]���w�
�X�3�_�G>���;>���"�R�&e�R��8!�>9nO(=ilC�r���~l�D�����`�K��(�C�^�[�����J p{���� ��\aQ�'�U_ߨۣ�]s�t�_M�)ٽ{��e�����v�=ُ������l�)�s�'[���<j��3ke��U��y͹�A��A�	�������F���5|Q:�:IC��Y���$�Yk��6J�R~E��Ĩ_z*x��_ZI�+"a��݆)�~>�ѳ���b�:����O]�f��MByT�%=s�ub��m�qF㥨8�9}H� ��u��� E���Pf�>������3ɦ�Y}d��y5��;.��Ҿh��O�6T�\���6km/D>`7����QS��@;�
z�b�u�����bا.[�
�n6=�
Z8i]bX��Bۦ=9i�h�/G����xN*����d���wU�����!?��𠺹����DZ����b7�$]5�E�DJ:j�H~��nk�����}�?�� �1K����ؘ���z�J^g�+�.�Oۨ��uq�d���z^���}V5�1?��7K#��CKb�4�N�r�n�F�
8Jj{Ж�t�U`)��[� �H|��k;Q �����G���k�r�e�#��z'��5���
LKvBM�@�w�Z��]j�ͼb���;�1�7S ��l%d�1�������2�(�W�c �`Y�J���m�h��&R�X�2j�n6J�Tv=�O�ͭBf���5��Ȼ��؛���:�pR���p �j�L�~䓺����P�n̖�Gt1��J�a"���hx�5��]݉D����m�Hg������M�﷨G�jg4u3ǯ���v��R�����Q'v:��t;:�Z�/�P�(�H>���.윻�ʛƹ��'-E>1�ܵTkrtD��RlxM3�Ą1Re�⩷������Vk����o���i��d{����Z>z_�&J,W��5�yф�<A����f^(�O�՟�⬿����عf�s,a��O�����{�a\5<�+Rn!�2%dˏU��	F�o ������Rxӭ�3gBʨ���I$%Ѕ��oۦɜ��R/�7�����������)W����=y��l��Qa,����U��YFuH;�)Zk�>�p�'��}Z��9[lj^OO|&18�Ն ^:��%m�؍�3iu���i'����7D�����NZ��8?�澒X�z"����N�|t^	k���$@@��/nBQ[֟	b��}Ď{;��o�GR{w�w�4� L鷵�wV'B�?�9bOC5��7Cӹ��?�r�DP�+^���g�zѽ�`���W�c���3�%�.֤�	/�0�H�ǥ�����K}�����Q7�����7V�~�s�
�܈L+��<�}	/���� :��{2��L��P���1�W��Q>`p�P���K��Rn��7���INH��6��L��DGF�y����8�Ǐ-\��+P�[�T>���$p�u����k/@��T&'x�z��".�莜z����Q�_�	*�8�
�������c�#\rV15DǷ�e�bj��8U�أ����5�>xiO�A���<"���e!܊�O�'q#_�~�T�6X�~���(�W]�{�Tz�����uԤ錔�UtC��k�:l�Ŧe��3���JoH��Ӈ.yp�6}DěqE�NK�0=�l�~y�kf�0�v&�`��I	w�̴��z'H�F� �/�gା�/pLdg�����h����wa,�2F�07�,8��rx�<��CX��� �*1K�h�╷�6@�JOJ�_�5�DBH$�� ��q�P�r�m�0/�e��y��+��=E�S5{^�i����X|7��'��J���@����e�o�ʈ{I����F�~�<�Zs�?u�MT�Z)��vr>P���+Ȁw��k�>��$8{>�}�θ�C�Đ�(�M1kå��l��.�b��P�〪�"�	��$���H����}8�i�\�??i|mU�#���J���DT>����J�Q�����Ii+�`V�E��#$TO��鬛�fz�]��l���X+ǈA���~S)�j���J�P��.�1o}齭郲D�q^Z@N�Rj�u�qy�.g��s�e'V�g0�aǜ,}ڍ�p͠rwwޯl@��W�^O`����t,dtF�����F\ϟ�ޥ���)��qM&�Ʉ�3F�2��>�{�\�z8����Mʣ���o�O�&S��'-���PT?��aB�/0a3��������A)�d�Jh�z]��uRo�qJ��l�;%��@3
`�*���2ύy�"���P�H�<C�:� ?��}}���.�6���1�L6�$L2��E�r�H��d���xL��%���7�1��9����L���$_�!�\��������V�DQ?��^����R��z '&��e�C�x��jb�tHc����c���LuS���,J��V2\X��འM�7d��C2�%�J�O+-�� T.y�����GH?j�4����~la�x��y����Z�_�c(
cG��	�8�����Bee�Xc)8���!B��O��Y�Ŏ�hD\/�0��������Gժ��_����k��\��{E�ߛ�T�ߝ�a�~�K����Se�dA^�$��;�NAX�>�`IyA�Ύ;c��#�0���d$*K������v�g6�Q�A�ti7
�
���mE�7����t�����a<!��KC]d�V�U�1������`(���Ѯ��+�����q��r�@WJ!�`���]�d��k4��۴����gw�x n���S���&��퇁Pt���k28���WmL��uÔ'3.n�*.>���Q]0�`�g_)�
5��8O��A�moǆ�����U�a�,n�O�c��� 믈H8���\�!�J��Oy�\�/��ą �0/P%vE���;xW7K�0�GE�����3�����fa�
g� �Bٲ��n����B�T"�k-#��pD���pߘ�L؉�����8E�i�Q+G�F]ա)"
��@ZM��:O��D�W[��<|ߎ~HT@��f?�7W��_!�AD"�=p/�!Y�2�ʊ%�rָ���@�i���ԅ+L����}nU��jK8e��aI��Ǩ:&����a���:\]r��C��C5B�f����Z-�{K�Hy	���4���ǟ�q�{��v�gj{�����5̡fb~X�Q<1y�������v�d�K��d��\�8�2(�a r=!9EN^$W"K'�~G�m�q�=��6��uT��Д����� ��
:.1��-Tƃd:�D����N���Xb����!�t�5�9ɯ�9�ׯjNUt�P�X0╞�dz0��u�oB�BI��p���}���^+���VY���
��F�;��zY�$;�BZ�m�'��d���������{�7R0��ft�p ���ڨl�[�+�е�ZT�6��8\	o�
=��*���� E����逓{���>"�u/��q��;m�B�u���r�k�J$
�1�\�GB��g��.31ճK�{�����_1��c�Z�:ȒI�����dz[��={���h�NG>�~]�p(r��plG�T�K�C"��N�����#F8
>Aw�g�=Sc�hۿC��HBW�Mp^��P82a�O�� W�U&�k��V�")�J)s�#��Yr�.�yc�dԟ�_�w7{]�<a��	��Z��`�=a*D���ݬ��^��{��UQd�FB����l~�4M�d����9�����Ž~�QC���G�������sj���k-e��{��e��q�|Ȏ�DwkE�F����	i�$�>��&��6!�p�F@��GlR$�;R��X����O���/��!��//Ym�%U0���t��Q*�W�������MI�1�/,��6���u�_��"��.��K���{
��u�����?�:R/��3�g�����e��=�O���}S��;�s�/O;�dtk`��w�:��m�TV�m����$NŰ�C}�.��${ј< nI��M�2c����o=�Q���aÈ�m_4ř <�������Y�D�<+�~���A�+ ��:x6���Ɩ����kᓦ�/~e���E!�qI��e��C}*��à:�t&n�֝N"�W3�Z١�����5</h��(ac���r ��iB�1��)3?�6����A��u���=%��&�C��������P^���V�D��,4�� ��B�k����]� )1s��8�� �d�����$����W��|�y)w�'�r˥����+{���ywr�Iɛ�&͕�@�Z�=m�����5�1K�ί��L�in1��DKa(^�
ġ�%�`��և}��u�XE����@��"k_)�x��+�jҨ͌g���"A�����񓁫�o'ҝ�a.�ܽ�j&�
�x�\]�i&��_�6�)�1QrY��Sc��	uEZ2������ �Y��'W=���#':��yT�{z�S�id�-ӗ�~�{���a�l���-GQF[���RL�M�V�5�]y�L �XO �x�;�^҇��9�2�B!2��(o@�|� �P[~e)��Ǵ	u����v)9=!�X�͂�s/��8�÷K����Hǫ�%�&֎�Z��"�+�TJCݖ�	 N����u~���P�O@��!=��Z�Ceth��� n$'R����W]/�!I
8i0����Tr�F�m�yJ��n$��������*�0l�{�(yt�G�k�v����6«=�z3ԣ1�x���h���Si`���&p^�LuM�#��4� jq$������Ͽ�i	��R���۔8�:�#��Ym���z�$��R�"%mO�?��ԝ*h"��L��E���B;줔�4:��i����~�i�;�rDJ� ���#�L���v�r��V^��^��.���cd�x=�v��G��R�,`|UOq��!Ȋ�6�QZ��*�0�$��op�=۶eQ*��P�� �|��������H���Wh#����XwO�c2ՐBj���K8�R{+p0�9ީl����8�R�j����GQ��!L�Zpr��`bu���#ߒ4��Ԧ�\l��|<7"|:Sb4F�����bϔ����31�gKVp�V�/�\����UM����_6v���]H���L��BV��� 5��a?��ʖ��yh(#�|<�lo�S��O�l.r��HD ɰ`��7L�.��H��zOW&��+	Q�S��S�؞^��"����{,.���	/#ǔO6�K�	�y�4���w�>@jA���N��,��;��;��S $"�,j���^kb��zpT��|�g���֚�t-Y�ˉ�4 0��:��3;�Ev��.�C^V��U�rB�����L��=|��x�2= z^7D��}0�|Lf�	�]�&iP��������a(�6y�/�n�F�E�|�! �$.�.��62r�*s�8
�m�V�ܞsXF$�b���� ���h�y5�s�;n&V�:�Dwk"8~�/c�BZ$�x�+���4����t�\QjE[��4�`)G���*DQ�\J��[a:v-�o�e!x"6���v�x�z����L"��K�([����g-S��H�%e���6�10���'�6�.�ͩ���jk��pCp����,��+C{�Y?�o[J���-�'�Lߴ��H_����4���{�X8��u{�BF�o��%�*vc�����!���:������*��C��ց��
�{L:$*%�nY}c�^���B�M/���3��)"��rB�j���jw"�s0���Ch���=��Kl���F��/�_"p���
�ǥ�.��R!�}ӣnT�MI��N�	�;G��ދb���$/u���|���qʏ*wǗ&������J$��X� ��d�9�w����60���mCJq� ��[MG3���az=:?�.�B���e��M�U(�VP����x
CZ�jɐͥԋ�Z���BvGM$�Ơ�]�˰9�g�������Wp�K� ���OP��S�:��,S{w�<�&v���m##�!�h���Kxbް@yBׁ�S��n�E#����Z��#�oFV�5�DN!/|�7Z���H���N�����9�eU�&�?�i2'���:���~��"Ncؾʹ��$�A�8�����N�~��ZW�rtq�-/��J���7�f_8?��fࡡ*( ���*��K*7J*+�9��� n��	Рۿ���K:vT%O���Q�l9�ޯ����3���%?��,/��Y?�]�?ΠK�bڎ�5�՞'.xqd���?�}�e��M����av�	�@� ���^V0ڶ-�s�u�_a��G1p���ĹG����y8W0���?�k������T;� M0��#�T�̩E@~�
f'�\�Y��N���_`��V�T�,.����{��ȥ����Q�c�A��K'3�8j��,��[���]��vz��k	j�;�R��3�%�Q���'�H��b�Z��c��>��v����i���;|��m�We�08S|X7t�T��=}9 F}�dr��zt4I���������%��f���~��h#UV���ª��5g+�R�y�3�'�8D�l�u����3Cѕ�ɄeF�\��1Z�B`������9�tZ���n�;ۧ�g��g�gӺ�TA�se�?����7�l�[�e�� ����Gu�P��VHlG�D
�D�A;�{�l�Rj��~�@�L��ի����i�1ϻ+ۃI7+��m���͋C��p����m7��/���z�|��d��~-�L�Q�9�!å�y��L�s<��W{ش��RK�:`O�ĥ�?�.�<������oc�$���ܜ�R��w�Lv�mR�$�� �v:�K��	T8���#�k�k�����p�-��p�%�g�!"gA�v�i V���j�id��M��� '��1�R���Z�Yw,�xyM&�H���Y�.�s2_�^������8�'
�we�:-wrbS�7rӀc�ךNm�PjC���=%Z]#<��&�ǃQh�v�8KP��ll/g�X����w�ҙ��o� ��£�a2P\i ��|�صA�5���7U�ED_�U�c �\_�``*��i�\7s�И��.���B�<�8d��t������S������`�A�۷@d�xϷ57�
P�yZ�H���w��u���_�̌їT�$kI�ˉE%t:��.���Q��=�Ŝ�t��X_���p�@�$(v3H�bT�?[	�C�<{�+l�0.`Ԋ�C��I�����̑ 3f�I�>x�Y���h���=�"����X�3l���=�=���ed�H�s6��?EjI��	�c��ò�5%>�/���~a������t�M��+�ra����Q|?D�	p~tkn����h8��s���}݂�[��1����8��ֶy�v�^�G�,{�K�y�'���(;Hӂ�y��Z�k�B�*��ڔ���.���.����";>�!,Xۂ��ȟ�Z%�'f���m*4���8g��FQz�7��p��]f<^	�a���vTV9�#�m"�����Q"T��I/�ǖg��VCFK���}��#ӈ��ō;����?��f�<�gJ�}�ڢ�d��!�"RPtI �y+p4ف�&���8�����`l�*bBT	P�\�L̎&��{#�������h2��gr�[�&��F�?�r�6�E��;�wKa�;XV2<Q���ǣ(��A;@$� �,��DR����Xc�oM�Q�րe�#7��M��YБrQ~V��$[��5,�`m�6Z��ިɻA/&$�Q/z��N���mv�7ʚ�ȿ��{���?z���~۩��N�����/�v1.ޒu��l�8cn�C�{:���I:��l"�4��As�O��j���m��s��~�(��vR���#��jXJ�nTr;��i���A|��ב�9��g�� ��<mrf�t)���)�EC��?w��q�'�*�̼�3�m��$S�JN%�ɑi[��(	�B�~Wi;�-�ܨ�6��㓙��jhN��H ;�9n6�9唟��$̳-o�Ho�df.Oa�j{[��H.��O�t)�E��p�7��8T��杗v�+��ۛ������`���D��p����x���#���j���'	H�c�,�)�^�Z$�rg��@ h�JH�8S����$m.,�/7i�f%<�{�ۤ��?���pC�r+U@˞jás��	�Gs���ࣻ�����v��_��c�AL�X���jEԙn@<��W%�y^.N#��:J\��&����-�G.W�g���&k��+s��ۈW�s(s���jPMm�3�{ ��P�|Z9尷�����M��܊�j����}�;�g�v��sb���V�Y >�*��{��@�3�'O���iU�W�WO��K���b����3����e�cm�}�x(��&Y�Vk][�Z��#��-���[E�.��@/���ڠ�s1~�w�9�t\�aNhc�㙦l�29� �����Ę�X$L��y���yK�ԛ��9Nx��V��#I���(����n�ڠ뵻Ze'm�D�sC%,0k�Ds@5P��d�8%��O�.��@�4�K6�
az��}�\�ā0�������C�܄Y#冁A<>���W�uS�7ۺ�L_���ظZV$I=�#r���6�J�WS=m��ʦ��p�"�������L�Ҏä�8��2�L�ԥ��}�_Kl����(.S�0,�o��'�0y*k�i�g^�� &v���eHK�Ic�K�53��xB<��kck����+��\�|�y�1�#�nG�n���8���hBz�q?�]�=+ �A�
�"3�K���WEIpCt�e�l�7��MG0��DU��0D���s������S�7���"\��{�V!:�b�'>�soLZ5���(���^����){G���)�'K��sӤ��v�&��4U�wҷ����8��y�Q������'����I��g�a���'d@]ߛ��v� �Lú]���"mz2;�a�ed�ER���m>㉻���J����a���&���Jo�:��Z�6�N{t$��E��5��#}_ؐ�gz���'�=>�E�t�!L0"�D$�aV��c>l������<����]�<�I����ξ�Կ���~�Y�nw}J�b6�8ʒ�F3��"���l!1D���+:k��c�0�>,\ �*��gl7 Νs`�N-��P�Z?�q��f���`�sϮ!M�̂�I�/��m�e��s��F��Íh��/w�yf|Z\���i0Z��b�T�o"����V(���_&��w9�n��AS
������9�eEi�;Y8΄"�4��Y�@NbJ{2��kV����;&���̢�� 5�OQ��v�uH�{�"5��?��޾��aߖ˙�ث�wb�R�-ĕ�A�2��n�\���o�	6���Ȟ�-�ө堬E!�;��2�����A��D��k�W����-/5�S~�h��L�}m�����2V�@�R
!۲pX��k��5���.��E�9c��Y�Ac$���&�����5b$J�@l�8��^�-k��ސ��th?0��ȗd�r	�=��Z�M������/�D~d����16��rq*� )a�w���$5��6�Մ�+�<yi��8J8m�$4�w6E��k�M���_�c� �4$�N@݇x�#}����XUsS�F~Xz�?����Q�
\���\n����c~��C��Q�k*ƛy�o��bp��O��7���Dx#�
=�վdߪǃL��3���!���շ��ŏ��t4ڤ�� Do��Cf ���@M�S��jV8|klBB�F(���nΖ��&	����''�c�,C<�~���H���W:80�=�/��f��������"�\��p���M�ϐk���B�^N.�ע4�W�5W�?�N7
)VzF[d�Y�P���R^�UE����$F�������*�����#-���1��+�:�'�I�y�h>11g��.�'~�՟�g�O3������4���v�-S�άC�9%�O��V���8ѕ��w��j��U-g��f;c��
P�KTâ��n>�r-6mW���
��R���ҋ"���D�K���2M�-b�����߶���qi@�]V8��/%$H�)o�ۣDI#���4��Gk������_�q�ZSE	57]�(���]U����d��qٶ�7�֐�[���)q�ԴDĮ��4���S5jSδG\H�UFt�J|I'	R�J˽	R��5����Q����9%�ˎ�w��Ǡ�t��LV�Dʖ�MpmM���M%(��m�-��b�М�S�#X���
���CK�ɥ�� ݕy�.� ���zGT�d�V�l�:ɂP�g�G/ue"F�S#@`��3�Bo�Ȇ�T�M22�YW�UZ�΂;`�Sl�"�N�f ��$��}Ղ-�"��M����YW��II��;�E�&ռ!�KW�i��.�"�׮�J����[��M&���Z�($Su��ķ�܉a���6JϹ*ND�P��I�%Z��u�3߄�Pdϖu��C�F$T2J�@8��2~�eF���zo	��X����,�9yR�4Z�:���� 
F �}����]º@�� ���v�nmUd�U��cU�q�na��#Izb�hdZ���L�S��[��hY/oHG8������釿�&�.�_��eg#�G�x�p��+�Z1�{T-+�e$�x__���`(� �2ӗˬ	e�?�s���������0���CZ�(������-��a���p��@l�S�MٓT���ǜ/�j,���]--U�s?s��6 �Se�3u�{�2R�$à7&�Yb><�Wk�
�{���\Խvt�@F]���+E�B �$��jm/6���h�č���F m��틕���G ճA��dHn����mqY�,�S��~�שzd�j��^���L�,�x'F���8������j��L�S��\]r��HV��LAP()��O?T��������<�*��/\�vL��m����s���I)Lj�����غT��?/J�d8�N�ȴ�B�~�S1�~�_a�8�1÷�E[�s�sSMG��X��[W����!�5iz�P��~��svm�A�%F�H��� �P�xB^Ff�k.�3�E.���wؒ�EL��
c�p��X������f��a|�t�g�z6Vx4S$�����v4�`��w����_G_J�Q`��vd�V+t��Q3�	�nK�M�p��_��S��t`?����@�k.�ZulxU﹟zj*��"1���BLa�ktdp,U<]��d��W��hB1�p��=^��� W��F�tA�38]��CH�b��0T�0"�����1|G���J�h�zPt@e9>�L������gU��1��V�� ,�I�F��U�7ߦd3L�}(.0}�{ޢY{��5 >xagps+��=��SD��K�q���>W�7h�ƞ�7f&J�O7�i&�����GSx�^[�0.��/5O�99�����g2��_��%������jR»	[֯ ��Iw���!Z�"�?��) �$�(Rp��o;e�H[>y_Kd�/qU12��OHl�L$A���T ��?hÎu�|=ѮU�9[�e8�ٜ�Wp�
���\���igt,&�6*��i�5�v[���@R�ٍ��lP�q�\���$c���������8�o�3�g�������� ��l��i#ビ�8VH;S�sƎ�u6cծ����u���9�	�]󯅀��Ը4@���G�H��j�k�.�F�!r)�E`A�oz��1��ћ�a�U9W���$ ��t7��S��-���J�Z�V`KD����=hT�z�+��t�3@���g?��y89���Gk�w�2��ȥH�����.��$DY�$� �Q�R�/����q� ��I��
6���k*��8�����l�N�������+���G@�f}l��K^X8�O�o�C#��Z1�Z����D��S���u�qg����RQ�8�Y?�����X^�q܎��ƫ���N���6�e���7�2��A��EsT��T&����_ƷIH���e�yG3��R�B��gyt�g��ϋ��{��&��2	>���bX��q��A� � Q:��0�O�]��I�GC#���Z#Z��ZU��{�ny/=V�y�LbL�$A���I,����+���%���&����OX�,n��%8f����#(��ٔA�;�9�hd�~~�R?��zġ��L�1��@h��3�.�b-�Ge�nX��f�{p�F{Y6滨p_;
�^���Uhc�L>����������q�Vi9�c95�6���6������>�Ƈ�+���+�ѹU�!���*!u�-�B|d`��on�N�C�3p���&�	w�YqѶ�Ȯ��&)N���ueK�G��|�^��DX����譶�g~o��O�ViJD�#���3�����'uun֔����Rb=�w��!z�.���Z$���&��/�_�WKԨ9;_v}���!�Bg�3c��r(���Z��8�X�)�H|�5Bs��&A� �5rm��߄���\��qV� \_3�C�Σ@{` �=v���Լ���d�����GmU��LD�p����l�	d��Zǟ�lzd���S#3�M�4^�{䠜��
�������
e<��=xC㌣�U%ח ~��A.�"ˆ��-�0��c���_�Bp�/��_,���t9<��Ox�,J��d�*�o��R-
����d`|�,86���o�t�u���þ��J{"���PAX |���t�[R��*�!h!���bb��B��ݜ&8���_C�9Ɖ<#��mC^�<	 ��c3�8�%}�/ƶ3��';w?5��0rងTՈ���7�ȈdZ�*7�H�g}�n�,�ϩQ\����W2�ip~lCY�Y`�A�x�[����M�\/��HO��W�b�?�A�w�"(��V���Rmf�u:a˼��4ȓ��܉����G������c��ʄ��M�b��8��N��')��Zqe�s%�x�?�qѕ�yl�IרGqlւ:�.N�ȗ%5��3[��P����~�����ͅ<*K�b����in��ѝ.��JU�ק`t|sF<]7Â��4-��獾�����=�3's)���C�%I9b���}������#����B����H��t������qЩ�2/����H v*���&�01���y�}N�v�ql�)�ڌ��6�
�^�ګ��Of-�̷���+)���u�gXS��>5�T����\�8�]���=�>���zG��T�C�Z����	?�q�|Ց8zݕ8��!��]ǰ��8u����m����'�{��h�{���>��ï"��/ctA����1�\ޭ]���U��K�r�@��	����>t#�E�A�y�D&��w�v3���o3̾��=�զ�?!�%������坊A҃�*?6�9c11��p��*��P���O&<�-��oe�Ꮳ�Z�-�[~d�s��
�^V���������ܛ�h�;U��4:{.�ͱ2�����|�-�����P�AHY�9Q��[��o5�.t�H<�ņcۦ�2y@CD�����@��jvQCW=-�P���7b*�[J�k�?���+hCͫ�pR���򸋍��	�=�Hn����h�(}?gE�MZn%�&,�8CIL�[VR��1�CBs9�G"��3�&:gal�Y-qP ��j���|��P��?ۿ
��Kt;h���A)Aבc����
�FxB�@=�4S�� �ot-Ґ�7h�bY�F�K��a�)��H��U,%ed�㜩���-N39�?"A�d3�-���(��Œ'z⍚p�l�Z��H�|�vFy`���o��hU<�U���L�F�n���,M2ΊM\���=>�.���3++BI3� ��O_���03�����s����0cϝ��=	����Qt���UO֧q	穱��$ht�oqh�9d��z߭�"c �|P��M����N��Kr���!���ʝ�~��:�ƘP��]���ؾ�K��P^�i����W�JIF���X�l�FNC�^
���W� /_��T��ߖ�I��1���(���!�$��-�e�e4}���\��")�|�u�7�p��	q�2%�P�&,T��C�#�G/c3��OtD�[�_V�El�M��4�:��{^��ܑ.�Q�k�E�Ŧct��(��Ѣ��ԛ'�����n�ee :���PQ�+%`;ݨ�߯];�&䫺�y?T�'O�k�iCk���!뾏���b�unJ)x��y�+ss�;��p�(<��X/�(M�_�t��{�/�#E'$7�("C8��+�l��ͥ6 �b�1[����� 	lnf��.�����ܠ�s�
I5��)���=;�(��L�{��nLn)�)!n�	��C�;�TM�v{%:�nl�X�56�%N��uYh�	ĸ�U�Pt�)4kQ+���ei���s�7qL���K�lS����+6Eʂ�(,4����"8�C�N��}B��R���0�A%8B�8N���K�eM>��{�#����"~@*���dMc�͗�%�0fb)F!]8�,�����?��$i2�5�����u6C�Hg�R��oE� r�����S����ٝy5�c����_
���q���֡YO��ɵQCuK�M6�VK�_�ev�� -l�ҩ���c�=\��U�v�ǠuOUy�R�!K��8vmB�@��e*�������k���Оk�fYN�{^yҘ �6[4	��&
|�U�qm�j�h,'�k��5p�`���sd�!�{�qř�]�|ؼ�=�Ƈ�1�D>d���M�P����s�$�J�W;]��Z��"�!%���Z*{k���ss����6'�|�a���1�Oq!��q)�r)�.�i�xPK�����z@kV���=l+Cش���>��X�~Λ�� ��c���ɛ���QR���_�R��d�I��:�K%�D��jxc����M����³�]��H}z)d�ͳ���>�g��<v��T%����Hፎã��'���Y��u�qF�0��w�ۺC |"�U�~��膳��j
�h'�5&yPe��c �O��F����v����B����hX"�y�[9���Q4�n��J��e0��6���W8 N�/�y��L�¦��c� ���y��
 �~��H����_TEp�������m.+8O�-��0Kj]����8���O'i�x���˭�?���F$�.¥�W+,����
묅 ?BˎDq@6T�����d��a��z�/F��ӦE��˨e�ޥ&���f�ʀ}~� �Ƙ립v"��"s�����SA�+��1�S^�w����q@8W�!z��T�;�pW}�n_�/L�Œ^�Q^�})�7!�O�r3˃��FA�j\&�&�$�N��c�� ����_�4:i�y��	���,1<:l����]bܱ��A�@�3��A2	�����!uI���e��bB��ky�m����}Z��#�oE��)!�eI�p�����jf�jO�ީ�=��F>y�l`D6��Q�N�;����N�H\�"z������Y����g�ݏ�� �OWÀ)K���<�v��?��F��v:F_���:�j�,\é�XD����_��*w����u�5
B^���Hα����)�i��	=�n/��%��[�i[��3z�1�T߅�f-�c����;�*��Q�,(����Ty���2�|J~X��E��JاE1��Q����̓B�V�Bs�\�7�sQ�y��1�����=K��CB�=]��_����=��[�Kl�ޣA�gMݢL��J��.�t1�]���	�Z;�!+:��}��&��I��<)�2s��#�-�G^߼b7NZ�z��5=׋q}�Wc;����F?�i�-��"%�H$yg���l�z�#��38-Z^[�G��� s��Z�]Ps�����Ǵ1B�HI�����.��i����P�c�Q9�BX3}�?7�ȵ��h���w�F��/=]��PHV&H-��C��a���ֆ���{��^�<��5���x�򟆖+U䗟�*�ۉ<<�A����7�����cs�m�T�Y�R���Є��0A+*ط���m��3�`��'�-�#��6-W /�6˗��ֶԱӖ"�ݑ�e�RP��G��[�������^����*�Y��5���N,���P�h�S'�d��
H�wA�+�/� �}M��Z@{��N��OS���u�;�0�+����sY��&��_8'*g'��N�.�
�:2�#2AQ$��퐳�<�h|�������7��[��O� �E��cT��+�����D�?$�����PG]��p�r������X0#;��㯹��@���$������*`��uPI~�99jm��T=�o.�5b�u��m�օ�5`_�b�x['���JFI��ty��o�	��tl��F=A6Q��F��`F�����D��-[��ha꺕3��W7��િAeݣ�V���&k�!�����]3�Ot8�a���.��2qۖ��` �pe�хC+}����9����s�V�)��g�ly�)��,v���{aN��I�ܶ�Vά��R�nx��.����{�l+�#����1qQ�R��&���N�8r�X��,T�siMཆ�0�<�'��R1�-��yA�I	�#�Z���ٹFA�Y���lo#2�X�0�F�}V��
h4=u�
���5��P���ly���m�d59k;�p�6��ʫC�/�n%��Z0e�b��w�Vu��3L����Z��7P.���7�4�EJa�+B���9�5�_�3N�9�>�~��dVZ��d�������)���V�)�Q�Gu���R����Rz�:���su���6�tG^Yͮ�n�"�qU��Ǻ1hv�Q�d܉6��Sj=B�BZ�v�W�� �S"����}�Sڀ�v��M}�B�$�eth]ޖ�̖�"�Z��A�w���l���%�"�%�\�缰�������no�Xh���Qo����}8��i;R?~i|��) ���� �����_���t���JL]I	{�������%vB�=ÄƉ4��zF���.Z���L���ڒ�/����[ۖi;��@*q;v�ʀD��Ju���a�Dp� U�Fg���[���u���Ř=*�@�l97X_�Q��Ô�Xˮ��:�⒳���_R�Wף��Xn1���M>8�K��q��z��fk��T4r)D�֦�P�T\�y�_X\�xV�������(��ں�Ҥ�K�x���9;��:�����?.Ǯ�!�w Vd,$�q��/{���i�ګ�Y�Nֽ�̷^b�<�kܨ�؛P{�K1�Ƥ��o^��]��:{dO���G�W��/�䛐v�!��_��yz���z��&ȼFx��d��'��F`�id��5����wy�������a���B��Q%%�I �Xb�"J��QX�E�%W�n�v��@rz/o�0����8���Ѩ��HJ:���~Q��c+]���j�z^��ݨ�vb��E���gZ���o��L����'!�cU�i>a���B	�Қ����E?.^��i����VD?8Ӧl&'w���|�#��]����%��ec�$(� �CG��|���F�9�`��.NeeHym�7"���v���ݟ����W�A��D�*���[о��oy�ܼ��nwc�,��J8<�S��@�f�U���<�>Z��swf���l���T.�H/N�d �I�.p���{I��ʃm^œ�ִz�Z�s�Q@�~� �@�@�E罥92ժ���>�P8M8_�������=.��JH���>&󳈃Ckqb��#�&��WѹXJ����!�q>}*�NFN/�ԣ�dI-(Pn�:U�8L�Z�߮��g�h���=@@���Q#&�T+%�s�9fͨ�/�?C��h�4/(a3F��A?􁏭���I*�jXӫ�e�w�`+G΀��O�c|��*in���� ��Ԅ���(`*=��(��R}58)V��X��ǐ���ɽ�H�o<�.�8��<��p�(*���-����M�K
-Yp��|q�"��g��!��У|����H��v�DDq)�!��_`2�9A���D��C�+�+*��w�/ߞZ�Ĳ�������8i�rm�s}ո3�l��m���z{���i�(q�|"�N����$�F�Z_�� �*�����t����JtL�$���l乜?�q,�w;�v�Ǔoa���b�2�0pno	���2�g����^��S(0%�.ǐ	�%}y����)b"я�,:a�vΘ�s� �a�β<��0Ւ���7��ù8I�-<�b����d"��hh�;���Q�H!FnTp����*�׉"�9U-�*9����}�+�5kд	�q�}��\��[L��z��9i*۶�93-��;"��]�����t��"���V�tQx�I��:>l6�M��IӾ��&l|��i��J��jilD���qZKmw����8���r׳iJ�M�ioh:� �ƭ�m�eI伋���E��惎�N�P�[hoT̶0��e�g{�V ���=D˚���
f6��
eY:�CT6�]b�K�AY?��|2bd�A6&.������d�E�Ğ�3�J��-���b �`�4Pe?6_5���2Ӆ@���d�EQQ|s	{��J�Oy��*D'�ԟE� �P�T�-�F��W�m��E�XjHH"3�c� M� 4ݦ���ĺ�_���Ɏ�02 ����S1�(���
� 7��I���\�8���ڇ�T�A��ݽ�I��K�MN~N`�s黪����*�F�\`�t�H�����"��`X@Ѣ�y)Mc�h�6Qh�(��Fbc��޲�c����I�(�8�U�Ч�k�GW�t��8&d�Y���LO��-(���pR�+:���kq�Ω��a�����gg���&5,��
�1�8���5���E��[p���@���G~�A�^�\t�!k�2!-�|��U�kiUoc�,�yma��g������,�"��=T�զ͍0�/I��n{"�NO
-��c�c.��t�晤e��j�u>F��R��'#kֶ�����+Ѹ�γ��YȜs�.����5딿x\����h[�}9�b��S*�@2��1���0�w��9e%9ݵ~�t���|���l�f�j=H�f{"��m��ȇ�H�J?��z��#��sc#��Dj�3�Q+�s�|O��} VȮ����˼�|����BP��_ڸ>5ϩ��e׃⣳�^G=4�!����Lt�v҅�8+ꭑ�a���J��E����������(�\:<C�R�T[xh���u�E��w&e�������v�BW��8.�M5o:��kf�(4�<��/�C���[1��yR&jDB���)Z[�e���<���!�7D��8DC��ǒ��=bS�nZo#�ۗ�f`��A�Uډ�5�B� l[)~��Af��)�p����}��5�&�.�M��o��m�J��bI�Z:��O�b����z�I:B�5>� {B�K�$�% �Ψ��� :��Š��K�:�}(��ݩ�%��f�)��>d�(�_Ԓ"lXc�A~H���u2���l$?ȓ3���Տx���X�ǎI������Y]����� ���!��v�U�5��xn�o3����k�{Z���}�$p��S#�!�]�rM��L����������4r����B��Be���G|��ZDx��+��TƢn����I6+{��G7�<d��ax�|~�Ӯt�.��C=�"�H:R�y��
'��ym�0���T�*�\�ozy�w�ѱ��Y�#��>�Lٶy���/+��w���Iȡ5z!�w���1�mZs:������=J�"���oI�b��j��/��.�m�'��6~����41^j\��H��I��t�EM<�F��KnQ3�Q�[�l��|hK���|�E���n��������JR`v0V	�2 ��y��r�)�xBFu�&���GP��߃W@*Zj�Im<nޠz�D���<vJ��I�f5�|�μ��?��SW��`I�;�Z�[��Sc �/q��ߣ<�<4�ʳ�K��ۮW�f�⅐RA�Ԉ�p�sm�X$RΗl;��z�A�w�ϩ���M0�<P���'g�<����Ta��g�W�@�!�$��$��I>�O3X�Lr�{�&#����%X�:W�`ӛ��j��Xs��p�������<r>`D�+<�$��-0\��~���n��4��7��Kץm�~��.��hp�'�%�7�F���ꛏ��Ċ %���|�����Q�b�7~[�Y����L���t�r#��Џ���,�섺X��8P,�5�x��X�Q�a9"���ȗ�xHM1�뾡��$����%�7���l�>qrjO8`�i�~Rw��2�簦�����[h�e��M������c�$�D0l�`bMF��iiE$��4���d���������%����q��X2𺼯�=����6�$;s��C���������8B+v��6�{,�rn.���C
<�2�Ϻ�����6��1�)|]ӻ*,G1����?��d����*Y`%=�$�ۖ�"l6-�"���?R��>�U�X:��xRN�$׼��>=E���)��r�i��_ ��|1;F������r���͓^���5��q�k�X���}9E����|�p�x�@�+_y�jt��ba����$Yz�VCy$$޸u2�Yl�
���d6�ƢFV\	��«ǧu��o��K�c��:�Z7YA���Gr�[+�}�/')�/~u|�\�ict��d�i����bh��h�Z05�O�ѡ�Iz-�M&H$v���G�8�׳�I�N�=�aۦ� ��<�Oa]0���ٹA�]�⓪���a��1	�?xd�w������Y���G��XKu������)���4�Ϥ5[Ã��$�j� .S���9�I �T�)� �PH�J�WZ��iL��� �(�q҂"�*�d�H1��A��ܨ���K���Cߜ	�Y84� ����ܨ}��H0�0�z�k�~���H��ѼS}5�q},���U���|�����@<�g���F���?	�/�\�K�:�����@��չґ̇3�G󧰚E���bE�@�9@�dl\Z�'��5ıG��"0��3T���X�����T#��fވ�X�N��?�Y��xQ:�;��H]�}\�-J����J��ddm�O^3�'	)�-81�ƎS���<8'�`��=��E���9�����ͬ�q���!yX}̆�1���U���\$����P��x��qi�o���:�4Y(�v����?� ��c	g`}|1O�{ΘmU���̢J����w�@/)W�s9��mȑg��t��鶗3�B��w�xsTc����і��D=�\y�Iv}ƴ}�CAkB�Ӽ�aٰ�#!F�l?�r��z�N���_0��T��^�-<�|�~u{ֹ/"!��=˨�)��s�e����lr��db��[���iI䎈�[�F�^�)3�`� ��b?�Jh�$鄅lK��%�����#��y��.���U_:����Z~��ԙ�>�$�/�Q{|�K6�o|�x��E���
��]�Ǡ�iY�^Aa���ᣧ:v3NG�P��~��O)�&W����g�U~��;J����3O��A��-Uً�J�\TKF���3��ߤ�D���"�0Ħ�;�1��J";~p{����xs���RZ�`P.�Y:���EkI�<��a=�C�;�_�eʹo��Yg�!6l��j	u�a�n��j3Og�[���p5�31X}5�ٛ'.̞2&O�(>Ήǘ˚��OG�ǌ�u� �I&z9-!���Cj2��:Y�N}>�vr �ta���3�n1x�b�9�|���:��`���»���=�Q&N���Y=i�6Pۚ��?B���|��0QKd����"n�4ofő�yû��?L�O��7&�Z�B�?��b�H���[��%Zn�}�/]�/-��2I���y@o�[k�j�慨��4߬Ƿi	C�o��ىU�[��n}���qȷFa��˨�8`��_#�ҹF�D  !�x��:a�^	���QE��� A:J@��m�%wb-��նЩ���K-UL�6�j�E�����yM�ܥlPv��&Aq�z���k�52i�)���
�GQ�0�o��+N?8���3��@=�3�mk'�i��7���g��]���eE=٧��w�>�:���b�R���9�	+�Φ���!�NK�%��P��� ����w��1ڹo�b4F�X�w�V��_F��s)�~7SR��@V���D���De�S���{���GJ�@6Lr�JM�%�x��p7����t3�n�_Ռ�j&)��[�y����鳘�p�Z58y�/�� 0	�i{չ-�ɛ��	{�k$r�m���N��v�$CȌ�.�g=�>H�8��Q�0	��M��Я��w"z�Mq��.�]�u���R��G.�i�ϼ�F�b�4����~C~K���� �[Q�Y��VZj@\�7<'$�_'�/����F������S���݂�?l�>:S/���/aR?U�N^���O*/�uL�+�8M)���}!a��eT�.�Q�P�uL=��ŋ�_h��l�"P34��ç܄��8&�_��4r�<q5�xP'q���Ð���}����L��u��K���<���@��4�D �HoJ|1�a��6Ǿ��S^���Y �Eƿ�z �U��f9���|M�N��w����l`�:yF�`*j Vgo��耑z��0����	��H�os��ڤz��R�xĈ�iƏ��"̵;P�p��h*N]8�w�=*�(I�O{f����{�E�CN��~r��|�������^����X����U����d��=��*S��M���e�@BB�����rS4�Q��˧%.�X��X�1rE^؏�����jԊ�p��ӫ�
�8�T�UZp$n)0�F.�H}�WI���՞|�ս�N#����"���խ(���%N�3{����$�n��u	��O"J؇tG ���O�f��ˉ�CX�徼�Q�:�t��WJ��{C�;f1<��۪��u���*a���/�蹜!F���$Ȑ�@��L��t�7���I,�At
���eE�I6ͧ= ��_��+�Z[��G��B����{ �Y�*J�m����@:�Z 5�Ө�\.�W���>�I��݉�5��4¸�6Xۍ4�g�����}���:���9�!��pWq�׻����:bhjaұ�>CJ~�����M��l��/��y���.�"��3�B�;���������_5�b�#J$�$,��Ym�W�Ob���lQ���X�=�{�̖�`�ڜA�Sy����#%Q �J�6��#/�Xr��k��R[�Β��r��+��.r�"s��`�֜�l40��e'I��i�Cjʺ�u�HDjm��4�q����D�3_�AD�v{H�ZG6��G�rc@-����.Nn\*�e�&̞�T �W�r�f�@���qc獔�ǯz{��D��6�,*���"���!'_!����MɎ�R��vbT|�Diu��V��髎СުN%���Uͪ�}ROS��L�q�d��55ػ�J��o���A
E��w%�3'=[h��q�VwB�{E�mà�	e^Y6tw�411��6]�V��r�6�L���LT�w	u���<M0%��:�e|ny!d��.�V٩��]��?? �����ݾٳA�w�Lw滐�h$zHX�i�L�餽<Ss��,"�sz�B�L8@���T!�;�D���*B}�'��J�Y�Z��EҢ��O~�[;���`��T���aԬ�L��&<FR�$A�)��  y�����"�i������R1E�Rү���$��Y�#}�b%A�5���y�CC&nl�k�/��� +Y���E����o�g����d�_nq=�S�������@�"	�i����G�:l�V��k�uu?����i��o �EP�+B�t�?�Y��g6�@�<���� sF�ַi�=���1�M���ݝ ��U����cF(����B&��w��`	uk�8v�k,�wlxB�RzSf��	x��Hk|����q#�����*�Q �"K��b*��e�T%6��.���oڼS��K?���
Μl �����H���^�Ć@��uv����>d��@(�\�bM�F�'&��e�_:{�QH�h��<��iZ>i-ix�a�-
>�T�/b���LE�y��G����1%��̟�Ul�5��>��l�ڷ�j�`f�`Xn|Hv՜�	1�m���%� �����TCx}w^P?v�gxm����bhb�#��TE�v�1bQG՗�{]ӈ��2-&�����a��>Մ�q���1Q��j�N����joh��_s�w�
O�wQ���,h\a]�*�"�����mٜ�%@��ڎ�ߑ�d�_)�{6�R��p�"�v��*xYiA~@l�Z�~�?T�=�B��[!G8�H�_'n��>�B0}t��>��+�!r.*��in�d���u�+��k�����@���� =���a�Oia<l@�t-iKmQ�&���0��ͷzKkQU1?�쑉� �4u� �/H+7�D�h�̓�ͅ��s)��bJ��9�3�I��Y�''Ĥ�zRc����[�K1����on����;xi�b�҇lf<X�y#d��y
K���=Qz}_16��ΥU>����.���`��P$�Z���c���i"�Zd,�M��|dH�ޮV��a��e$�k@�5�sd`VG�������3�:�M=�u�VO�a� 3�g>.��ಞb�{��2�dM>��n��(�Srh��b���řA4b� ���j���ř"��4�����ͅ���jH�	�����קΕ p�+��D��'1����`cgk�����1�J�r�Y:�n���g��»*�R(6�J�C����?��]GO�/��g�Aȟ���k:�v��	Tz�kh��A�O�� I�X<J,oOE$�0�C������U_�?����4`����'2q�Z���h�V��:dt��5N��Q��sTx��e�Jj|�Ê����1%�����v��X&���Qճ
��4KL4 }ht\%�ȆT�����Tݱ��[`�s7C]�^E9���L���M>>�6�P�#�b2+Ԡ?�"a
�F���l��%�"��ou8����#��\�ڑo�:n<�' ��<S������� r�{x ��<cb���U����F.��HX#E������G֛ly6(Kq�J�^ɷ�Q%� �y��e�KJtXrݎ�X���T3���/�7�c��zf:�����z��,F}�����K�~B�c�F���OW�)�O��ѽW�eY��GA#O`���2;� ��&W���ynkށ��,7u����^�^3��r���(�����c���G�Ao�8�nhf�ѤXO�'�7S��-�"��|�a�v~!�t�,s��
%mX��.��"�� �lg���t����<�FIB
�'^���T���9��|:��-�f��N'4:�U&2��2T0��PX<��4v<E��d�4��j �]������Nb��Z������
Œ��{z��K�A�d���5���>��G�j�����ܕm}m���9�p��Ҽ+��/$ݪ����è�QQ�Z�,�~��U��/|'���Om��3,F�^�z��ˎ5t���{pt�hc�B��#�s?/�U�Ȏ��;�(�?$��+��8,H$�t��5���E�}�	��
��0R�Jm��-к�`:�;�3MN:"�Mr���jE�YV�j��x�����G4{�xt���L�5De�H��ڞ�Q��x&��!uA�4�N�ou���0Y�D��G�q���[���B�2��"9�Z�h;!q��#�&��[�bs��px��WĮz�;q�mv�h;+�2ıT������݆�QăH����H4jS���T��Lb���~�U[�&@}뗧9,�9��[A76��7/5�iȐɗ'k}z]Ǜ��q��{,K�u}�|CK!oB��n6D?������kwJ2�é����.�J�S���������Ozd"l__�����X'�ߊ9z��u@ڂG3okb���r���=��ݛڀ�#j`w���j�)�|nw�:�V���ƣ��Z��� �V!yƄ�ٲ�F9���&m�~`v}`&
���ɂ��qT��t8E)
��i䧋7$xC �%��t�Z_�VQ�ЬW��im�aEc�N��/y(��n%�5e�cP �1��o�bq`��1x�dP�u2'�[B��`�Qq@�i� fyL�v�[7��"�dw��XB},�b[,���Z"j��C�����f��>���1���/��bR�L� 5��5��5$ihn{�T�	v",h=������Zߗ<�@(�Ԇ��/�N>aa�� �!��Y���ɦ�Q̱�/�3�@X����l�l<�,;S��R��+�v��v��O7�;��3��t�6-�d��b���8-��L<�pM���Ǌ���4|��j�ͭ�������C�kM��n�c��j�?���6�~��Pb�3������R.X�r.���&�����AA�d��9�e�&����Ɉ*}?w���wB`�7�]���I?��N���>�W��1쪗s�n�AV 3�=�\[�獧�&�ss��5��M_lͽ)&��$4�����=�wr�:x��e�����DB\��t���E���_���@�E&��9��}z�N�p��bĺ���k��;�q_:�y�yg�J�u�������Լ��箇�G�j;��L�I&
X�3�"t򦅹�-��Th�5��*�pC��x�D��fz.�w�P��A��e�6�ܞ��Z���wL���@��!�}�]y.����(D�V���hNA>O(׆;t�&�=v*�j�e�=jx���J� v���R�,O��r���ǽ���3d�0"��C"�N -���405,�7l���I��,�U�uA2��AS.h�W/�JLP
th,���Č_n�r���m���,�b�g;�*\�j�7Df�3��V4M=�N��)���һ�<�k'zć(�R��ўP���e>����{*q^G�˳b5��M�0��	ұ���yҤb���~e�f?<گ����J�<�cm5Ɛ���=�_��0�a�$��Q�4B�	�����X}�R�;�W�����M��|+�� ��4a�/���W:og��s��<n;bL�C
��`��v3�޲|Rv!Ճ�3Ͽd�0��JЍȏ͓*%���rؕ8j$�[�X��l� L1Ϙ	�Xͬ�ټ~��s��h\Z9Y7|;��D�u3����������@����/��9�q|Q!ڭ��Ԙ�F�ߖ���3z�^��bh+�sz�v�p?Ww�z�;��6 �2y��V�?�7w���Iͫ�kNs!�缈X8r}n�˗�q�B���f[��C���BOHg���S��)����|����v�YGL+c|8�i@�=�S��]�3np��춸�͓&E���@�7׿ǑVHL���7W�ϻ��I�r�fj��=F킻�Q#�U�8>�:?��Ny��� �c�|��'ɾ$�^Cz�R���c�~�{����D�V�p�y����Ŷ9��h�ʐ�J��|g���T�S+���(��-
@p[#��ʹnt3���G�66l08��o��*�T��R^��g�'��d/�ݍ[�z��n7i�|�M�S����ȚZ_�E��Lp%�����C����#�Y� 5�fV��t�v�IS�R'����LwF��֫X������U�����)c�[�Kz��� ���`~�(�V[�L�rA#`�<~/�}s*�h�(�ǿf�.hc�ɵ�^�b<Ն�Q�ߖ{�V�[4l܉D���-��"��wl��*��vD|׻��dx^%��߅ɺB,u�o�R���H��`��P�~��U��.B�˖�̊Ȃ�{s �f�~ 0#��0�T6�
 i�(]��q��ֻ)�&K�9^����YoJjm�;��wTv�vB��PX���j3�<�8=�l#r.oq�W�M8���P�7bw��������|m��B!h�a��7�U��XFW��<���<׌�M�z�[��]��Rqn�@�y�/����2zv9$K^�gη5X�b% ;v�D������ZY�ɜ�J(E�¢�\��̷�����7�QC�]k�{D��ȕ��$�>W:�5�9dw���n�dޞm��P�2g����/��fF���is'�Is$�-��ذ-���IX�c�����Z{J���8��1� D��\��~ر�Crh�wsػ0w'��;��DZh �Do���C�����T��	`=ea�bڟ�D���E+��j��TKX�Ci���ݘ�7��	����/|����3�q��]�s���7���.�������[`W�)�9��`_8��{w
M�+���HU9_9���8L�{Ί��g��.RݘH�*�������s���~oӺ��dq��q�u����7]3�l����6a;�;#Ϝ\ȁ�^S� ��M;��*3�|$f
�!}���Y�V���*.��(��x�rϙ�EgG{��U�g��u����Amd-A�N��9KƎ1;l�W������e��=�S���wu##0�����%"��o�q{�Um�N>��O(�����0q��$��;���
�<�l�� ]��u���ͺ��2��(�<yHa����\є:��I&������8M˲�����ϡN���"c@��(�.]�?��V&A�����3�Y������y^h�B�
	�c6��ت<'-��b������؇�
�"���rS���i�_gM��z���ԋ(�W$�L�,��&�R~:`Vڀ�m�uQ>��̩���¯��G�u,���P����+N�<p��fK'Fb\�pU �aٝ9���}-�ޑf���J< �[R��'w
���2�[�z�[5�U��tq%���E)*�pz��{H�o���[RL#|�}��ɱ���~��j�{�WRGf{a�^Z'�ob�]��jB��Υ��%=[QF��B��TCK:7��%C��U�7S��A�f�"���:\M/�0�-���l3�*2�f����7`��m,��ޕ��S��X�h����F�&�EN�t�~�g�q6�@.�6r�3��ng���L�;&V?4�[6)�B�l�{lRYB���eW<Pl���}��/qʯ1�� �rmj������dY�η��a }ɻ��w�'��x�}�0F�:$`J���S�D�ZB�.���\{;�)J��Lr����D&�=��q^n�9o�#�t�2ă�<�Mm�9�A�fKY�V�a#Oݦ���ʀ�|�5�|�"�'��J��r��a �LE]b��j<R�n����C[N��JU`���6�=���ύFSOx��`w�i�zu��;QG��#�85(Ĉf$6��ghU��Iq�,�9�h���m&��Hpܳ�Ӱ8���+ZW��c�A�*��3�&����A��H��K:���g�PF�:��j�| �`ښqO�}��1�'zB�W�[�&����.���biU�Wl��Vs��k�橍�����[�������X��J�p7�w�?)��C-⬭��lsp����`��3A¸ک��۳��Qm:�˱v�^�����v�;�	��`;f񯤮�.$k��42]K�f�
r3K���f!����MƐz;k�Dw�Լ�&�G�w	Fp��b�g� m#���i�`{��V��t/��x��D�s����N��H;�G��|��kzu��8/���7�@W�{�+\������6��p�z�7��ٗ6��zA�y	.���=5C�Efn8xU�5)QN����¨;��8����~�֮��f�l�UC3#����
MZa��*�I#�$�JgD�_��	F��<��MW��أ��6�m��6n�3n����vhw�1��m��C��e�˗��Y��Oe���/��Q^�&�-n�T�,��QF���Ǧ7ӷ�mo��m���)H��Ƒn˰'��^�z�c*�De�b ӎ2���	��&Vo�g v^c�v�o_�]�'�����y�i����!�m�ـ�I�NBR]O��w�dF�;1��_J"F,���x2��eU�U��z/�H<jM�L�ېy^R�.�(��緉���� 46�Gޑ!^+��Dc�+�Zr�v��t��Fy����F���抵gPǡrz��4X��Ӣ�bB�z��-%�؅{@���#.J���۩�='��j��gL�0�I�V5(��Ӫ��i��a亞���(��I.��hXc�D6o��3�ИF���5Cj���F�xZ�Y3�͐hpG�����Z��bǹ��_7�z)'ʾ+Щ���Z��d"v��W`@c#��6`��u�//��|j$\�#�~�d������ɧ@
�\C�4���<�|jNa�p��v/9�� 0G(:V�c�.`۰���pT1��q����1f��ί�۬�D�kkP�XD��-���,\�����1��Ađ`3l�Y��o*��X.~���4����a�����˳+�{-�d>ϣ� i�߄(�vZ�9����Oy<w��Q�������xun��_��VQ**� x��pw`Mb"Ud9������]@sƋ���O-��U[t�7@�Zd���i�6LQ��٦79�Ő�a�0�f幧*����*�B�	�k��fF�@��u�S]�E?e|~y8�>lM�(��D}��Ʈx
Vc�௼�:� C�d˫-�pGyߌ  ���]T��7Cl� ڜVn8j�Q2^�.�!"���PaGTs���"Mݴ�_�X%@r����9yHaE��:�Nט��R��,���tY6J#�	���kl����M������X=7���a��L��Ex������"E��[L��(&ԇ�����Co^yߞ�<��{�*�@
���Z{�����Z%X�n_e�)�
�I�?D��}-qb�f�9�6Tv��H�O� ��m{ZZ"��o]����. Nd&fVY�t�"�MQ�;��	s�f��{��1pEz�f�%�c���T�.F���~z����'
���۸�����K����6�3KQ���+��TӲ�0L��X:!z��UC�1X�фU<5�����#������m.�P� �yyT��ڢv�Ecҳ����Մ.|�g�(mD�.�7��`i���)oo#��I����
�8l��b/	xV,~���ܦ;���� �vč ��ܕ�(1��;�NEIi��}+�ƚ��� �g��:��M'����m�l�g)屓⿱����0 �bG�t�B���<a6G��Et�y��f�̂�RҲ�+������
�å�uN�W�e���)���9D�vи,�D*M0#�rU�ْ�B:l.��;��.L���VS��E$�f�/��R�L�sXmH-��,00dm
r"��(��+Z'R?�	�ֲg ^�N�3F,����Bg�vuMQ^����ݧ�.Z �4'#�\ng��˒��^q�ȿ�1ss��x����}m"Ӏ�����gv����_.l���R�Yqz�ў�[�IOWڎig:s��uj�Mm����~e�>Px��^�O�"��0R�<�#�1LlLae��޶;5������wޡ!!)��o�ne����ʺ���?�1Iu2�?#z�����X9���'rh�E�k�r��{�vd�/g1ѶX����,�o�cR�\H kl�cG_+�|��&�:���H�Uγ����S��[#����#�c��YJO�4�EЙ�o��4"4Ȏ�����Co �%��������K��`���nư"o��0�S~�T��-!���,��&�����vw���(�\Ő&fHG���F�j}����M46i�si=jYu��?H��h����6f�����o@��Z ��l�l.����8�T��x�c}&��|��4F2�8݌����L�|��Q���ؽ��(b�>`���(�,��S	8�d=�D/hh��yk�j5p	���"�Z���5��^a���������T�����(8h��d��J���J�|}�U�2��bi������C�4^��T3�,�r�H���Ds��5�5h�g�L1��C�2u�D���е@@`�ɑ��%m_P2���Acp��߁���[&����z霧v���vIb|���y9I��?9���W�{J�I>�c��h6�h�,w���?m�䆚Q��U��G@Y�G�
�X���1'��D=��������^L�Jf��p3H$A�����+����>:�2���r╷^$�R�6�˘�%ȵ��g��Z��z��s��˫w����?�S=�NH�C���	�(�Q�H�����,������o��-ԋpy��_�/�n&$���ZKu�-<�v�2Y�h�#�Q�KUA��q��<,կL0)q���
�ڈKß�w�Y����!���=�{GfR1�TH׊�&��F0��ƾ�2&���#�>5>�W�H�XgN�_��xv�74uL/d���c��<��s�QJ9���P�\�<ϱЄ��r���$��r�=!p'Vr����}J!��c��p����W�C�D�9�Ѝb���(��ݶ��e��M��L6a�*@-0$�B�7�����4)��o,N����)�� ����,��g(yM1�a�4��%&[�uR_�)��[S�]�7Y�g���{ �V(�Xk��}^��͓i7[y�2�;?��ܑ�@C�����{�ѹa�i�
`�3T@A�ߚs3ԓke��:��UA(���]1�]{8� &� -�N�NV�n*�Uk�n�$-g���5W �c��S�)�﹀?Y<�m�c��ƳΞ�E�8���[�.�6
^�L������9��?7䆭5B�7�b�����j�왲Ϳ��s�^(eg|�����Oy�bl�����/�1n�)�}`gW~\��e6L�{�k'�E��h?ԸZ�B�L��B��[�_�w���	˺M>�np�x�*o&���ׄr�(q����6�����Y�G�1���Q�k�;��@���*��)�c2*fKo!�E��m4x��p�߹��]&OD��/�?k;��3�B���b����I)h�y6��X�=�)�]`��**F�KAB׵�����˩|��38!Wa88	�Ǳ�	u��吓����Ile�.u1ؠL����q��.�x���qġ�S!�����v�z�pv�c����Ɠ��P���mb�Y��dq���Y��Md��}ef@�!!�Ⓒ]HdF�l�_!�,�Sw��[Μ�/��]��&�}v�:��~��d]�,�\85�*㧐�9Z�]G?z�����>7S2�WwY���M����*Y�S)�����2�#w�J�2�瓦C9B�Y�4V��"�i�_�]<!�[�(��ΊC�yU?�Ԩ �y��t��M��+�ѤǤ�ڽ���v��c���������i	��B�uE���-^%L��-i�̤m�v�=,˭��/�jS���<�QzMS}o�xE��J7�k��~H|󛺯F��5X��҈�f��S-�q�(G�Ju@n�?[�v�{U>�����J��L���[�MQ(;�{}i��O3�
���1�̻n�N���g���l `�Ʃ�8`�c���4��G]=%�I��>�i��fMn��y��ǉWKĸ`�����J��1o�x��(��d�7���J���WQ2��T�$�;���?�+$t�jj�~���7����4ҷ(i�喁����̖7ԍΜ%��W|u�Q��Y|jgcl�WvM'u���P���������ҋ�/�*:���8�nm(ڮ�g�7[�j��B��2��''��\�s�ԧ+�]��P� 0��A�<9�06hщ�}�Y�v�# Fx\1�@S�����}Q%1��F:���H$i���@�[�$�ſ}��93U�]Ok��ډ@�UN?�l�3����0���-�Ct�u�aط�d��J��Їz�d6%���B�_q�Vrr����}9+�/�4T�|-�F�C�ͽ4[��LF�c|-��z�b�]nu�bۈ�!�\4�/�3�/F�J�5[+濙Z�b��j��7�G�.67m�W��a���堙u�^M^uD؞���BUHL�Z#�
6�v_��I3�[���xb�?5s��ub�k��ݼ�����O�⤆�c�*p����pU��U� �P��6��H�1W]�%�9���zdsX�u�H$��7<87Y���t����������iB�� bv�X�n �՘#"		�߳��C>�����7���fr�4`u�>��̕�3+克$|�*b7?��r����㐿�\�wsws���XX�`663r}南�<e��sA��%j��WI����FlQ�f��n�X��o���3s��e��_��R�Z�]Z9���O���x���������Ma�HE6�<e�ȏ"�o!�A=��X�{'S��-�(�R����<�5Ծ��n:�c�x����r����6NHc�T�7'V���GZ��z�#@�G�z��INw�+{��D>�B������^0�(��>չ�,Mro�/+�s��r�EtRH���E=J���p��H���������hoMo��'l�On[�������ݪ�T��r��Fd��m�ٲ˨������k�Z.�!(f�H:���X �5����m%DP8�9�vSZ?7s��0��h����M�7ҟ�
�~���↑���e1�dL:+)�u���19BӼ�s�Qr<R���%�r��p��P���M*���&дiQfQsm�Qw�$f�ߍ����{����⹰Ôm��^'ԭ���L����Z�O-������ZQS=Ҍˇ*Bھ�Ey��Ul�E�l���D���T߳�֋��*M�H2P�K�}�kq�27x��¦���'`�F�����~[�8Oo1�߮�2��M��~���'��f�.Ӗ���~��k��To�2A���/��G�z�.B�;�(O<�H	��-y�~Q�+�_wߩ�}~�tԈ$	��v�ط��e�~�
��j�����,�	mVXM&JНt~���$�����Zs:�}��wD�q�ƎJe�ҹ"��pH	j�R͜�eg䂶�+$Ʈ��ME���������8��s��ϒ1������&'�,�e,���`�W��Q�\�=��l

���Y���G���>�N��x�`��v�b�2Ds�%uZh����RbPU+��5d�X����BzM�`Gv��w����/I&�C�d��z*�j?[���KVN���Q"0�y�5߫�U���g����(D�DE��ΐ�^��0ݝ��#s��8�������'*]3��I����V\؆�}����!�r��Q�_4�)��yK_=�|�������������=j_��ni瑒c��8�VX)}/�%�ћ�SAp�~,��o�����FљSx�~6Y�����1G�~~=���$��
���8@P� '����}~w�H�Ѱ
�v�Q����V�>v�n3��x=F��GQ������"�!t ڻ��oi����j��2�F��g��@D ���%1�;�̂�����(�F��|��n��5Eu�!$��7A�q���ʄ��N�Z+p����)g��=��A�b�=����rM�Q�2o.]�P/�+GE��=3��!�@6�~8�q0��$�\+�K�tɕ���hg�j
�6��@�c!{���q�v]D�"�� ���g2e捇��O�M��TVVH�ď��^��'�R�'5��pɕ��U��YՂ�
zk���W��y�XR@5l�P�N����~3���Ԑ_�~ �C.w�?u���ч+�K� ���@?�FK��������оEC��J����c^j?��1[��Lc�N��W=ޖ�N�6~b�E&P+�(����v7�J�~�6	���;$��������������+r��R�mV|c��-����z:��7r	XasC�9�o
=�<�u�E{�q��ee#��v�K*���O�F�1�p��׺�6�HvV�yu�G��4�{�]>���D8f���h����1�d!А���P��S�GU~�_GVPP.�
�X{p�sQٝ/��/,�#Q�(6љ��������*-8$٠D��դp�)���Oy"��,Q�d�s�I{�SU�
�W��60��Ro��LS�p�KS#�j��j}.�o`Xf{=n\۩�D$N�߯XT�!ͲRB\�݄�&��,6}F�c�������O�,D�N6O�2�;�r5s�<}�ÒHuN�u�ã�\�֥�S�Q��'��gr��� )���\!ڟ�ţ�q8��]d�/lw61��}_��=n�E_�0�Ÿ��բa�Bpܜo�A���(�sF*V6-P�� K�i@wm2�^�P�m��}��� ��
�^�Y�p��ϰD�X�loGYuZs'Fƚ��P��f�M����ۻ�#s�I�CRk�`DO�r��]��w��L�xA�oOO�&��
u��<��t��
�A	Z}-�}��"?�-E(d@H� ��p㷈���t@��US�&�U���uw���X}�d+�}�m:	\r��<'@�Q#����:߇��W4�)��S��<B����������0
P�}%�.'"ˇ�L9����Q���������Up�6b
��S�Q����x�t��) e�j� mZ�^� ��Y�=}�/���<�,�  ��|�Bočj������G�-��c�Y�e�����Z �2P
��NH�:ovo^�ؖ�2/���4�Y��V��ó-Y��L�}�l������B�`M������F��d^a�{F��n`���F�C�E/���/)�}'7�]�֝6{�}�zh��-�6_�^�Q)��D`��]������l�g�x�D�Ä�����n+�-��%ݴo\�{S]oG.Q`�����s%�~A��k�Q�R=g��t�V��E���G��թ�]�cô#0�<tW��qN�e��K优4��|�n9r�����J}$��M ?�մ t.h�,�<T�*b���e�*�_�gp���?1��@�67~��#��ƺ����T�D��<��o�F/�����φ�`�Y;̫a�c*Q��A�쿿Ӈ9r8*�|6P�Ӏ7+��|@:�	�۬���v����L�1�i�g�^��K_S���AMȿp����?�"�p�f�O^��8��jѹ"&���\T*��6W����w����NA	�>��k�Q~ldJR��q蠚�t.�%ŝ�NgD
���8��%Z٩:1 ʕ��/	����V]�q�0x�h��B�'�̴���f��TdZ<��{ۘT��m�O��B�.P��U�z��X��a��B�e�`nR7D��=sJ��r��=^�Z�:0qO�1��A��O���y�9��,�ە$i���ȼ�\�1X�G��B�zb'�.�Z����<���ao�������q.:#��T��,�4p>�B�]~`�M�M#.����~]��!��W�'�i�3{V�ʢ����41��(���4�*�5�����[�:V;��k��nd�J3/�	E�7�wHƔʌN�/Ze I���E��Qbw�&ݩl�U�A�wy�nI�L+{������F&�ej��z�HNg�}�!���&���"ߒ���Q��V��7�R�� �����G7񁶝"n�)F6��x��c�z�¡�T�^��2l�>�$M0�w'tԽ����Uux�.�o�Q���5�G����-_�`Y{�
5��L��ʂ��gy��.��ď��2���P�,Q�B �d�l���H���X���y����l�������oE��Τ��ㅆp�-v�s�ֺ��[�wP�B��µ�޿4F��fK�e���I�h�Շ�TR���jB-�]�T��?�5X��h_��⁉�%�
ך_apo ���gn�u~7{��?D��+B\�:g�W	7��^BG�~A1y,����h'<P����2��e�`%荼V'Gr�����3��1#&�؍��ب9.����V?��8����=��q��):!\I�'��K����w���ӑ���iZ,h��2���z��p�O��� �3i/� c&1Vt<�Q�J]2�[�,�a�r|Q�\�ܜw��u����EI� ?�
x*�!v�wĄ%��*G��;�-Q��߹�����qr��튃�9�/l�֗�rH,�:���ʅV6�%����İT�����&%�՚�U]�>�ia�3�RM����z̒�sJ�v������!bqt3�tJ�%�2lxV	sS�<�ݿ���3p�=F�^��-�<2��_:��m�����f}f�`֊k�=��D��hE��Tє�)[���3�頃�7
�I��Ï�:�\�M���E�H��7�Flv�M�6�Dx0�M���¾Ph�2wk�x��e�������D��%J���262�*d�������j�RފfXR���+U�*v{+*��Wi��������zԒwjNi�g��n�M\d��>:��n����=��z�=%�>^BLqb�=�"M����,���j�A0�?�oux��uۉ��ۿ��l�g�6��4�v��e���7�wѽ�a�>����r�������K��
�"o��	q�<�_+��ž�5��~ӯN'���ɢ�sg^ڈ���/k�]�^����wÄ�AK���FJ�����>i�N	������܄N�d)�m�.@D�r�<.�Z�s�%�RDX�- c�ܑ�)��.��⋩��_6��xqJX������44���ғ9�7w ��M�Fm�쳙�֊�#&�>�	�q�/�
��{���sBw��\B��Y��<�S�.���1T� ����xO+���������M�鮛��m�^���?��Q9�������%��]���A����լ��n���MP�Y�8)���(<�f��� ��%HYo[_��֙<N^ �%�*b��:������i2�kw6�q��'�|�����`�UZ�O�UC���ͱ_���_�&�gYl�݋�B�a��_Ú�{و�C�:-\�v��򘘚�.O'����O!ͱH@����y�ز�����+��(�ֳĔN�f�0b��)��w {LN�jCʹ����W�6T�Ec}�0�_�/u���恜W�&ĵU�r�2&��M��#���ĵd�Te�`)��"J}����2��2��>�]r�:nt@����`��`����\-7d���#qj-�g��ek4�)�&��0kVk��j-Qv���&�w|�˰��2����F�t�I
��ʡ����I�\�����'�"��� x�2-qVX��A��:�w%��F�$Z#����<�FPH�7@/��'�*lO�n��Y� �/pt:�l��#H	�ɦ�	j�T��2*�����,����ֳT��`��u��/ƤA�����kBI;���]�����(Z߯15=0�ǄJ	����"��]z��<�0�RmWZJ�<<����V߲��_���ù��E�/�ПϿ(L$t}�:O��%C�7L�&<Y�{bX��@��##n��m����t똯q�612��6�Uq�xX�O�[	_נj�-�#�� �"�7X����NP�K!&�������s�|��U~����v�>}f._��+2����{Y�5�`i*�;�/F����ؘoJ��F-^�Ia�G6f���<�>Т���{�L��u9���qW��o�b$��~�Gʀ�Z �� }F�=jf�@�ޅ^�����K���uË~Nm��H��1��.�����)3X�}}i���3��x�O��{D���b�,�&4��N�(���[u���=r���2����ᢶ�ڎ{���q��П���+�D�Ip��ƀ6W�aT��
Pk3t�Eώ�u�h�}Ԇ<B�F�	���M���D`]_��p��Νs��7]��2"H��y��L�z87�Y���PS(��Y�O8H
�x�����'Պ��
r�w��/4���ۇ�ިe���O�>��5�g��\�0�1h(-�ۧ��������I~��b���������E�� `G�\cG�����Ψ�pffCU��~U�3�O�=\�w�����O�$i#}6!T�����xP������ŕ�B��΃��;�J!�L���5��C��cw���;A>lt;�Ո~0x\��A���|=�9�
	��PX��J����)�+�M�f �.�¦��e=
���Ʃ0.�H�L%��J��7���G�ja��,j� {k������z�~FQa�O��LK��%�2�JS�
�	E��dj6e�`l��@���S K{�M�����8/m©yO4�,�e�n����8���4mZ��!v��ml�K]��G
Z9F��#u�����i�.�����yR��*%g�!e��ka��<KX��C�\�W��e�m�=*�N���u�I [�q3�*��U�������O*'�W�ބ�����TN��Iww�w���	������8��\��=k��aG��@Q��5��Ta��4�-p>��AܑPo���f�0��ߌ�D�"���7�~X���qe�s� aGE�t,N��3,�F~D�\�0'�~=�w.y�f �w%M,+y���'���)ZNR�F|t�z߯��.ub�2��iR���Y`��Gdv];U(0���%��6�@����Vϰ���z���HXE���� @��oЭ!�XEH�b����Op9(K�"�mk�^2�}#�t��	�2z�b���B�A��wգ[�o^tSx� �^, ��PC���V�* ����>�%����>@���߰�>��=l}x��S�&n"���p��c��e��n�Ff.pZ8���,Xu}�zK��
K�EH���;�-[���G[G9�07�
 ��+i
���Ȝ���C�6iЅ�
�Q
�#��;���CG*�i�α}��p*���3�1���_��
��hڛC{ Ò�D�Tc�~:����*����}6� " �5e�]
�kn 2�b�3���>K
�&���83����3�նF-'&�p[��T��\d�ș<+8��8b��_xs�֐��a�����L^��`
��,���{�Ʀr|�[�-�F_Ł��fQ��R/��r��f�wo_��G�(�z���d���*]?�Pg1KT�Մ�+��r?��&�-�#}�0I2v��	�b���J��9�p-%&z����Eeu�����/<���k;cW$4A�$j�
`�)�ANN�_F�W�8`��d7�*ゞ�
P���,.8C?/�K3ϜcWd<�$�/�T��٦����3�0�l�f�� K䡷������ٮ����ٺ��S��Tێ�y�9P�*�r@�Ȱ��1&wTw�~	K�CT�z:Fek:{w�s�Lj�ib����m�e�F�L�kWQ�+��î���&�:��=�U-̓��]���#f���ۿ���xrW'x�W�&i�[kB�(Rx-�<�H�� �s�����/�%�ő!���]ckR���؄���M=�;SXD�Y螚WR�<X�q7H����n���6���TX�X\CF�b��/�k�
�7�{��&s��z[ %��4��Z�,�Z�Y�z�ւH��@k{��6q��o�M`�M}�4Va؜OP��.,�}���I<rn�V	����w���2�8*2���9d��ZܸW��.���Q@�Ǜ90sJ����k6���VY��������1����a��FR��k#�غ���G������N
# l���(�*�r�Sv�fǅ�9nkq���]��鯬U�������g� M�&�-(Y�XR%H�En3��:%A7�QRŘEK$D�
��Yq|;1���ԗ.P�;u/����L�M3݋��B�{����*��/+��"�����YR�8ʀ̂���8�u���[<C��k��6%���-2]`��D頮潠GRb� ��y
ư'	cI5�e6��sI+��MRr����|y��7$=��=ha��c'�[ܬ�u�T�-������jd��ӟ�\����A��w��j�<^�>����ck!�R~�Y�7���i�SM����������)�ďZO�~�����%�<�]ᤲ���60#��B4�\4�V%�e�Sc]'�x��̫3��F����� .`B�=��ܾ�OOJ�ŷv,@�\η�J�ӹ+7ל�J�H��D(�38i��i�n95T;�"���$qx��C��c>��.�M��K���;�ŀ�R
�=�9�<7g���rN�U`+���O!nOSH:iv<(@r{g�5��*<u���G��z��V�$^�I���ѱ�f�����j��?A�c�\�<��r��r�J/Á0���ҟ�٨� :�dܰu���Z��8�f���<{Z�ssez������1����Q�d�MO#������*��;x8+�lPq��·t�n�(�GV����k"@�CxbG`�Pt�e�am'��i�ޡh�V^�mF�#��q�7+��q���[]e�l�;7Hb�R�����K*Fۣ�:6*3W�a*2��spJs$�
�L�m)�S�~z�i}�w����F��,S�э��|�d/�TZ]���yt{/
�],�_?Ф��-m��ei�e��%��A�%����b�{|B�uX���l�j`��`�����I���]��_<{
��8���AՂo�/A�pnT�^6������
D�u8�7�)��{:Z�z��y�:;C�;��:��_W��I�/�_Y&tC�Y �4u}���}\���@\w���Ų�_�jX�u��bVg?*t �!G5o��ԫu�2}� �"�~	aW�+�_���j7E��#���PVb&�멩�����/{��OPdᱛ�S��H�VP9ߧ3iK_�9��O[G ����;FB^�ſ��{a��������/��u�	�Qyq��T ��(�ˏ���.%y+�<5�#��!n��ҝ�6�H�R���o��)�7l��g�grԱ@�L���NCԛ����B�&�ʘ!D��f<||��J�q����N��ɕ��&�ϘLHA����-�?Pΐk[]��x 2���d
��[Aˌ����VJo�(v;��p(x��f��ӥ�
;��[�!5��m8���~�d��o�E��/=M��s�^�Á�E"�ZD7n�Jf(4�7�>Έ�ᬽKej|;����~��g>��(�"ZV�h/���I�
&�ɘ>�ڷ�Lz���s��/9ZWlZ��C���]Ӏ��Tj�����;�,C8Edt#G�,m� �d�h5��W}.裤��ĵ�t���tۓyȦ����
� ��ܛ�+k�;E�ƫ_g�b|^m�����NjX{��a�s3N�Wt��(4S�o[1��<��������Z��,�O�������S�� ��C�Ps�4�����ˆ�?��W�؜��wi�ܞn�.�+NEV�_m�W���`k%���������l�i�G�v��ڒ���S�o���Jn�Bp^��nYpS0�8�;�=o�c�^L���U�آ�e�ͼ;s�q�gW ��Q�$9X/�*]��}�uw絎���%\i�c��F�/�ё5=ކ��Tǧ��BVG5�(&u ��K���>� ���꜑���%�,�8�[�ډNDV�І:���o�n��4���4X�f�:��N�]�����7:q.�����É�c�z�_�[5	��kj��k�N��]�r�������B���8�PJ��i�tlW/{J�}> ����,����s�Q���,��eAAK�]�;LW5�x(y�f��^x��"֫X�O�� ԫ�X�R��C���qh�ց1_�p;҈lt.p��f�B Q�����\������IL� yd���_L�a���BA6c��49����=���hT��7� �]��G�Wϒ����e��p�ܟ��wg�eI�ܶ8��S��w k�8N���c��_7fӤ�'��JnU�6��3��H!/�^ڞ����Rm�L�akH�1N2��Y���A!g�v(��ӯ��s���_�Z1vA��#�94w�0��D⮨��޲�Ȅo���4��=1�X��u=<���'�um����gk*d����"9��������Cƴ����,��1|��%{�x^��n�}�s���7$����b��P�6�a�!���9 F�?]9:U(�stH$r�ыNd�.���7��|�ƾ��}?�"}�9�,R�@Y��6I�����V��-;Y$J���0������m,9s�'QD��Ҩ؀K�����t$�~�K&�M�a8��B6��� t*#U"�8�&0�
�틇�OGC� Y�[�-��>���~�$�#H �V.������kH�-��EN���"x?i��}���A�b����h�;�2�&'<7����<\��~�pر�cЙ��-�B8���O�]�g�-\�XPɌ�$�QC���L)��2�1}�`�18�x^��晽6! @����A[�2�5�c�)G�,
�@���w�5� 8y���Ն�Ṟ'�W�͈�=���w�|Y)�}(��gU;��0��O�ZZ0�w�z6cp�D��@����=�lok����-S�Xt/��8o�}9�+��Q��,F�mE#��g��<i=��#2�9� N�ow�R��X~�������{�T���~}>�������N�6f��'<��p�{~�-��50>�8�r��F�>;��I��S����J�%sFV�Y�,���LP��|gs9oL!�!~�i�;�[��6cl��қ��[r|��}w���ǝ�
%��^����.��P������8`��Al*?/���r����KǾ�7�[!��H���hl�f��õ���L��t�ܣ&��ȴ��TcE����E�n�-�6���@�ާ�/�4��V;��k<�x����t�I%J��k
�����}��=�X�l�����?�;�MQ#}5[�^��)��m&��-�)��_�T��i6��!�𘘝!A>�.Ȣ�%=A0���9�M#�E��D9^O,�XXv�pŨ�\�:'E�Zn�1AC�	l���}�����N����s��?:4�bj�vFI�#<��ͅx�
*��dV����H�BLݔ��,���h��.��<|-��=���+�׬�	�
��%��@�Zpq�������J��Q�@��<h5�	��#)���?	:��ʧƼ�׭Uw2��Û���V���,6��)����0�kv��o,�Ӕ�ٴ�(t��.������1��FRh����zKJ����w�9�X[iE[Ogb����hZm����v�;���G����殕'3��D�:�fg�K�������{'B��~]Y���ך������P��YX� �1���R���I����l�� y�ۡa�ӎNv��O[��{ �wFt�����%��4�v���#u�K4�j��M��F�{m���Y\��OG�DN�bb$j�`ah��o|1>=P�s��bW�����H��.d?`4�D����n7����` �J��>��:�%f�ʼ]�=AÍB���a7gv�6�/)�A}Ü�h�H'�%H��|B�����tI�Cx0������fQ�G��fx���s�c�P	�������A�9�g�����4|���d�
ߡN����Zr�k��dk�v�WoS{Hi��='�b��ڨ��P���.�N�擏r>��?�I�?��UA�)������B�@+��R�t��
��X�rl���gw��W������(s����e3�V�n��WӍ�O2E�Yissϟ�(P���x��oqqE,U� �d�T��R �=tW��&!���ss���Ǐ���,9=̉���w�t���%^�])E�n�W2DUo��Z,�.@1�N>�T���9���"=��Rm<�4�b��=�e�)�N�p�����c3���oL���i��03%�ݞc|�N��_���6������]�&R�=����ҨZ�&,��Z9bpk)ݭ���L������u7�sr�^�&O+��*^j�"�,IZ0���J~c�	Y�1c��
eA !�5z؁�!�Y�����B5� <�$����մL�/d�/!�"Wc�	#��D��6y����_,������G��w�B76߾O߼O�!z���7i�Npq�B�yd�ć7vz����kF���!uLo�-�;$@5G1`����{�����a}��D®BM���[ �7���TV�f!��\�_H��F^���)���0���G��?{:�up�����I���م��`:d��"���@e�y��Z�/���G�=A�'���9`8����u�Su�j3�i�$Ŷ)mà��C~�]�*�~q�+��=��؀[�R����hw�Q�s�\��Ű�FE�:�ڴ����D�'� Giq�v���o�����Y��3Ց8J���Ǒ�I������]�}#rf�[���#� T隔Xr�Sq��VT�*�o��G�mA�P��٭��a9w�������~!���~r���w �̭���r}��E�7|�����-�-���w��4j�KCߒ�%͑���j�r��>i;�5(8l^�b�Q'!���Mڿ�@�	D�xC����K@!�ߺ�Y�ꘝ�kz.=����od�� ���Lk�3\�����=>�v�i
�bہd��?]�b+�=��B�~*�.����92���X��&���wS9�Tĉ��㙢�ڄ3I��.t)� ]���B�"ᕌ�ޘxY8ei�<����KXu��5���Y;�|bB�81AK�[и�)����m/����*7m*7N�T<$�v��Z|�pu&ڂԀ��N�r��+�����U��������3�܍�|��
�Xo��.}JF ��̂Q��<��Ylg���s%���l�D���l���;����ГVL�k����pu�N�|��<U�x+� ���=Nzv�^>���8�8\Ұ`�ɝ�	u�65l#�K'��!2�m#��*fN��(b�tC���'��X��Qf��.����}u��"�|�زҡKDe��K#����4�E1m���H�c�ٛ�^��(k�_���޹9>e_J��(o�zQ%;�0V�j�f�i�����]�� m�R��	� ۽QPmY8�t�\ T�y�$�㹡�v(�.L��l�
%`ԑS�/��r+����L�Z�fut���`��e��`�5f�g�g�(��?�s#�\���0����ȴx�%G��/MJp�	�e��p�#�e�-������ߌ�b�3_��eD����%H�"6YW���H��aj�fwDpS '?�����>�YT<��	p��!�r,��Zc�T��X��0�8a���i�O�_G�p�2�5�2d$��BCm��:L�7q{� �����*������P���ۋ�չ}���iK�2�\W�ZSM+�1��uW�w*����B�IT�q��#�V�`s?qg���M� z�JbL��`����e��4��Wz.7t}��0!ͷu�e��H)J0�CRT��'D)�����;,h����r�u�n'A9���JN2��NF]*��e�3�#Gt�A�E�u����y]�E��?������
$f37��Α�n�� |��<,�;m�*V٨�ŖO%c�K�f7Ѯ8p橆ăy����M`��X���L�8K��͋��	)ӣ}��9$.���o�V8���	�+����F�#��Q��ƥmpv�Q�����jØY��KCyi!�.���<4;7O��%�Ո{a]$�I]-9��{�#�p��ϖQ�J���~�<}'��$��U��<㞄�ٿ�[��36��mCJ6���c�S��Q>i
PAe̮O�W��<�Ć�����ڞt��(M|���{7�0#�1\I�~>K�˒�g�(YC"��V�|������rfѪ2�t��UGE���=�Ġ���Y�� k֖���,�c/�#�[����;푊Vx��YO[t��%U"��DX���u�t'��%8嗲���VEA�����u��	2�]5�T�#���a�9HD�f�ﮕ1����g@l	 R�wF������X0C&"X`�i��w�?*�F�h/"��}��j�$�|�D&�q�I^�=�K����܌,?%M���`/�]��Irz����௭��SV#�JYn�I�wt��
�*�(�Q�@��3�r�j�GM�Z�����c��P������U}���S�eC���u~�zЁd�NT�l6F��+;Q��Oꛁ�}�D�)8����z򋻵a?3�n�GF/�ȬOlT������!T���(��a.�� :���2�)Z��'h3��(��5�yvҕ=��"4+�>랐�Y�W@�.�{��V	�6�mp�
��d�d�rA����^�c1,T ����x/!�����!_��COG?�\{���OT��Z%-?��/ ��Z�y�;QS��B��pp�,<��=Rzz����s7���:nCM�V��	���n��kj>i�
������ <´`�[˩�U� xԾB����2<�WUTRNb�L��j
7s���Ǝ�1�py��;NTNC�����)/�>�`DY=��fԦ�*�M�G����D�PS<BC�`����l{|�@�2����:c!!{�NO��=���l�?�	eXf���y�� �&�h� L-6�_�L�/�����M�ܝ��[~���
�j��Ԍ2dW�2��8�k*gX#�s�{W��d#{h0�sx�Y�o�"�u1��q�[8�I�����/h(Һ�/g-�N���!�XL��b�e��6���{<�������\���9�h�����4��Tǐ�����7��'j���{�>�?w4��(b�_v���DX��>>���#I|�5뭬u.�M�װ���x�LJ�H�XF�wf��c��t���zG��RD�od�&сro-[�^�Ȑ�m����[�n!a��DP�X���	B7���S�{����0�/��Z#�؂��n����h���=�l澦�TE��Lװ`�r ���M�9��-����K�>-=/*(�Re*�
G�3���#��_ �X×w�FJ̨>��w%�۲1se�r͔j_%e��M�	05����6���[��Q�J���Y����T�=i��QhL�+bJ#�-g�8��o�����l+���~b�2��C���-���V���W[��C��<#�9.���h��W `-6�0o���TW]�t}��wB�H�vj�bLB�	p����_M%����DƤ%�^�[�f��4�̒B����"sz�I�@L�NDG��cnJaG��P�#͜l\��4Ў�+�%�S��n)�+�ł@jB�&@L�*�k��Jvk��}�$N�a�l}:�+X�<v���Llbs]�6,N��7В�s,�������I�ZGr�q������2���xvS�S��5V*Y��F���V�02ަUۑ���S�ؑ���m��O�";��2�D�X5��&b�$�;�ylv@�	J�ag}�Ǫ�U�S ��gM��+�)�Pr>D�zQ��l��\=b
PW���_3�Zh�O�I�<�շ=iE����a���O�f½y;��
[�r�!]��2F�z�
��O����^fwK��Ɠ�E:��I憂�>oƛ��?ʹ���.��UU�_!J�|�3���T��Ȅ��XS�C�A��9@7H�}�%���Y��&�)�i�a*�"���sAl�b�rW�����"��������r28�ht�w�M뼹��c<��r���K^ ��F5��(��ݫ7�-T�	�D��<��a H��4��A��t��z<����ux󓂎�۵�4��>��G���<�Sjm*�ʚM����TV���o?���%���L���i�xǧ���߮41E����B�<|Ư{���]�:��W����T�.�<�;x� �,3L��Vu���\Y�N����n�U�����&� ϑ�}�Nx=lc�-�i�/	���x|������;n���%A2�ρ5�f/�0� R9u���f������q���;f�x��l�����-s�[0C�`���px�Nx�3�mU��Ⱥ����A��}�	�*��dE87���o:�@����;*V�mO��ǽ�O�
pBd1��]v�y��f�Pα	��)�*��m�@#��h=��H���1L)p�NL��ax��kϿ`�� �ǯm~�����+�ɐ�> _���mo�~k��ίZ  ~�_zY�#��I��s�!����`���	D���]]��S�m%�|���qVk�^�Fb���ͭ���8&�{	�ƽ�&J��MUtr�ko%F��� ����N���_]g��[��hgo��+_�����&W&ј���3���dK��V*�4�܈�f��>���84��P�x�)A(�G�^�*7��x�\��	�=o<�����zqŞ:F`U��$���-�����m��a��ı��I�I�:h�K`�~��>��d��:M�|Q&31#���Td8���
IY�b4��\6ng@l���=u��>�/�4]v����Cr�mA��4+��8�eO���/���gb`�%B��9���hp��D8s�Hl!�)�8�%�1�������l/"�`ْ%���?������������޾HTt�itq)�<�J���n�܋��4���ڏ5�.��9V?�	��7��=�?� 8�F��ky�W^�@��G�.X�~��ߥ�n�S��FnT�z�Ŝ1�}��3+��r�� �jۉ�eq����jڟ���~ZO��*�KbR�^��D#p��/�&ݷ'�o�Ӭ@�*��=g��nO8�w��C�̯$�|��H�L���J�'��8>n`�����ˡr�����a(����9�$���˼�5ރ���sPm$�T"K{N�~��,��3��u�H��	�U7�t�Φ��y��چ��lj!c�rɳ���o�IO��P��"6"�L�bs8
^�F���	�n�u��๘*���-E/���,t�����7����g(�Ԕο_���R�w��z�����a���<��+c�Hj�R�Y,"BE�Fv��C���H�K׏�(�D��E�Ð����s�/��L��'A߮Sv�h!R,���!�:�Vϳ]��Y�!���B&����C0��F�@��Q���;xɚ8�sR��GNA���q�����b���S-�ɟַ^2�+�|r���+\V�z2rY�4��N+��朘>�>ùąc� �{=�.��V�%�p��]�����K��V������h��C��rW(�?:�w�����-㍄@-.8k�������bPukK;��L����5��!D��>Ӄ�-���d��V�|~�'���H�M�*4d� ~$�X(:�Fc�l�%{%E̯~����I��a�gZY��s����>��@���\�#�*��hP��
Nͼ(��`��	.�zp� � qr����Cl�/|�ru��$����Ü��<��~��>�� ���;^)�<Y�3��_pj�,��ݥ%�[�U��a�fE�����c�,�"Q3 <,v�^����kx�B��3�,���)^��#�����g6�����;�=�8$������lN�q�U}�+��,�ᣎ�4 &��1�JI4�j�v=�l���<A	�������G�f.���C����6m��]`b+�r��Ǆ�<ʫoT��;�k��/��3�^�~$/ª�7^ѭ���)�:P��
՞D�F������O�b�.y����W���*f�81i�bH�ւb�_L�D6B����giCy��9+�Й�F��s�`����~=�r�Mf��x��H{y�9�*wB��龏%��_s��XO���dS*HP���c�t�QS鳴�x�oY'����C�,Ѿ�O6�Q�{^X
os8@pY�j��!�*���1�����F�9�G� xPNw`����־�Y��ﻌ3{���� ���n#�a'�	����)A<��S��ٳ	�e�d�[�7D+&K���*����i���G��&r^��4�������7������C5 �%�Q��z�7csJş]t�c�	�d�YnSpÄ��a@�{���ܩ�����#'��f�근�@��\`S���{��H7��	Ӝ�<�F�� <kXʙ�����0F����0����1 �/�����~Y(/
B�>��\s�}um�z�Y�2��|�*	"�HΏ�1��J �����H�B/c��E,T�텕�q,�����C��%�����ة��b!��9�fϠ�zc�_!\�~B�{ϔYv_�o^�!�������F���Z������U�o��oՀ�Ԏ��� �0O`Eø�J"�^z ���+�+p��*���+(?�Z�'�n­V�+�1F��j�p|d]P�9/���w�R���2NI���&�>�����FD�! �1:��8-.T����Y�箤>��_IMº�b|�W�ג2��SYtӜ��|�������ϒa����Y�ʸ^Mܢn���T���ˮ�g�BqW��/:�,m:A��7E�<�=�6*pi�#����۲�S? ɏX�J��/0�*�(����)����Z����p�'Ⱥ������n�V>��F�K��S:� 6̺�v��	<�����]��Hx7���l~C���l^�u�S�n���M,_	�rV�����J�?�m��_���u(�i�8�D7��w!#��$��{�9=�j�b�fZ�Sp�t�0(���Ⱥ� q��N$��5�K@�;^&C��S?��ƔBAsB\�lq(�ĝ�)	�wo��������*�{mkCz��'�]�����'����}�q��#^�х�iF�[Y�~�ɬx��X�xϱ�ry�/�0�\0#D�%�O�
��ڬ�b?'ϱ�DSc��7����;�X+y�L��:}���8 w�C�5cw�ؒ.M���7���sZ���d:ѳa��*���L�Y¤�����X$cP���S������A��@�y��z�ce&WM�3:�H�G���՘�$j�XO�������T�AjM�:=�`-?iM][#c�Z�|7�3i���UQ�.[4�ё%��9.$�Tk�c��b�?�4�W�c�l��=��븪CU���l��Zh�E4G�v�oٚG���`ª+`Lr��έ\,��Z�nܝWr��n�� �bp�h�	��Ӥy�dI��EN�5Aͳ�u�D���X�K���K�3� ��jt�P�.���� !ɇSIq�,\o�ߘ>�=NZ��q�����zI=��P�7����c���9B��1_���Zz��a���\�Bl�6oPv5������}\Ծ����<H���� ��#�g�N�����@�F�h��{��0�s C�YZ�5�t _ޓJ��	���ø�Ѧ�k� F�,(��%�-.}|٠�����DHB�)�?�d��L�GZKՠ�-����@��9dy�,&��<�*P|Ͱ���'�:�"Ƃ'D�?�����!��p�C@}��������>\����^�f�$�s|�{�Ȝ���dIv��yY~��g"�&�L���5�R�{h����������5��n>�=݄$=r+q��1���췘#b��������O�g_m>���?R��e%4Ӡ��&�Q���{Ըaǀ��8̈���-z�	�\͠S`�T:qџ�� �=�#[���`���T9�DUM�����0�͙a�RA�������o��_�8�'0X��ܵ>�P��U��F��x�	��F��"�(��!l*$�ZQ�"�EE�bmZf�Gn�2xM3
�q�l�*�$��^��]#X���s�.W��NiX���|��.�6­E����Cn@
0�1�}�>�Yf	�s;ށ�Vw��  ��G��H<�|�,#��
C�H�#D�1Pץq��i��2���/'M�0Ƒ{?�J��3/�ЕM,<D`�}Ϧ��% ��S�ܝ��s�K����v�� !�p(ʋ&��e�\�>}>� &����ˉ8��9���X���u��J�u%19�kr(
�P�0��1#���&>�"{�r6���CB���F�H��S�Ag�#�=>�"w���ei�Q�p�[oE���I�H�)���p?xJ�����6��*�oEƲͧ	������kƶv3! #E͑laʩ��jx��(=�Y{���ݳ�K�;Tܨ�%���Nԩ��7�>By*�.|>���[ڍa�]"���F�e�W�fj1֎�GR�,��,�o3}*��Z���#�����R<��RP�\O�k[7�P��\Cp�R[:�t��-G���olr'x���>`=�>�pП����<�;��e%g�A��9X�]��HH�0�n�GOZ���XΚ�}��+=���"I;����נt��+��sE�e�'��U����uw�p�f�'8��$��<����'�\����Y�����P���W'���[@�ƭ.>�F5X�Ϗ���kԾ�'���U���^x�#�u�N[�ˈD��D�����8���v�w�v'��D6���~�U�n�@=��������X�
�8����!�e���H�1��sH���1�����x������pz���G��➶e�mN�I���W�8�r�>�d�(�hz���X����X�
i:!h#<��	Hk�bA���v���J���n���"XX�����>� '5�T#�~e�kd�1TêV~����bI������A^FwC+���.Ç-E}}o]�����[���,	����6�'�i�p �ag<�iz���U�$`Il%f(�@����s�ú-�Y��ӱ�gk��'�|��yڿg�,T+M]C]D�,7�@G �VQ�3.^|�[�UWJ��P`]��r6�bl�%����Xt�/���c[e"����~�5��IPpd�o��%UP��DpΈU"�I�W��6V��b�.�ܝ���jg� ��Q�y�=z�%�׎˝��w�~�~�u�Erg--�&��)˱ɡb>�͋.���N�-�t�����f� �k%�*6�{ԯj��0�_a$c���E["�~�z��� ?��%�q��_7�Wg%���P��.������h;����p<'>����+H���j���g��J*!:?����rtw��*��T\��l,*�JD0�x��$�̗�̯���M��IM]#UtUش��!�;�����~0-y�^���-Q`7dGx���]�4��ֿ�Û���[狀��D�UY�,��M:�gk��6}Tw���(�󝤻���{�=��>��'_g�����u9�RB?fG�>���OF:X#������?fU������n�`����3��̉��4ާtSЛ1�&�j!���\���Z8p�+�{��~��;�[�DŻ��|s)&�KѰ���Mݞ��p� �e�-�Fܺnݺ��h��9��]F�F��I*=/�h��o~�*�ɧ��x�ަ�y(���Q�Q?�{�f?>7��k����Y��z�M�=��yjOJN�̸W'6��ym�W����9��s7��#*^��0���d�M���h
ZG��9KoIV+	��q^��~����D^y9��^�P�'�ɸ%5�d�t�{������Z7M(>c��?	�,���mК;��y ��SL�¨��]�g{!�鷲?ǃݗ���=��9$�(����T݋�t�\�p����~�VS;��࢞�M_�� e���B��\�� ˵��^�ڹ�}��E�}m���J��vN��y��!����1�8f�۷DZh]l��/h�~)e�0��(��U惩�l��-^�[U!�p�Bc�w�*Kk�Mq߮�D�dN!>��ŌƤ�T!ZzdPs�5 �-Fۈ��1�$��ɝ݊����ĉ��8 ^\b�sf��4�~�����s������**�T)� �I7���l�n�i�$��pU����i�I�2��E{ɸ�D�������cyw�)���g�$q�0n�����C�׋�v\鎏?�,P���U|yL3[t��c�
�O
w�y�b&{d��;Z��g��fc$�J���g�S4�v�Y>͵��8�M�4�=srߪK�}�G���+���)�Ϳ�)oM*�:4��9�Z}�4��q� �(TI�̐�҂JW�U�hO<����l�lW,�X:�����3WAU��� o�~Iu��4�o�
�!�ǫ�t3�W8���?AW*������\['�*C�ث=W��o&�+u���#�<tF� q�[<�@�Ӥ�I=7r���3o��y谛�B"��j>��7g��O��� N/2�,�XR[4�:�� ��� *��`�6��V�-��`V\���GK�Q�r]��Ô0��P3D��"2_c���t��E�o�0T��^�V�{�5��k�h�2�NT��D�Ì@��$�Z@���=�}���f�%K��$s��6��`|�h7,�"�h-W^]�ws���s����i\!��j��t)7Ok�J��ӂc��o8�؎?[sA<#��/�2�Z�g�Z���e̏���^T�%�2ΚW�?qu�s%��~�4�NM����A��W:a�7څu8�ܶ��ţ��,l�}/G���N�w�_FJj�mDsϣ��E�}�W���b�b���|1�I�J���Ti�rpАØ��B(��D�@K�u�����6�6O�ᔽ\^}�--��T_��pk$���d�0�{�zǲ��݄lT��6�i��sR�����|���Hhq�!t�d �61�"\�����v�����I(U�B8� l�z�'�a�����/xQ>���H��}R;r�}��7� E/3`�����б�Sk������bS�?]�2�����x�����,�1S���o�����b��t��;A��w��$�u�Z��s�Qh>��l�m�P+����}��-{@��[D �:�6���q�f掽���o!��ND�D�X_���o�X��D���JmÇ��B�b��5�!�3�C����7��8Z~y �,��#�a��H���g�u�;���1i��b������ޝ��X��.&��ʇ�2ڀ%��^2i�v���~;�������w��j1͢)�5��6�} ������kP(���g�0�t��Rj9��W_�12hR��S�S'�0؅�a�,��A�J�F��v�d߮���2���n��b�T*��#l������0��C>������ּ��4�m���l�H^���?�
��z��	{��������g���S�Z�(�����a@.��h^�D�~C�ע���{{�
��$"�v���'��Vp>�te/ ���kh�T[z���I�y^Ƭ@��E+sm ��x�y�a�x�1���l�(�7m�D��b#�A�!ƣ�������6	%5 ^g"��ey�ѥ֍��o�VQ�Ct����0�$3ˊ!)�c_��<�b����@��و2���j`�K�`��c����>�Sf���L�Xv�#��)��\�U� `_%n�w�B�3����>�!q��X��H�r:%�k����q�Q�5�!��0�F��^�;�>��܎I��x�5�6�l�����߄��l���ߌ�$��)�"8�P��k Am%�W���<���~�=�E��Y�;D�������G��_��|sK�*4�b��=l�ZK� #��پ�rb��|6)ػB4��:k��^���MePt��&IRnG�������z����X7�-�:�@��֕\ը�b˘2ڽ�{@	;�K���(|a���R��g�7,5�
�<U����̉�ؔ���u���v�IP�uՏ�u���B�b&�G[4,���
����r�**�K����G����(��@X����..ȼ�����̴���E)����%R-��?���j��Ӹ��\_K{R`Wg�!m�~�yeBz�H)~����k���2��߷��u$0�.������̪�`������US��lE�Jm��-�As��>������t}���Q����ʬ�S��N� �g�E���: ��H�d��Z�[6Ϻ¡[�/��A(�P�~)OX���G�E�S~�P}%:�_�4��憴h'��Ɠ]�ǩ�C��{�:̺p~�W1������S<�ky!e�+%��9D�ޠ��P`��;E`D�/�e��`$�ڭ"�w��{����T��{!H�쏩l2��D���n����c-�-�] �Ύ�yfv8,:�3�*���$�D�c��P���r�&�0�:5�@�|];��q�g���A�m�Q�b��G���1g��R�Δ:��D��&앗�)�˭��i�e��ȭ.��7d�(y��El+`,�Xm2�-�WW�"
�RN&�x7��4�#���c����]�-�;���������L���>�D���y ;nx��v͘#�Q�{���
�&u%U���l��&��^���L��C����V�[ik�R�P}Kk�����q����C$��J���e��`�⢼v'ۊ�s��A;�[5ʴ������W�0�o���rɋ%*��k��Q��T�h}gyſ�+�{�Goܞț.�-+ i1��G|Z�u$L�<�����@]�[��\3A]�R��-��yR��ЙT���&���Q�N��w=�>6~�����c͒���}P��-?h�yM���jeWj���1H����-l�>�E����=�Ky�ʪ�@��m��[�uh�{.�����SjS�ލ��S=�IP�y��(�+�o듀�P�Z����	����N�7FQp�~��j��8�,S�/Q�J�pCH>��s��_�.�I=Sb�a� ���_!I˿!��������m�����z��Sv�I��Z�	�p�H�Z�w���q�0����V��e�)��(���+�.�-�%c��=�����{��U,}�U��
is�~mi{
7��;��L�ʆ����dHI^��&^��+�9KN@�q�M�X�~E-\����;Jy�D�3�|3�w�R9�L�����!�hڇ�a��jc�p@ ؗ>����M!M�f9��������[�1���DW.yt�]r9����M��,4f_f��C^�
�?��?��%��F�O<&n�S�nG�Rl�g�EX�G)u�9#�CQ�	�#��^c����*�+�>����wH����0�6_�h�RT��E�K�ϳ���'�+<�ZK�)i�RWs�ux���t9P&# �����\�T�����A��Qm��%�/+\��&���*����=�J5�<~ms�Q��
�PӪVŧ ���䶇R*��������`���S� ���<~��_��O_��s�r�n��z����38[	���7R���J1w�s8a8d��DC���~	����Q�!�
�7����~�&��H��X*�liw3�O�0޷�d���0�f�!���P^x9�����sŪ\=��Y����B<�#�F�C���=���55:�O�o
 `�_�P��0�U����8Թ%n��#LoS?�s�U_�@#���R:&L5�aa+~PVl�{��E�ٜk|�@��&L.y�^��tsy ����u��:iǋZ�1As$�cK���t��
�T7�d3�Sh�.��ӣ�j�JM�^lm��c�k_���Q/�)�p�T�\f�Ye��N��0�]a���xG5#�s1�*$a�ԜL�����"�� :��FY�����6v�%�ò� y��M6��:�j@T4)JF�'�L�bޒp�;Q�o^c>�k���J=wЙb�k�	h��<�v1ω�l�DaE��Q��� aM���M�me��,[p<��
�ē�p��"b�1G��x8�M�r����j�@�����~I(�r�g�=����W])�5��~#3j�
�g0�,\�;��W�Aj"���(:)�?߸�@1�1l:�Z���K��n�D�N~9���šm$A�O/����5�M���ov������f���p犲���,��o�G̋s�y7.�oj 
7�����z�&���o I��������Kos�ˍ5�=���Q�pu�?�H�����F	l���-���+�ꂐ�C1!�`1�@�����ӗG'|���#��[l��詵g4�HpK��-F:[w����t��7`&QEv'�3RRey���eb9/�wl7�7M��]K ʳ���aT&�.E(�%8���7����##`���p�!��7���(�D3�k�y�+��vX<��U�cb�w�;��˂�f�;<��ZQ��l�%�)�R,�!�g�qY����;�ɆIMݠ�e���`'�s %�{:���i��B�W1�-�=����["Au�a��01�Y%�)��iZ���N���^�ů��q���P^ۆ�����=&�,����R��4� W�����-�g)���i��UwK���!B����?D?p@�2Q+轅黲H����I3�:�x�g�2Qw�6�4��O����!�kF��MM8�5]}����"ae[�ן�5ŷ.ωT�$����	ad�YШ���G����&��c��n_3e[�sB:�xS���VV�W�*�V:7AF2�_�.�V�ݓl0MJ�,��q�g��̯ߺ�7�N�����˦���J%�?o��4��8��ϗ|x	4��4:Eq�6u&�8�M!3a�&��ߏ6�cr��@׶l�Z����ξ2��jN+F�����P7��O�,H�AW)��
�vV�?�^W�?A�d���*�#	M�T��~�n���/unr�V������TW׆L(a[����ؕ�L�����/i�H] �@�pK���Ll��@�
�qnp�����^r.���Gx@�fN�c�`$�^�)I��(	�0>C�:�(�Q$e�g����v��u���w�c����Ȕ�OG@'��w�}���������P�މ�;��yI�j�2HIq����|g	�"�����m��&8���	�u�"���k6�oT�+{<Ź�C	�3@`~N!P"<��<�)�FO����*�����n�<or+ �E�z@���Q��ǘ�_�J�%f����F�f��\MWʯ��2���%�lR=5��WLE?q�eʢp�E���,�(��'��w�S���28�Oe"Jk�b�B�v�-�u��B��� �*�ʈ�1���	D��Iȴ+C�@�jr���������}��*�T6��/;v�im��!��2�++r:8����^{���䜥�}NN	j �P'0�XbC�P�b�AAD�<��l��̖��o*_V�������|^�<6��͏�s��`��#�[�Z9�3�MVp���2j�zA��VF4{''Ev]��0�+^����k�_Y4}>��|�1�?��A����n?�^C`� ��,ܛ���-��t���?&02jK�\߃@&@� Q�:�G���c�����8����)\�%3���4�X��z����B�;��Qz�vѫ=�yK�O:���o�G�y��C'�����)��<;���o �,�3�'��=��������_:\��E�p��K��)ܳ;�8��o/|�O���.�j��Xg	��"u���*���Fg����L+���gY�s�e�\��x��?���� ?�O�X����3X�)���J�B�V럯��lrsuSH�B+$K�]{�+�ci���q��= 3��Uf#Xf��rI����u������T��rܓXX�d��fʵk
--,"I%G��90\�%AS�m����u����� � ��wQpԸ�3���6k�5��>����/�EBb;m}�^�!�������`ׇI[%W����z;Ŝe�(�����G�N��	ER��ɍn��dV6G!Q75l������B폤��F���	t��2�\
��y,a@iݚk�L�K�Y�#�ӕ.��`�M>��d�+H�W��N�+4�Ɍh�م�eAR+s�w�Gȝi-%B�V��܂�-�1:,�Q�f��ly�	����Ѣ�#��\�a��5��\�!|$K~w֓ï�Q�\��&ϫ=�5���<�|;v��l���cr�-�z=*��h.��&o�X�-0�v�����NS.���~��}��:1��Y�P�z�l��%��Q5�=�d"��r������i�x^���\���]�������'0��۫Y��F�hU"͵M��Ɖ��~f��Ê�	H1�ѻg�v�HJ���	�g���7��z"�zA~���ڄ��na��V���I�!�E��L|��o]G5�ώU�4k�s=H��h㪍�������=��x�"�x�!���K�˸����b�V��������.WP�#H��?	i9���O�;�w�yyX�uG�y��k�+�2�"<Bqk����]���_��I`��`��=J�^O��rθ��H�F_>}6����*���4�rӊ)"�yɰl����l����=�@�ܰ�k���j���mL7�Ey<��:=x� �}��o��@�$x5��Z2O�1�a1�#��X���׃��L꤃D7��<�f���;ܕ���U�jմ!1��B�opӝPF���{���R�`��K2�!�6&s�n<ŗn���o��\vd�>%{i &b���R�Öeؓ6�v��Z>rg����^�d�_�[/���),l�����M�U�wyM���͔F	 *pJ��9�W��s�#Rp�J�6�@ H�gr�����ր7�y�J
~qx!1���sx�{rq�|ѬN�	l��%7y|������WE��;�Q܆�o
c!$l�np��H�� ��a��w,���z�fzx�'?����{�v}���(���4�m�2��X��\�Nx�WfE��)������Nv�>���=]-2������t�������m�:��~жN����;w0�㨪�=U���V�����|���@��Չ��%K�"j��)M�y��f�����ۡ��
�x�S��9Y�&����XK8� ��Q���H���b؟>�����;	��>��>/֍�`�(�PP����;��,��E�NL
<�gAob��KdɟOs<s�f�z]��|���N�
נP���A�Pʂ��ھs�)�n��kH�9�j�k��yD�U���8��5<��T�lrb� �����sA��<�X%��u��<>~�u�B���@kl�r��	\�v���r+Aw�}h��X8ai��A�*|\�a�q��ء��y��@�#��wg��*�Z�x���z;4��`hWU|��,���q9j�d���ud�={er�L��
�i}}�����s㛢��fވB�d�a�?�Z��Cܤ��Cl�Q�=Bc	!V9����3�̙GA����ĵ�e�c�jy�bF[gGV�S�=HC�2�A�Z����3��sxD\�R=�O�h�X�_��W� �#����/6H���N�MU\��
Ī��)�5�$�}� �%�f�+�|�T�:wf~�~�(O�Ӆ<@��^? �0=��q��7)u��-���[��������,���LA���{;C���ّW���Z/�qy�Up�
S�kcӻ�-���7�T��9�y��hh�_וv6)"B����S*s��ae��8�ߖ���o��]�堑����B�0z��"ۨ'��Vk�CЋ@C�����4P��|�����~8�	�a�[Vկ>x���4�o*ǆ��ƻs<JQ ���5���L�0�B�S���-���D�2N�.����XA����uo�Q�ט�Ӄ�!b�Q�����;��mJޕʁ�]ߵ'�v'�n�%(����Ny������2b���g�jr��	jf��}4��j5��g��iT'��5�!��m;�S�F�
2:T���?�
��԰؀���  -RD`��@���K�Gt(�^����0X��!X���kZ�7[����/��obdU�^��c�Myj&�R���t�m�@���/Eʓ����J)��Ⅸ����3��0�I28A����'�o��MV\o��f��#�=O�g�xn~qQ���i u�W��9� 0)��0q\:Qe��.��~��=z�ꡎ:�o`gi�������ȍJ�@�{��,�:���a����W�I���E�ZcDskp�y�=�vn �8���N�(�w�Ԧ�ŵ�5�.@fZ��`�4���1�[��D�䠦oX�m�uV���M�S� V�@�L�q�@�L�f �����=�� ;� ��6�OLsh��L�_r&$C~AH'�p���x��^Fe1�|��Wn��6x�'e�?�?DǕҤ����۲�'��$9oW�8���j~���e����њ�%�r��>3�)�����4���đ��k��:Ը�V�'��4���L�2Q�@W4Ҋe�r�<��.yt��RYL�SK�������Ƚ�$a����y�o�� B"�����g�{������h��o��+�_�*e߿��gN|��������k����͇_�b[t�(
b�ȩ��;�Nf��E�����������oae����P3�hK��mIGء(�Jg���G��*�Hn��e� ����?#���9��)ˬ~5zuxZ���Ʉm���yxZ)�D�8��e�?�
���~cu�ن��o�ь�_�K�k�i���x�%��P}�L����>�e�H� N����ە9*e6I��!�҅Н�ԸT�NN�
fW��^�_��~x~I�2�(x��+i�Ԍ=��h�wLCⴗwuS�~<'���c����
+(�Z'"s�ut�Ѿ�z��޹3�cٌd�a&jcj��k��sŵ#��a�Ǟ�
��&�Kd��2j��K��7!k��4�4�����v��V���$T<��=�R"W;����ꪇ�.��_��.Z{�i{�&��bY8Uw��{%�dU��߸oYU��#���J��h��a���Į��#R�ߢ�N+ѣ��ȗ��� y֍q�R������x�����)fb�=m�Qݒ��5;��y���
=�=e�=>U�k;��~K���E��( U;Q�>�?v�U1��z�r�Z@�Մ��0˵��MV"�]�4���dh���|�g�ZNQ�PH|��q��{e��U�P��Lh�;��'��w��U�hi�20���fCj�LH0N��Ά��l�����%ܫ�\��S�uh
�1��]��V#�?|n���U��;���ד��,��E����r� P~t�S�f%�>�κ�d���mDm�5��ꇏ��I��±�0ZD�ZСl�ߘ$�id1��QM*�l���c�փ����[���7c]o�c'�l�/C�o6N�L� _='~�6猽�J�b]߽d��T�����\S��)O��W�ڧ�zt���4����$qjgͤ_�[�i7����ndi��n���zB��gA_����?�f���6Ù�!6�+�f!S�%��
�������]�؜��<i)2��z_������Ct]�}��i#j��Tz��.Y#K�Tи�]��e��扉���O���3�eeS7���,�S�+[Ok��M+�ezCs����^�D紥��	ߢ�ծ76_�� u@���ӮݣwH:�#'��*��GP1r]�&��L�g��1���I��6s��|���mug$�'�:���������H�R#0mF�8�����e*�کi!h�x�-���Fx^������S���X�5�xF�N������A�����LI����_���v�q:q��IW8�7`��w��Pq��Q�p܋T]"�Oό]�u�����és��<�ܗG4�+�+�}�N�����!Cj�U=������)�;e�ݙ�;��u���|�����e|�'����v����y/�.P�Cz
��H��K0ڤ�%d�@H�*���8�P�w;����`�����R�m::���|�2�%��q���T�*]�B?uX�{���y�3I~&����v��zB$�9}���e�g#c�+�f��7���pL�f���2���.���V�	�T�?�U�F�N��f���mtx៭g锎cF��Q������2��2�>�&���8M_ ��4�Nٚ��j��$���gD�F{���(��>WSSsqO�h<����"�3�N�N��k��`�n�a�Ho�9��фj4���GT)(Gmd%��稗��T/**�1���`ڠ憡���!c&�P�t��<A��WM���p� M�:�E%j�͂�����ܸF�w��$Y�^�&KMYd"�b|����χ/e���>>bs�TZ�Rė���AI���EB@x)#����������D��i�gI���-�Y���O60�f��T��~I�Ǳ�B���$P넦�c ���; ���#R^C@}�z��S!�`�"8��1�tok��]I8N]ˋ0q��oO�t{U8J��%sQ���5M�w���Ͽ�$��/>��D6���݌,'��^�rW�/�[���
��@d�li+�Gi�-��s�*�Q��OÔLo�~5lY��\�/S�\ӄ���2�k!MMZ�mh!c���g�~"*qJ+�,� �!>o��gue�N�"9�i�n�͸�Á뭥����7�e�4��x�B�&3{]ek�v������w|4bo�*)S]V�(�J�$�ZL�|���1/~���K��S�� ���ߥ�:�X6��d���G^
%��?�6A�@Xf�vB��y���fM�<����欏Y��A��N砣��n~�KT'�y��3�m�s0�:�/���{o0G�Z�%4�/�3�P�AE�c�Y`�׺Щ�*�o���ƶ�%������+��9���Cdxܖ��b�U�u]��":t�����A"^���J4�헂�%HK`�~����ʚ�W��m�z��(}ݢ�����&4!e��c��L��V M��Zoc�y�\Dx9��N�(�.C���H"��הa!�X�����agV������##Z�/��\=�`�֐A�^�!�2:g�O�닀�W��D�٘$%6=�}�rt��4S�����t�|;KJ٬�!��#�+4�i��7���6Q+ ���_�����oK��p�ލ�0,T��Ƕ�ZV.ni|����a�C�J�SBa#���~i�s@Q �\�&a��,� ��	�I�u�ӆ]����,��:}ռe�ճ'�Ȗ�p�H���������Z)��r�����)��M�mk�� �x��|'�o��gb���Ol��*�s�ZY���ڮc�b�o�齔zˡ��]�U���kM�wt��u8�ýj�v�e�q�s&q�6ʅ��ڼE���oq���b�l	���}tU��D��1�A�4�âЭ0$�� �nW�:Nk����|;�ɕF��}w�ђ��I@(Q�30�b�\�p��_z�?������N�F�����na��������4����ݽ���Q��͈��k�'�+`���}�Xl㘙[	�_��f��\1�1b��k)*2�Lp�]��J��4z�"6z�LE˶�P��Q��xHI8�޹��ƅ��}LO��/9����8qCʧ�I�s�]"�!h	��^x�3�[ևe]�0����h~��p�2���y�	����0}�w8|��Z/��uhŪ����#�u�SY�G�f�f��rg����:�K`���Ծ��������uRe��1!웮�४U��r ��K��5#O�Bp��C��f�TM��d���#�t�B�>�_�6R�m�4s%Ŝ@��$�R�/�֓�p����YM��`��K%��'�߱
�Kʌ�ۤ$��,~P�.�`Zm�>!��<RR9ze
0�&e��ez�4�/U9�)�s��w]PL<���s`��W�)�(<�P��$F���]�����L�d[Ǆ���6��@�t�C��sц.� ����S�,s	� �U����d�J�p���ر�9F�RoA��ga��ls𦊊_'�0�+�=���*��O�)���L��� �&߰�HǙ���j�<>���	�d��k�As���iͧ\_��s�*��c	1#�^��y�>��)#���=WJ�^��U�J��=���4b�\�d���7�j3Y����w�w�rԗv� CKU^rύn�q&2et���S�`n�.��=14Eי����?#&U\��Y��	ۤ�E:4���a�T G��ѱHC�_����4a�u�F�n+4����:j�rɦ%�����A2~z~���\]ʺ��
���}r\�y�:�+�$�2�Df�,۴�w��4_�-v>Ԯc�jHl�jG��Aͬy�2�DA���%��I.��s�!�dW���vkf�j|�q����%%�;ʷ��]+�P�d��}ˬ���|hmn�_��xPrJ�H��*�:�w\�	����q�E����2�K\�W�1��hG�w2�������ӳ�ڊ��h���I�X81i��¸�����t��~��qE�`�U������>���0�141�Ck�\�Gzg�i£ SAH�H&�D����F��xҳw�Y{6�H¸䧉�_�Z�T:�s�x= mH�U	ԛb6j��$4B0G�lը]�*�~s�AzP�3�W��r3D7��ʮ��܅]c�%��6��
���P���\
��z����FY#�� �;����4���.��-�$�yo�tY����_4�8vDl1� @MK?T� ���v�]��� �=xȚ\(�z}�;It;Ϝ�~o���]�����/~��eT.���T籂�[�i�mW:N�{6�(��+\Z���!t�V�Bw;Kx[^������ii�v�&(R�ƾ�S��Q��K�P.P�vR9��(����f��x���v�3�T����0N�>?�q�ɽ�\U��A#@n�vk6.�j�.�Z��&���s:���iۓm������v/]��x�F(dƢQ�y���a�I�q,S%�?�j�#S+]ݓN(s��h�,Nk�O���-\(0���F�N���n���Ha+01�����A����y�*�L�qQ5;ZW2�Iw�H&��C�N_r��D̑�'�W�J�WnC�K#l#��x���0�_Ef����I�%��:f�#��Uf�|Ȗv�xF���M�*(@�����E*�c�"��x�<�3$�����q����Q�j$��� �FbJį���7؜�"Y�9ge'r�(�r��%�ۨӿ��}���r)4��<{������
��Ö<�+�2��/�)�t%�w+�wb��gjlDL@���ڴ){�UA�\��dG���`�[�ߟC�$Ҟ� �%ŢΩ,����Ʋ
�4&mS��CZ(�B$�]�z��;Y�����#>
k�k���T!%b��� Բd����0Q�(���d�'N݌�OHh�#\˲d�H�Vj?OJ��ux��LX�J���<���cw!�f[��ܦ�$��0~�	���4��vv��Y-�O��M�˵.Nt�1]��,=yu��l�Qu]�L&Ð/p��O�pw�BsG*t���}G�6[������� ����0V�R���4���/"Y�ך��V$}�jcmuϯgDr�ȗ��D��A��t>��E���U��fu�/�_0�(L~���8ޢ3G��ԍ�7�;v� Í��+1S�ǪCΈ���7�>�� Ƕ���d!�1[_�şR�p�[�E�nC���t䎇�XF��њ+��-t����GAa�NWg*I���������@:�V�1�Y36B����3�	�y��K<�X�|����p��\60��Y�����q]���*3;��D�¿8?�E!�$-���k-�@#p]�	����},�w#p�@u��Yĳq�H-�	�a�*3�^/Z:�ʑ�W�UN-�^*G�Cڡ����I��zfj;�l�ټjo5��_F��H;�F�ݎwN)ߞMd�Ԉ����=8s̏���u�cP��~'�j�9���#�팷�.�8m;68� � "]6 HI���΋3<4k2=BIw�VB��5�ݝ�-�j���[�^�2r(�N'$��b���V��,������ј1�)w��(��Xt2���XL+k6/�  %!�<���5�I�qu�ţyk�qǢ�Yf��ػF��'v��@c��g���a�1��7S�����׈Cx�_��0����y���6�"�r1-����B3xP���4�&_Kv<�d���C��#�g�Ъ��v��;J�lL�K�Po0��Z��c�m �Uy
��St@H�,U�{�[�B~��9ڑv?�[n�j�ϋ� l�P�Cf�8|el���>�H��\���4��Ϫ�����O[�*c`Lh��|Y6K-���w�l����MX5�*��eU���	ǯI�b�ݍ�&�t3KUj{}���b��8l�e���J��ō�D�ڢ�)��l)Cʢ\0&PO,EK�ą9)�8))wy]���R�<N@γࡤ���D�.N5u*9��)�;�z	�w}5�!8e�N6��;��w���mNf�D�J)�}�g��G�$.�*��"O�epFm�0�PQ� ��/xnϥ��/���������[>����Q��T�#(&�;ɛ�X��Ҍ0�n#Ѻ�x��#�^�PYzS�c<u(�N�5� �"F-�z�;�N���g��kt���l������_d8M|c����j�8�<Di `B��Z-��<Bw�;T���D���+&(/�N���Q]�uZ2�!���3rмmA�tX���Ӵ�U]���.6F���+)R�;^���^P]��:@�]!4�K��^�r5�(�夐���\R��GF��{cX,�zm&�M������J��=��B�{�:I+�����>,Lo��3��l7��BEFěg֍�s~���])�|;jK|e��j�شܗ$X��ߊ��z�V�i�,T�z���Ij�X�4z�\Q�+g��0!�є�3���I4���{"��Sh� 6ã�
(� q���9��+���Y����;K���8eK��l6��xZ��gBj6�Ǚ���ͧ�Y��1T] �1���HP�y1��aD.5����~��Unu�I��j��\����O��l-�����B�=�g�%��~;O��:��g��M��58���M&_í����T&���a";T������6��3�,� Mf��>E�����8��Vl�H,;�_N���-b���P͠�3ч�t�{K�5���a\ �w��R��<(��;#�y����g�J�-���q�F�x�yE@��ϕt��Q���0&����DO� <�m�� �}Npl��/N<_!��Ђ䟋{��*K=~��Ve+tD���A��Q�-C��q�\��-��}%����=�:��^[������9�qZ3���|������R��|�Ē��%9�^(�9;*��) ��ԉ���H���^���h���O�(���90��+Ǡf��p�M���O���o���H۪��o�{��
1X=�We!��ۈt-�U�"��FM*{ o�Ti٨��b�6�J8ȴn�Lm�C�W�R�N�wo��E{�<�JV�y��"��P+gCB+=���0:���tw`T	=���/��B�C!|2t�Ԓ�$'�G��K�<�8nG�J&���&=*��]U��<�>��e�!�^�q��-}PqE=�ϭeo��|��%G�=4�:�~��8-�YP�|u���#0ͷϤQ2D��3���^ߛw��- .g����F���S�.w��k��Ԅ�$F����v�}���1 ���'SAhz�i%�9d��?�y]��������!,-͙�'aK?���j�C�]y�`ʐ��NfAZ�B�b�/=ۮLn�
���W�iɏ�W��R��� Sl���LЗ�L]� ��eĴ�jM�h8�H�FR|�I��{Ig�VZ@����;��D�h�-�1�|��=�F�����Jj�}��Er�x�!(4��e�LAv��D�ʾ��:h
,�U��r�׌��{�.Mk�`����A+��zC*�[�(�f_�n ���j[Ⲉ]n9Pi�]7�XW_7�~,#�1W_*
�&�.�s�.X/��Y��^�	�Q\uB�:�7�m�n�!P�r�̅k���f5����23��;M4/�����%�������f8	V�(��6����(q/�n��] 騔v�VH�$�D�|�ricP��"%���ߞ�$�p��f���:{�� ho4�*����>���e��n�Bm��B[ �w+,�z��Ma����O��}�H!e�g�+L��9����b:2G�8�����n��Ղ��7/ϴb��QS�(h�T���f"� 0Z� ��ԗ���\�A�L��L��kј�V장�%Q�k�k7�k�©�����쩍^:��m�ɰ}
I&^6@L{i��n>@��E�y様�u֏�g��s_��~��A��֮�E4����9+�@�W�?"�U���ɳ��Z ��}v4!��ws��e3P���xu�el��kEׁ���PBٔ�k:N �E�S���Ƀ�苮��@���n��4��2wDc&���lu��n���3������H�H��@s(��r�^p㎬�n�xs�6j@p��-*_��=ե⧝*G�k�0����M|�6I���-��ˇ�5�SE���|Kn�]/(��t:	�=8Fk�t�"bm���f�P=������.��^�AF�Q��W�nˑ�=C��&����ۋA&�7�)6
�]����DMO���u��/���iNU�>����l���∙�Y���
�%��8Lo[����t7)��	�@2������<�����k��}��\��)	L���=���܀������]���Xvh0���MR5Z�)�d�	"(���*;l�f�?����LL N\p��W�r:�Y�ՇW�V��(�Fީ꒮�_g��r%�����]^�Q��R>t��?����yѹP]��)�_�7K�����v�H~�?�
ߤ��d����6[VU���^Q�;t�6�*���]�R��b'54�k��d'����U��J�tP�X���5����7�23T��~��?���Uҕr��g�m�J'K[ ��h67h�d�ϧMs��E�MO�+�>&:���&�sA�3���Ik ��y�MyĹ��=� v+m"���Q#$KK�X��+M��a�?\/nۿ�cS5t15V�p�<��L�4�L��h'������G |b�T�?9��B�놛�R5{��!1WB&g��_��B&l���9�ko��U�j��������{
p�An�px��������� �$�a׫��ʿ�3�͏�,��5�;�ٞ�ς�T��a����D��F7CS�@,,�Mq��в9���7w���x�U�@���>5[1���G���0��x��:ϡ�2R���^#��^3񪓉�Q����1�P�@\(��dl\�J��Ab��3�RoGRNj8k��D^�U�ϋE��;7y�D�<Ad�1�t]�b��*�����+�Ħ�B�=��>���R"�$X��7��j�g����'׽��k���gd7u9�:�A��7��r/��>;����%���+�v��h/� ���H>i<EƋƉ�q�-�l�pmRysJ��cW����t���Qteb���V���r�3�]���g���'��S�$�~�4X4�����6����k%G����#�2�������vM �Y���l�}���W"��Â!�x��w�!��q��R�M�oN�3X�WRK9�	�Ms���'-�A`��`2%ʭ�'�n���:�z�_���8��	�|g�mތ=�K�!�g��q>sOKt>���-�;3��D���Hᢀ��1�ᐸ -��ҩ�u�o�m�5�!A�.�ƕ��Ǹ>g��B^'�F�CLj<�6o��^�
�hC-��K=�qB��%|�h��X������D��[�?Ow���)�p|�m Pd�Ev�TG۱�¦I������e�(�DX��H�$����}��cߏ>|�DO;9A��!���O�N������O��*��'�8( ���e^f2ATS��
86u�Q�9���_4em��"�K��K��kղ�iv��o�@������?'�R=F*�HH!<�oSj�dOϦ� OJ�8>��Q���F"�L���[K��	43hJcs/N4���x7�I��.���?�9κ����D�~.��9��z�C��`b�!w�йsb"����7��I�쮧5"���J��h��G�Ѵ�e���F�;�J�G����Py�K��l�3��3x��F>0*V���\=6�"�=Ȟ�Oז��TyJ�MYi����TNp�:_�a�ȨD}U��\U� S˅@������3r4��S��,�]g�&�y-Jq�$겁W:"^������Uw;����5ǽ&o떶���>�����L��&��/ӏ�R��R���k��x�hͫw�Q�+U��N�N�a�?X����1/nm���'�'$�cH�|}�0�����(&��7%'�#�J�qd�(��l��ez#y�&Ȫ�LcQ�#E��a�� �a":�y����f��x��5v�%�c�>*\l�<�� �i��I�_D�"�G�w��Z7�{�h�������.��bM�I�/��-S�u�N䧢�L�B:2���߼]�lm?o�O�\�MP_�ȡ��tbݾ�b�[Diӆ+	��6�Q�>�� d}����S�t{����ZC9쟌��eȩ���d�s]�����C�{�1�u�8�#�'��R�b������k��<��U�v�6027� �u�C�<fa�����'`p
#ğ���G53�t=��QwF��G**z����L1D9��#S�KȐ��$���7ɇ�'�99��R9���0b[�.W����v����H�ϝ�m�U>�׵"��"�^��-k嘉������n;�;��6t���k@o%��3|�r�A��#_9/UJ[�E��%��*�a�h}Nw# 
���<=w\z̋���_I?�A��o�A0�B� },��'%Mӥ��'�s뮮��)��F�/���Ұ��s� ��F4�� �`�H/�X�����#6K�ab�7�IF�kZ5;�-j�q�v�v��$����ll��,�t."(��D����_ m�#)�l|['PI/-?��[�4��=u�v�}���%
Fr�AV%��CCQ;�2&,��*��MD�K��a�)=�����!�ˑCB������$2��c�vב�\T�QI�S��s�n�[��v?�����~YO;�(__E�r���@��z�]��r�����zr ��`ྴF+*yr#��t�+3ޞ�7h�Lۺs���
�8>����ǽ���?I�u<e
�z�a�u�p���m��
���W��y��̃DH����Ƿm�}emo�R��!��6��*�Ľ�n��G� ���.6J�Bӹ?�%A��^���2��r=�(zo;>������sCQi����^��7�8�fc���}��UK��jr�H�e2�(�}�ώgyw��<?Ⱦɾ���ew��)3�1��E{�]h��ڏ�9k�$�U�)�����9�!�Hh\3T��#u?�x�$2d޺�xw�?�ؗ�����O��E���r�5U|��{�kT&�=ӑ��s��H/�H!s"��y��,�Y �VW��9i�ؼQl��wd��b6�,��f�=�7oT˄
 �;�?�l�ΠZ��R�o�K��r˒u����  ���ڄ1������"��u(%Qr�����+����<'�2'�o�MP{��5���X�SUЀ&n�ȻԞ�����xd?�j�m��6���d�d����g?��yk�E�����M�sѕkr��_1X����?/��+-��aV��y�
����,���+�a�z6}�}��I��BޑV<(?��]?Oy���q*�	+�M5�#:�>L����eB �;y�A��-<���pkLD(�!��ٴɐ�dczA���
���� 
��m�2ʝ/��t�is�B�)�pB��	  ��0�,FǍ�{���cp�{BݹOץ`�������XM��pE?{"V~�G.PFtG�g��gí�U����`e`rI;����tmlNۃ\������EzEv���?�1�W�z,�>xR�A��d�b[>*�R�6O�|f�hb'磫�,~��_��jxv�}�ȿ�+��Q]��2ѡ�����C@a����D*:��hU��z��������+H4����Tp�Wf�mh�SH����E�G�p����܆�<�^�!�Fh��1yE�ԍ^�~nЙq��	�H���V�=�|�^��U��9�<Q�c�5�F1�-�a ���X@2�"vv�Ł��O����m2�S�Cr��yVx\�Rerw>6BBml~Zj�e��T��3��O�b\��U�{8��ԡ�נ��6����+��f}�A�UY��@'��S��C���v$bʋ�v/��z����9��Ż���1����Թ2�R��"V����Ոv��"9�=Dg�lOs��O�3ĊO���:�3�������;h�	��e֋��ȝ�>�W0�Y����W\��2�Cf@g�U%�;����	���!
��,E;wo�x�:
q~}���/��7)�lG2"Y���������K���Ȳb���"t�Y�`@��`j=^x�Y�k�����}59�%iV�ِt�k-��O	 ��:���`>�^y���G0R� ��}G��:���$������]�G�@|��N�o����vc�J
h�6a�݈�O����c��!ZWۅ5z��ڕ�k�G�B�i���v�Ytۉ(R�bA��~���A<-)'�i����qPA�	G�� �*�X!�M���Rۂ0�ת��Z�^�ܡ�ɋ�|�e�:��E�(�8Y��gT������t�xA+k4��}]}�	7Xr`�8�K�v~Bnl�[^����D�ߴ��E0Z4�Mn"Y�M�D��H[P�,gh<B�]-�>ʊ���B�)&�������Bb8%n���l�aAaPC~�	��4�gj�{�*'�8��͓ލ����2�$����{(+GA=���ݗ�&5{�0�qP�\pH(�l�b�ڹR+ ����=~�5|��I��tR�M��m�ś��O0�t��9H�V4")�#��.��\ﴄ*X�WN�ޤw.c��B��)r�a�?qՊ*��Ҩ����($6��\[ �B��f�����e��%?��1{��<��	F����O�(K=���)��nC'P�FH/r#��͠��ͦ�"@��7-���|:xz�SO<b����?T�����8Y(�4�ȇ
ؾo��8��Ӂ�{FLd�����]6l�.k9��b����S�e3�����(�7��ŇȬR)g�Y:24���$���}#j*Pf�d� ���k]��	�z@��lD�<z,/�۹"����p��R4V�Ƿ2Mn��N��%a^�<�^�}յ��1�}p{�8�1��k����j�_s�U��L��}�ܷn�T��-pDk��Bbd���c�D9-Uӌ쥍@rl���nE}Z[�z�qۃ�i%���Ss�Oo��X�R�7(sr�4����!�g�&@ъ�q�/0�'v�<I���� �w����b�,Dy�����g%ۥm�q���e7��-$$�<���!uL�x&ܺO:��UZoyP��s_�uW	#�Y���f9����{��۱��w�ۥI�ʔOOI3T{�t�)6�d¨M�0�Y�O:>C�R�m���X���`�=5�����ˌ��u�c�B���pmf%8ġ���I��E˞n
���";Y�H���|Xv��k%g9^�������}w�f���I��pF>v���96Oנ&�E�#�9�y���yW�����Ij����O�eL�O��mwPW.�R_D�'�MVq��+'4`
Gz�&5��T~x��w�^7\�e�W}mT�z^d������ƚ�c�S��%��
��$F�pj^~b}����P��Y�e�-=�Wo��"�@�ڔi�T��s�/�)~�|W.��?o�Q7���������pYCM�ɕ�,�'��bTjL�����,���:����X��ǒ��?�u7�J�**�|�ύͯ[<�&�,�'�Ҧx3�(�|���g�%�d���VT��d�_?��	HU�Z�p�܁���|�0\���׿iĸ��動� l���?�L���)���*HbbBI9��~���d o�&���[Q�#�����Tem?Z�ã�ۢ߅/f]shtګ���\�w&�9��i[j~�~�$@j/\h�
|է���
]LH��6����������(��`4]E��2Iߗ�jr�t�3�8�*1�r�ބ3j�c��g-��5�OU��;�����ΰ�J+q�S:��V�)Ø�2頀в����.%��K�J�i�������V�����|1�'vɧ���#��O�o`��םN{���M5�CWQN�B���ۭV�8��Z���f*����+��f� ݒ��R��X���ªJr�`{ț�-0��լ'����CI;\�=�L�@�!i�<���!�jF����n�_�I�-�U�v,��t����8��(�����̣LG9�?��]�Fzw����)���*��4�..�䍻�F{|�5�z�m�ڸ�e�zC|d:���ek��$�H�o^5��}V`
���~���H�T�N]�q��|��2w��Z&��\�a6$.*�p#��C���̋WKJ�Po����ʞ���Wh-�-�t�o���E���ֱ�oˮ���u��ΞL��\q���Zt
,�Jf�T���h#���ȓ�(���=��[�x�5|��[��yb�ǒ�|:$N'#������ʽ f�zR����-����:�ɇL�ܱ��q�J�ՠx)�Cd�SR�I��}M�чZLֽoR%+�!�q�k�\@vc����B�K����?�������"���m�$����hJ���Xa`-TL�6�=j���L�N,V,���L�s��OvB�s)���z0��DYc v�5ڹu����~{�6�U���<���ˍ/G�h�w�?�%�b��ӗF5�Riq�F�b��`O�Y<t�
f��-�9�63��.�6���p�j�rrd'r������}��Ǭz��]�&�2M���B流e\~@�܄��{�K��UWP5���G�_Vc��5��C��L�2��Ռ�
����]5���r'��C�-��4'��\����$�U4�jD���V��U^7�
�g  ��<���w0��/[A�ί�U�򷸾Ң�M��A�4�����v��h�Yjd����o9�� ��Pf�6@z�C��R��h�r�� 7�z)6G���ƘW����ũ?C�2ذ��/'Ǖ�G>�.� ���U���
x������#��]!���.��6��-0#��Wl��.oCm4�F��ޯX'��Z�#oDb9��k�|!CNd;�^�ѽKiiK�6���X=ֵ�ej�-�7���q ]��W
+a'����2[�܎V���^�J<�n�^��4;&G�l$EH>l�����.��*�"���������\s�>wB�[�4���|��o�Q�a֋7�$C�4��/P���8������^0�Dlk�?�,�5۳><	�M#�oTuf�:F��v�%@V3�툰���ei��p��
PSA�6�q�R�m��b@�?ƚ�g׽�hFrZ�k�4z)^� r6.����'�x�Rڳ�ҟ�E�I�[��&�){>33�ZOE�2rL��9%B����bKx{���ڼ�_w�@1Q�ty���G#�����.Goe�@!�\rfh���{/	��ۥ:1��A����7󭙠�De���P��x����kS<�nT���6t�����}:�h	vLL�״9�̞�m���pˈ�I}�y���
lc�bs9�<��l+��Ϩ�EѨ�6��͞)yMq����Gbȫ�gkx��O9 <�-��0!�����T]�caV]��x2�������/�{f"���WsIw*ÿ����{�x!aAP�̝�m��7��:{�%���R��w_�@៍���x��q�^��'kg.BL�>hYLTU�OD<�M���}��L 6(n�|�Vf����]��S���P�+n�ERg!a�b��"���2iD�z�&�8��үyV8GvN<B�YYp>|'�W�W�����k|d_Got�>W��`/�B��R�w诊�6��/6���~
f�+U���K��i��DLc�H��;E		��V�(��V^�1���ŋ���{�;+9z7���r^_�'����|��|�[��Z4i|�ԸO3.�"_�:B�TF�e�6��Q�|���L�z�N�����p��ݍ:ʹ"(�~�����G�'3����X��|�4>V���X�!	C������]Ѡ�E:����ӅA�l��ŅX������ϋ�M��	|�-�1�>�W�Ý����S�'��L'��|��d����i�9L��qv�����g<�+�Jt�\0��>6��.1�F���Y�K4e������{��m�7�&��?��G ����ܙ{L���j)�>H�,\Z�]J)~t��i�!Z��
��l�nK�g�0k5�]N��}~Ѷ|�6S\{?�����2�@�9a�7��`S39|[��ҥ%G�B�I�Ȉ�vF;�~��ܯk��0�I����tJ���P�����T	xx��LԈz��Q����Z���ޙ���ʿ���Ne$4�~uD���=���a��
}l4-7RqU:���IbCw:O(ؔ=�	`���A(�9�jc�˱�jH�F�����(�H��E/�����&�v��RUwQ�]8QI����7�tHh��ދA�XK�)g�&j����߯�[�Fd`��v߳� ��	�U������,������v�����>j���L�v%d�n�4KKS�͞�|�n���7�;�'��C��y�o�c>�/��c��'��d�O6��J�ܷ���g�N�t�8٫R�i�!�xW���$��N(y�� ���S�P�~�@e�.�=2ˀ��e�4G�����o�I1kUL#���-4�.P��C���Z�o%�<���n�Xf�&ng�f�5����� m�?���u8�[/ɌVoL�����8|{�-]���P�ӊ�����ZɖzҵHڃdbO��l�[8�@Tyxޏ�m��aT�g��F���V̠.a�Y��Ԓ�]Ɵ�S԰���"��N|D�x�s��,/��4 �--$��G�Y�	�*�W�����+H�Nѝ�<�Jw��1~��5f�ł�Ò�4�H�<�	ͮ���{XnK{�ߧ� �u�w6�ݽ��BO�칞/U�Ÿ(R���^x�5��eq_mM~-� xm�8�k�{,��,��ծ�]��}��J�����t�p̕[e�;=��0�K�n����ݠ���K,��ȕ���l�ߖ��J�� �5�d�8�����޻B�\Z�~��N�T#G���a�9&+L�C�y��ϧ��\uO�N�x� !����}Wt�3xN�LŐ�Эz�u$�)�ͤX�%p�>���wk��/N���^_�{<~s�U����h�i��0����Q����L��˵�2��&r�\�$ ��?i�U�&s("��g��Z�yQe�Z5�.�Ǉ�z��I0�����OʖM�ߧ6�,o�/�6H(5yg�<{/�XN�Ѩ��^n^�[�tT,JS���n9��]�w���H=�� _Ͳ�s���ѵ��^���{h�!���&�B++��W^�J���!bT[�r	�q{�C�s�|]���|�>�\�5�R�0�(#C;����x���p�כB��C��T\�ȶ>J5A��a</�/�ٴ�,�ҫm�~t��r��
�+0�Pl�)w����r4 惰�J@;�u��m�lu�7^�)�ߡ���Jsk�Q��C&$�K���^�6�b�n9���|g�(�'��h��&*��F�!{����i�n
+�6n�����B�W��l5U�X�'�b�{���i���,�+���l$K6�S3b.oa%	X���&���Օ�w�<�"��k2N"�]����|��_u��d0�~ �4[���*ǜ������m��uL>S�k�4Ϋc!��^�*��K!m)pQ�z0�@�夰'�c�*hYr�'!� �dS�)Sރ1=��ʦ�M>�l@8�,����f���?�l���I�zq�F#l��%�!�Z��ϓ�U#�ʏf�"N2��B%on��M�)|v24,q���A�dT�A�Y��J��J/W(^R@��E��U�Sӎę���T`oؙ��"1���w���0�b�i�4v�x�U�:xw�٥�;�à�@� ʾ�Z'K1F� If �Z%�N�9�җ%��?؆ߩ����l#�/�s�)xi��"Qn��Z�n܄�q��5TYn�5�Kp�n��a,�sg�e6��G6�#��l�����J�
b�*l02u#Q�@���d���R�ۄ�E�s'
����x�}2��)��J��%gS��˻⩅dY��PZ@l�-�V�^��)�I)6z�����>U;�Y*V��h�jtfЛ$+x��T�I��S�,�jl-	�pk�p����\�/���k�Y��ER.)��m����Z��σ�fS. o��D�`c��ﷃ��G���p�S�O��;��X�=�=(Ǹ������!�]�EU���J>=�Bt��Q�F|]ڎy��tW�=��8�=^J�����S�(��Mx0M���P�;Y��a���"�}�@�܅We���D_���b��"6S�օ�!}�ꀹ��L��奢"�C�����8D��ۋ�0��@s�89OO�Iʋ�'�߅b:br�.����:1l(^I�րu��)+U9MLM�Ѣ��j '0Fz���@nx���V�}Q�-�hs��1X����GV�P|�8�0�Ɯm% �������4&[�˱�+� ׌͕�C`C�P�\s݅3	��!:��2�����KE�� �I��ހ�G]1�PX�N`.j�}�ų�O�Z1R����tDp���!̥�X�K���1����AD��7�['��4���_��vƸf�fS�T>��q�s
�^��pƅ`a%�y��YQ�g�-?6��mL���������K5�m�4)Ob�6w6uI7Q�_kG_��2�~��f��U�^9Dh�]�c�*���Qp��=dǒ��*]�/TN�����iA�!ݝmv�:0�Ʃ=b��֪_!���-/)�Su|��F{�'^V�����|����t�6��)��C�~��'��
3��������CMSOЮ�bp��36���vh4�n��6��/
���:O�R(l�W@%��Pc�䦶�A��/�Y��x�pAR��Ms��UA�ה�;I�KEl���K	6��~���|)�ن��@��b���{�E��Xo!P�
t~�B:���N��D��p>�A )b�/c	��+�^Ki�m�������l�}�TR����Z���W��څ�2g�h��w�]W-��q�xt��A��w�����xn��	�΍���=O����S��?�vD�y}P����/\ʼ��T���m���O��S?p/q��]��,��ة٥!�g����Rg�z=���h�wjv2F�Ɂ(-_B0=m����
�-���>�Ҕ{=4V-k��~]��f6%A�ޚ�GV�Ez�f�<�������8X�_ezI��%�QgZgu2�]Y�V��-��}�p��p)U#�,�p<+�Iڛ�X�_������hBɻ��&sJ�������z"�S�)�ռJ��6��xʼͭ�3����)"�o��4�v� av-�H��,|LQ��5g!���ڹQ��J�
��9������+N�4���6 ��X#��>�]<����C��+��{yhV�p|!&��%�m=�+����_�`;0�
�����q�u{ JE��zY�Tbge�\���@U�9oq��5���s����ާ]���`�����o�i����к)��\�Ffa�W_�6w�1.�=_E]�,6��$8��l^E���sPZ�f��L�R��6q�������` �o-��/'��R���dA���;+��\��`���7vPP�����põ��ҶN�D��:�tO�V���߻��1 �*vҡ��i��||o�=������`z�ۇ�`�*Lz�^E����":�^𹯑̅E���_	(�d�@�dƽ
�o�OK�G�6C]�[��F&�?O.����p׉L@���T�ebs�i�����|z�1z��t��V�"����!tmW��qtz|/�P^���-�N�V�a*��g+���y,�F+�6<1^8At�%G@��m2,�y��N��gc� 0���_,Hn~֙�F�m��L��y����!��B���LR8C7h�S3�h��A����i�j�gu�	<r��$n��U�N=���x�s:[���F�G_�f%5_���P���1��#��E�h�w$T���E͛x���tÍ_�5yTf����N:D�Z��_�x��>^�bm# �L��X?Y��/�����)�s􌜿��+S������@Ϧ����xX��Ly�gm�L߯ܧ��"
�`�2ʭ7f݀
�'J�ݤ�@��[�+�OvT��r<jV��k���&�CQ���(�CS��a�8{��<}��t����b]oQUh��0[9�����D*�p ~� .����`��R}V��(}�/dY����::K�ۍڨ�"&!@��g�EO0�U�0��B��B:k�S����#H���wE
��|u�-�Q�����uy��7������C�/�^���cq�MP��6�POr�T�A5�/��0p�k<�@K\,cRW;�,�.�,Aʣ��c�Uf�V[hV���C:�����������+��:"��c[Cƹ�1����T�'�{��\d���c�V-���Bħ�nzo
�+�rg\�ٺ�����ro��LSՎ�1V7"��c��)�F2?9N�8T�[�6<!�v>\{=��K��w�S��	�kzz6�R������$�vy;��Op���*'x*��P�����z���'�-~��Eܗ�,��84̵��V2|������d/t���x�g�/L�DR�k��W;s� -V��� *l킅���շq8�h���AȞt6U�t���G��g�A�3�-f�U��=/�3[�F�/owtKhE�H)^��l��*���
$�����Jפ.
��|{�7E���R4�����9z~9�ي_<c��ͷ�%�"!gΓ_G���e�� ���z�A.�Ӹ�P�C;�J����v�>�i������H�чH�(�SAD�B�r�!h�����6��56v$�T.H�����\���E� (eٴzVZ)���+��dr��-Ɇ�<��[}�=��:,ʜ)���	�ٝ��ת�z�c`�*	�銘EFsz��d@H�ʱ�5ic۝�c�aQyE7�q�#þ��^-8AV�+���qtvs8�yC�D��0��>����U�]#s8_��s�,m&V��t�Ԫ���J	Ф87Xе$P�A4����@�n�Oח�3"Vt��w
h��p��?��*�}o$���a�U��@��<��!pW�b ��_]�".�ǥݿ��)�(|�5�1]���N圹�h{�ct�}�6�"����	g%i���/]�cl6��7�;d&�:�6�P$�/�+�\^h�lŰp`�Iq�ϒ��"��M�QZb��F���r��Z��4���[��������Tԕ���x�s7��RR��ف)�P��wA1��t��?(�����`�:&�0l�B`��Rˤ��J�R���x �LE�N�7�/Tx��םL��!�.��缇=V �2�q�q? �5i�;�e"W�Z�'����x��Ҳ���iM8]"�81��֣�|̼n��F��q��.��6{�ͅD��؍	}*x�GP�����!]�~�`/Aa'�ߺ�TAr���
р�0&�P��lSY.h_�T��Y5�wy�CX\xZ��ɢ��P�!'ع\�h��:� Y�9��:��ۧ*���<iSm3^xKI��(��
b= ״�$���bȶ����!1?b�e�4���f��p<bd�~�|C�Sg�!����	�-~Vg��.��-����|ط�����=H�$�Q!��()�qoJ��<g�X��t�_�y�5Y�q��!����V�^0���*����d�6�I��󇩨wG�RK��gѥ7A�α�o�8�
Om�0��J0]Y}w�	�H;-s��`B��;)Q�@5�W����qݓ6�"h���SC<�$o��E�W�e��\�"�M:Y��<6Jߊ`G���e�������[�����}"�ȥ���b�V�5~~lYE}I,��̨��>��~h]�ᱶ(�XL�O�HdGe�G��ER�,�Es3a�"4k߁r�E�L�6��S*����"m��I_����N"�	g��[otQ��Z��9�:G�<�=��B�Fn�lΪ����Łz2�j��ͭ��/�hm��4#8���kg���P̆*c�
��_��W��?n��{^1�5���{�����&^8K��mk�m�o_�v�����(1y���Ft����Mc��ˁ� �h;/��<I��l(���UX��y����Qxῳ_2ϑ�F��� G�[���M;]Q+҆��&�rR`Й@��A:���&� ���{
��������y�ivh3m ������t�*�7?6�����u�'^0u
p�,�3��`kɏ	VԁQ�_Б�<�+㵽-#d��7����.B��[1H@��4���R�ϡ�]e�n� ��\�GJ��Vkԩ�������iL����G:Mܟ�7�Jg[(H�dZ�b�B:�`�6���}�%k�7�t���E�_c���I��l"bhG.b�F-^ЋSa���gu�<��ߡz��HJ�锰Fl|������z0k�#��G1�t��9��H�ӈ�G�=BΖ�}�L�Q�W�guӖz�E����@:�ݡ����7a	�,���K�u�1����/xV @���,�����@�Q�tx�K	��UQ��5P	d�|XZ:�Ϊ�t�٪I'��w��W���c����-Ǆ}|u�,iU܃3T�J��Y?��E�6���u���%���&��ap0N#w�����.�zù�cr�����>��<Y�M�ttD.�sjs:\�)�+)� qa/�YÓ_n�y������3g�!y��H&�)iuˇ[��}�ek��cR�=���;Ge�⪴*O��c�%\y��!l�,8O�3�n�u8�n�#�$,���ѳ�!F�喿�4l <VK��0,v_���G`�D&5�~C���T�>0���-ϼR�XtI���U�<��y봆�I���շ�q]�	�Q�t/�Sj��"5���%�N��9
�kG'�kwx�bj)�[�I�JA70�<�|
-A_6�ǖ}�� +��C���-�GB���V�i<�Μ)(�t(��F��߇�%G��[���s]�3�((��D��a3^�eo�tl��hL���W<<'4�.55M�5�^� �`��Ka�,�|��&ӌ��NTڵj3s�Y�XEkM]�HL��n�Ð-�z-���V���!ړ��:�,���A��/�?p����S�Ŗ�X���x:��@<*�DCa> 8c�%����K���[o�z}%8���G�Oy�i�P���9����{,Vz9^W��.:	X�6�*��;Nbx�r�r��S����>6�/���Jm)�أ"�]C���z�\��|N<�SG� �
c��K��X�~&�ξ!gl�(�$T{�P��&W+�M�W�ܕq^(��Ģ�"�񏅤��*���=��(�G&���I41ES_;^��6��W�衢Β�gʹ�Ͻ�P��`�/�r�|��N���x��L�$�l63&���Ͼ�זX��$�(�DW���[9u�-�P@#m�MUi��؟���y��O�my��1X�ZЃ�e@ ｑ���j��u`��&�js>;� ����:mI�i%e۽����m�Cr\~���x�n�r����EA�������ȅjj@�~ɖ;��Tp�\͓L�`�J����n�RJ	��������(�97�8�i���%�>�M@���EJT��.�ZO�����B\�:�f��9�T�-G�h�����n<����r�����FͬG#�e�p�����yV ^I"�b��Sx��~*��f8�f{qűz���}��z��m���;�<:�p��U���@~Ht�$��%��\�r�	��+Ck��%�؀��u��脄���,����[	� j�Z��;T���@ȼ�
�����!ي��W��%O��u��]u� ˉ��JZ��fHG�JJ�%AWK�+�r��PNP'�'�t��������T�&���	�i��~���;���+���Wi��
gC��x[}b�Y��ocGڵ��q2��0���׈w�Z�M�{/�y�_��9�J l";�=D2�,'DnJ
s�N��p"h{���V�9?���}��@��-M�\����߼Ǻ����˷1�k�����ȵ��_�ͦ��s��K*���/"Li<�]��D���uI��VFE����)��=�9�T���[Ή�)���s�Ee�ߐ�$]�/w;.�?FS��ܬ��CI�D �&�*I�H:�`bz�"��0�f�cm�q��\i�&��K� ���zIآ:=�8l��z�}�J�'�����!І@�
f�z�quvu�&'���d�=�h�5�^��6�d���?�z[@��Ӯ'Y�������e��rĢ���yZ�͡�,�}�!�	ekK���W֏2�aw��9�){z	��!>Z]O��gV�>�GD�䊻 �#�R���F2�� 5�z��9�rpF�y�n�b���(CbŸ
��
/"���iX�ht��<%�xe����z�D4��ڭ��5YcEZ��Rx�g��(ޫ��T�	�"Q_:�k��5>��RW��2Ue�i<�0'M�@Ѩ��j�+�MTg�Vv��#�Z�P�.a�q�Lĺ�R`[�ﵤ��`޺�b��>:Wݵ����� z^H�3�ߝ�d{����.f?��Nh�'1E,��'�Ef�R`B�&�S���,�����{�#�|Ș<��v)����.&~�G��}�# NA�D�W>�E$��H��W���fv/Lx�{2A2��P�T���eh�&;A��7�JM�e���$��~'��9�Y�A���Nw8� ����r��Wv���]�����<�L3XG�78�n���2S�E9eI�d���^~��W�a� ;����-	;��K��S"Ǖx�t;Ul��!��/���tr4���� <p��z8 ��I�x��m<����|�b�Ò n2��b@i%��bl�4�u̶_|��:}�B�[|]�f��D(>Z�Y@�6����0[]ҲY�0٢����W�_���q(*�!�r�k��+���<�.I�̛����0�t+o4j�]��=�H�>Ӊp�	� ����������
(1��k3"��b�戁#I�>�}5o�l=��Ā��qrc�F@���l4%D�I/�(0��c��j����Q#~te+��J�Eq��)E�����t�ja9��M�X�lk~1l���ʑ�$���-�� �pE3b������hU��n�~=�����SK�޵�¡�j]'������.�K��aZ�_"�8��|�,���/��b��a�����Y˛	K�R���h@f["fLްZ��T��0�z���50�˃���IsgȆ���`���� _��ʏQ��י�u -2<������M[Hb8b�$I�m�62����2=_̟6�jvEv���3�s! &�x�Dc��2����g7��@�iX J�jp/6(��Y�������;:�U;B#* h�/X~f�r��o�δcQ~ �+a��6l�`�����f �"3�g @t��O	kK�{�]�k�~L�������Z�Lk��}9Y�E�'B�b(���C��\�2�+��G_՗!��<���d�&[9�n�l�h0}ywgtF�_���B8��L�?f�'!t��|�w�.H�0#`�ř>q��_t7F�E�5��GoW`+8T�>������}t��
ͳ���V 6uayI�\
�h�G�(W���d%D4��M*՟ˍ)X��d4��A̒g_�M^����TW��/U]�|K�4����~�4iC��]x}"o���i�x��͸�u�%��n7@��ɍ�;����f��؇e� �C�ک�ϒ��ؕ��&�WR\U\>�$7�8N�\Ï~B�LQ`��`W�~l�ʹ��	������x�1"i����,�Z���ĭ�ZV%�/Xmv�3��	��/���)�*Y%c��kYuTd����>�N�!?[�>�D�#G��	��*��Sy����:We��w�[��+|�dǜKk�'A��Q��p�T~˴V�7��*��c1[c��q��;[��tY]�X���)3[�;���Q�<�m�}GW"%Q�/���K�w~|����f�f\�R^C�����^��,)j�_�'~^ ���Ts���� �,�X�l�w̢�����~�e��(�K���]��Z��C�R}��T��a�7c.�&�[/g�	Hڻ�j�dX	�n_�S��bO���O���2�5�C}@�Q/q偗�ͤ�/r^!Q��R,�	<-�d���#��/�!J{<��	Hp�U/��=��(�]+8C$�$t �U��$  �5x�u�|�4[4[�$�H�t���1�>���R��ρ�����`\z>V]�qFc4�q�;�j�%��&�A�4�b��w�-�){�n�fh���e`��T
q"����O�F5���~	@ޯz"��Wl��D=��߈4n��X"$aD��7�[|k����O$R����@{�o �&9����^s�"���i�=��Yz�v��Ū���ܩq��s�-����M�xJ�`�i8����lcFV���n�'7�)<�"$�o��~!��6�61�]���\^��d�Hx<�:�/��M��@�sCm��C��_��O4XA�A�1��%_a�zI:Xr2砶#F�~��W�&�� �pz;<61��Pυ�<`St��L��N��f�Eb0U���U(6�rQ�� ����k�|k\�S�
'{�+�[rL���Hm�ӗ�>w�M�ć�3�J�&>M�%*v��/�<���.�ݘ�+Ģ.����lG�^�F �NR�p�b�X�@P3���Y�P؂��^�&2HKר�w�7Kfʖftǩ��W��/��QQ��V�aH�Ҹ5yR�UT�@}W��`J~_��1�_G[��ܴ�)JS�p����*Q������'V�w���{��R�U6�v����@x�T�h{�/un��/�P����i������`LC�Y�����1W���-�i�� ���P]����]�ɰ��VM��H,Z��X���M�j��I��
S�xU��_J)5y8�INh���tM���u��II,ϻ���WĴ���`e�^�3���	��m�4�w�M6k,�Ϩ�<U�7�l�����`a!�U�$x'��ȄTS�|+l�0y����@o%��Q�W����!������9����	�O%joA��NBޠ7d���$%�}o�����Lr�´�o����ՄB�B٪��)��as�`E�U�[��G�+^�<m9ņz`�8�ӟ<ji�X���G��B����F?���`6z��5�L}�R��n�VaĒ���y{�LO���<E���Df�M�>�M�x��`��<���3���y�^N�]=�K쨱�Ȥ���#�Aa��`Y��9������i��r:pב�k��g�*�*���Y7⽒g�f�=*��*��vḭ���K��~��C�I,R���!$Egא�w�A�qP�j0	W<�{+�@WҒ�]J_Zh����m!� 4/�~�#�-���,����w.`X�Z?]U��Oc�������O
x}$Pq,{
Ds��V�®�p#H��B�K����\����[ё�@�IA��+{����o>��2��Ȁ�n�G�:7wXJ��'�W��>a]�pN/�
��\��@�D�{ �kj��s��9�x�]�Ƣg���ބ��	q+Gӝ�,�w�S�<�ypg�[(�d7�����c���$Y
9�:N��'�C6�'+XY�0+��$�Pn����&c]$�� �s0�V�CE�(!��i���)\���C!�!�H?F((�/P��웬N�j��;�z�~<�E�j�����MtP�9��]z�����ޞ�:�K�^��lBv��Fb�wxvj'g�p�,>����z# M���6e���"�%�6����~{�g݂1��>��c|Q�¸�j�u㈑��I�/n�W$_�Z50�)/*�Ì�����{���(۳+����^`I��%~�Na�2
�2�D�p���J�O=�H�ջ�n���o��B����e�;��j�u}wQ��'�TU*b`X��H_ri�O��͕? `*,���Niew6�Y]�P,1�� ��+�ss޶6���&�B�z~p䮬��3��f@���l�ZX�X�N�����Ї!b���g�%H��\���`�����c��C�+h6�'��9��xS�#�=����������q�� ��o=;.xq������<NW�4{��f�ԏ����X�'���^"�+x���2җ�J0��� �?�¿ݚ�U�u���,�-�#9��cf��L�w��c$��.�ܡG �;�-����:j�暴�S3��7R��Wpvz8��vӠ�g��(�׳���]<7��Ίq�p���s9q鮧�#[��B���#l�%�Hočs�4��H�(��_~����3�'��8�gb̳T;�gq�=x�4to|���  6�a�o< �z� ki��i���K��>�bv��}��C��fs\�7����[�ӹu��o �����Z�08jr�,S(av׼ϩ}�����;�|B��Z��4���'ˌ^�Ԇ���@�@�EϷC��G�i?�+ز�fӇ�R@��8U4�Y�>X�Qa��S�)R�o����銔%=�N��"A��u1�J*��-�m٩��f؜����$�C��9��of�`����ˬU�C�G���r8�5$���8�1x?�S��nPi>����Xt��*3$O�&6�ˌzʈgs�d �� !e��rA�"]ĺn+\:��B�!4
�g��|�����C�-������*�-@�P��
y�Ɲ�p? ����S6;S�UY��U�S��A��Oi��~�9���֝`�c}ߣ��e&/^8�VF�;pȍ���]+��\=�ɟ�.O�o��QѦ+���I���=��^��@ZO�z�t�Uw�e��}t��B���������-�m�1����5�n�j0-�ıϻ�)˖�Xd�M^Z ����v�*�(E ����W0.�YC�L�O1�n�{�2x󦹱.0v'�8���NG��ң&ZHU!�F~�b��NqLn�0�yV]�c�83�M=���4�� `���8��Qw�J�A�ſs�u|_z?���"/J^����g6�X]6:���F�
�%D����uD]@ۅO����4�z��fO�kKbG��>�D#�bF:(8�Ԯ��7�I�
*�����9�7�����=!��~�(�T�5WW�熠�����+�Qu�́��eN6��|����x�/�1���u&f��J�|�2����/'J���V5���@-�g���b�����v��I#���i�LP8�tb4T?|2��En�U��HU���S��'ֶ51��@������TAφy���0�eƍ%�m���~���>�� 2E�wӃ	<����6m�Gˊ�ŘIq��B!q�&0��i�%�'Ƈ#nw.��7�J5�XU�ϜS�^j>��fļܞ-RO��|�t��ͱP�=�fS���@��������fgh��В#cǨ�5ܰ�)��V-;�5��������ʷ��{�nz���)��aF���tz�	H��,�C�݊@q<��V�)[���*�g�2��A��d�n�L\p隤5������Q����]�M57P#&t��6;���C��~(�xR���}ac/�9�Ww��3��?��+9\<=�y�����;n��j�#�
�M����8�R�����f��^4=_����Je��l�O�"�3S�ɻ����y���eۗ�1UI��`�D�ꌐ�&��G�ɥU���9{�Q9�.�i�����j_��j�Z5���h��bWq#�1�?�@��6��ߴ2�$�dw�5�԰����/A�r3LB+)�!�Y;��<�����E2�̡�:�!{�
-FI�? !
��+%���p`����t�䍃��9(��z�LE��6����	A�}�����������J���I<�NÌ�7P�ڦOm��҉�k-��N(*@q��Tyt��C�恽�㏎���L��$��v8�>��s�n�K�ϻ�Z��Zs/�'�֔�٥�൫1�^M ֊#J
pė��4�xT�r�:��"��tPv!B�(���Eۏ"�9�d]�����1�|>I�n��um�4-rF��X�ef.B$��/�:1�|�3c-�'�q���L�X�F� �>wR_?�ew��z���'_Ǹ�9-Wd4Y�6@�M�r��Q��J�PA��{[�����s���n����0�|KQyDO����x�E��t��o<��	����h�����n#	��CI��b�axue��R���ֶ03Vi�
����s��tpG��� ��������7��ZNg�d�3�r![>�`���� %�a
T��A�K{+��83If�F�ʬ����={�{l�\(�k�L5����M 3������x�5p+�ħ� x)�%J��5�3�����Ej΁k�d�tWb�L5ȶ�	B�u�PrĽ�!!�M�eQ�ӈ_���޻Ն�ax�x��z�"u����l���U:�a�eĪ��j&�X+�~�)���Fv���#nd��+�)
z�ve.��ƊP�e6
F�?��106��u��k��4R�r�����������T�����(�&V�TZ��y2��]��SX!��m%�9ͫ��s�^���u��������8�4�O��f�q�V�dKd�[�1!P5��D�:~_��\�>Aw���(�ڜC�ٳ����T4��q��w�m��v��<�QN\�������� d�/�&�<��φ���Y��	G/��t������<�5=%�A�}���TR�{�����늝��jځJ豜rE�v��>/zN:�������Sybǐ���0 }'�|���c#���<���uc%�z�;ёFS�9ڙ�����rƫh�<��"����Q/=�;ExZB�5�cޑs^�K-n�$!�3$��axE������{�*?�v�S*v�i������r��R8�P0�z��@�e��
�㈿��ΔhkEI'�a��MM0h�ï�˺�|'4�SY(��!>2�`o�dA�i� �I���W>p���5��S��1̤
Y2�E�Oe�) 7�ȢZ���e�D��4x�8�?b�W�G�P�o���O
Dq���E	����z;=��nZڠ�f~��D'I�B��,
�X�(a�'����E\q���	�N�}��	��(�Z3��OJ��C"L!����uNM�e��>���opj����$Fr¥��3#b#+������\��s��俓�!G�Eh�y4D�x����!�/��
6_�9���x�����/>�\����m�.��ēH$�E��l��b��XsEQ�c.�6
��6�4�a�}��F��%d(!y�e�B��TP[&M������k�Ƈ;�2��]�p��vǰ�_)L�{��?C�����e���IhWf�%27��rf誡RL�"A��6	<c���"��c���E�����Y)�
��B�9�ϝ$�~sÔ,Һ�wa<�3���C���2��J��AV�2k�sJ��<�@7T/�no&0�e�?�p�51>@ܪ:/���td*��ȩ�T�+��ӝۗu��W��0�I ۫�*Q�����R��Fؽ���
k�ҼE牄�:�q�}�t��i��_f�]�y�CڇI�V=��uT��v�6�.�L�t4�o�]'Ku����r7[V�|���!�3�`@ō��{�'jK�s�Fw`������s^�}�=V�gؕ�n�*U�������1q������g�M��j���Ye֌�-�=���/F)����M4�'�_{|��P'+$aA]�����6����q|��'�1��t�#�Fr�s!���o<`^k��˔4��-�	ɶ㦡�u���=,���i�J(�
T�_��q ��1N�w�� |�r�Q���HL�~�	V��񉏌o(q��S���%k�Gx{�◬g뢩h`�Զ��iӑ2`<p�)�?Y��oM"�3жs�H�֔1�%���8�w��w�#�ԩ�i� K��O�,��׌8�J�3�E>���2M�F���#wvUr���x�!�,�],%�Z�C�V��"�EweͲ�3o* =M/{��=!����Yg+��z�4�7!���i��&>�����H���8(��w�u�Go��rGt��g{�菟2�V*�O���;���CA�k{=9d����Lt�Rl4��f���������p��0�y�A�X>�0=�Gf=hSDE}�%<� �V2�9l���z=n5oH�;F'c��ߜ���\P���5��ǅ3r��҇S���n�)9yѦ��_�a��I������ۮ����2[�U�����k��sD���Nս�Z�={ќ�{�헭���yGBb����d��V����J	��(�3ϦK�/Q����=��H)��@��O�{{h�C`�QaM��R�=���F��V����"�?:��{<|���Œ5�8��w����y�K/;�+zO>���D��i�@D��hHάq�Xd�����@&�/G����#Z8��%�tA��eMNan�#�h��Hn�_�����o��ʤ��""If�G��q���30�4�0݄þ�mX���͉2%�>3�����5#Ω&�I�[Sl���wo?.U�l��_�X3{�Ks�@O�t�w󯒓��vp�S�j��n�f<�*��KgG�!Ø����a��n��#%ς��SvT
?��FHc7W�Kݩ�E`J@�������~�w6�)����m�#�z��P�6j����6$�l.��*h�9r��ƌ�mi�&_K���\�Qi@&�u�9?��J�@(�μ,�N�
Jͫ4.]��M���u�\kL��T�(��{Ž~-c����C�#��ό!��iWp�.c��{���͇�)2�<����2����͌���$����Te=�?U²a#���A�E��
-�E����hb�<��D�:$�����z��8+q;�K��]�1��p���Q5��j��&��Ԥ�v�٫yn��;u����3���V�M���͔�G]��y���;�����1?����wK��S�gw-��t4Ô1���r� Ǡ�TK�q�va|^���?�N�T�z��7���H�p�Ke2[�v���h���p[H�H*9��pC�
B�s��S�w�]�?,Tn:t����
m��c�e�s��(c�)�7���?��lW��/W\������x,�p�}�dݝ�]r� �l�Y�h�}���[P�����F���˨�� ���!۰X�s��pK���VZ��-��QM���u̖{�[�;��o =���|NJ{���Ŷr��*<�G�lY�7��	�a�k$U^'J���fg��;�6B[���A��]��t��I�|��#R
["6Y�n9�>/�ŏ!��O��d�t�`=������l��Gʂ��� ���o��R�nkl&g8sz[�2��iۃ����f�u����\ݞ|�Y�0H�j�����$f&��Bhč��ө�)�*n��Z�D������o��>[8�A`�.�)� ��#J1�������?5��r����`����+Z������f<�Ѵ��t��u'�`y������BJx�B�,/�+���sԚ%o(�%�ɭ!�N|��XZ�h�waj��-�-�{ͅd��IĢ?	_P��4�feweH 1.�0蒂��uUT��얗f�� 2�i�r�yOL��$���xl��"�fUU ƞ����Dj6�!k����Ef�f�Q��q>�F�&D{a�P��I�H��R	�N��Jn�����x͏鼞'��j�<y�(��SN`u1h��)�n�FԽD���xb3�d"�?��$��krA��Y�A%�3�P�A��.N_�0�V��Շ� ��QQ����k.CY
su�`7mb$��n��VE-�P3ۊ�N]���+VX`�����*�ar�M�͕I�"��[��A`�H!����)SE�(9>/n.�QJ��|��'Θ�c��`����"n���Pq���vڃ��I��ڼ)|��5�w�Hp7'�
���b`����p�����]��wH��bH5�K����>��UbnFnf��h��?7�2�H������1�4�'�SyI�Cg:sWe�J�[Rnu|��
�b1��>@��g]j6��w�E��A��\]r�ꛙ���'y���4����ˈ`H�����A�B�\�(�p����K��!aB�����D4�r��K�r��݇6�ό�1�R��a����|"Nd����~bUC8��1t�����1m�9��J�]W���aB��n�Ž{js��H�^�^'�
�����c����Tا/�����~���Q����B]y�^�Y@��65I!��ie�|��{�}�ڋ��1~@R���p�!�V���i-Ή�l�01*�J/�%�L�8��c������>�xźϘ�s�R���_I�/_��.!^d����O��'h�al-���ί`��v=Tp+g҂���l�C�aE	�^�W���H�#��Z#�!t.�Ӭnt:W���u� g����n�]�2 B�G�Sj����K�+FEH���;Y1�K ����LƉ���X�]��0S�U��R=�V߾t�&J���^U���]��*Yɑ^&Ehh5�|��S��M֕�k��ww H���D�ï/�=���Wu8�{4��}Ȇ�^�U���a��7����BX���Ϋ}����MM�Iq�;�[s��b�n�au��������<�x�+u��&a�x�<���b�]���)zq��z��ſD����E� jE��ë"�XY�l����e�"B[Vw��>#�W3�����<*��F/3��ť<s߼�ڏ�9�k��7����9$�LQZ���Ql����/5(u����턦�]vܨ5ɖ���i$��{�Ztt��=Im�}�\}ڠ+Hw�s�� �^kvG8N)D�}?CB[�2s�����r]31o�}h�x��4%@S\����^T$��"��ba���1������I.N�΁JX�zF.˃����eI�ݷcq�ӧ�(T�)������+WkF�4��G�Lɍ7�f_��f���h��x��?�л4��G,^A�V .�u�K��;bL�e4'ng|����"_��!_�H��\��~�&@f܇��={�nD��p�tJ���e�S))S���N�����d���y,��T�Yl�D������*"BP��3��WNk�J%�d���R�����L�bw��0܄,�%N�r�� ���&/�6;�2삞�lA%|� � ���x������g������J��P�o󾡂)V(���f�_~\-U~2�pQz�f(fȳx�GG�6��>�'�Y�簬��G����F�տU=�K��>��Kl��=�����N������xF�Q�$�'�����/�����R�P�� �����c�� v�&%l�7��8���.N�(���t�y[0 �� r� !���$
��˹�vZ&/ib��3AfV8��o�%��/�Ԓysfa�j���B�p7!�H��jivy!l�@��A�!�1�S&Lب5_ �c�k>�G$����x��]>6f�&-]UU����5��G9,�"z������T�E�!�pIl^�VJ���GبG�z�04�R�$t������c8T��Ff��]�J�t�9Rq����Ɣ#$�w�-~�tڦ�&{^����(�c�C����1�Э*3�o䌸1s��M+a:��w���G�ŗ�U��k��8�!y������\�"�:�$a�RD���;�l�'���1�~���F�f�w����z����.�@����Tÿ��'<�*Æ>��K�����Z�t73�k\�����Zg���)��ÝHߧ��aŒЌK�O�<7��f`u�и^G�8Me)��"�T����4��rFJ����s�W�|�\y�w�Ď@���&2���������Sg����P3*U!����a��g��>v���c^�vןU���0�4i�#W�� �����s�$>J2iT�mY��מ}�5Je�LX��W�(W!A[l�A�%<�s�O��II	�Dx3E=��5�C�.��K(H`��$��J�(�����،�,o�C |La�V�Q���A	s10��q��y�,��%D�<$F}�;���`�꽺LX�x��E���vl��U||�F��%B�^�.Q
����Y��DBT�;���?`��?��F�_0pB
5Y�P�Gt>N_��pP���*,��h��]{���~5���]�=�����.������I��� �:�?vo�]�$,4A,0���J\v����%2GP+���{I������]I���� 4!#�@7�y:	��g{��q�-�2<�&e�4� �i���B����5'�L�����L<�#|�{��g֐;)��f�3X���&1Cc�I�4��=@�r9a�Q���\��l�5g�,�D�����

)��jQ�t �3r�Tm�B�kx�ex�Kԅa��qxC�+�v�����	�Y� xgA�p�c�b�~}{G�A�(�u �ba��Qr�w���-.�,_�-3��a؏���=Q�S����U�!�uwBr���6G"�Rp��ͻD��l�`:O?`E�v�Q�|���?@��Br)Z�������eP��8�h�F �Vt�bS�Aِ���c�V\ч=�S@�����Ͼ>Y�a��-clQ���r�b�큦��4�L0BY�L�B���44Gg�;��`hn4	�'$`S�32&w5�Ne+�f�]:�w����$�\�����by��x����E�<�?��r��(�׈�PW���N�%�$4QooH�_Wu�u9���vJ�ne�'�9�nĥ��¥��0���!9wh0��3�7�`K<%���e���u��M����X�?�p}ʄn���^aT��Z>�	KP�I�EǱ��cS8�U�	I1r��?�40Q,�s~g46�MK��\�%*��#��B���|����Uy$^9*�3R$�'@�hߋY��
f��(�/�����d�$TJ����'+�&� ��\�J;�����*�R���K�e�Uz�d�r�C��'r�Π�#����6}ݜ^֫�SH��w�����[%��}Ub���ʁ����P(6"��J��ccE��}��kMP��FY HD&�;���L�FC: �Xt,#rY
o۩�\A���B�)�ٜ;CL@	�V�Z�i>����0��)mB���Ɯ��A��/��wF�B�{A�h�Q��Q������/���i$����k����90\4g���R�M�0��3p�a �$�2�v�s�H7.��q\+�ڽå|��bB�����R��:��^i�N�;R6)>+p��7���=�#-"VA3����ؔQ�g%\V{��Տ9�U���2J�Bl�D<4���[���,����j.9p�Qv�����CX�:ߋ�Rþ�]ÝO-!)�@�zi��$�#�;����`~���[_�"�x����i��M-�Ļ��̾mi �E-�&,幓�9�Զ6'MPL��fð�}v�U��j�`��}]@�V�#�o�+IU���G|��أ���)�n��u@��bI��9��uZ�J��I��_&(�:��2�v�{����Kh}��>��_}�'�i���%�
>�F��Ę���R��u�^�>���5�����l�I(A�H��yJ�1��dO�N&��2r�;6z���rV�բ�3S@3W��t��m��B���Ec�%�K ����2Yu �_#�%���yG|ӱ�<�Ӱ0b�CN���&CZ�x��M:_Z"S������*h�����S���,��m�.�׭�#���PQ����b�~�)��kPS�D��G��	�H	[L�[R�M��$ i|�w'���� �ҏ��Ċ�I��6.��u�Ì4��Q×��Y������H��9mS���^���=Dŏ�y�<ILi⣺T3H�&!�L� y�W�ت�s��?h�A4�yk����Ve��6�����De�g���ȧ-�[��'����1ʙf�5��:s�1O�W���!`�1��(���n��08�^��F��y��H�xk�CMP��������yF��lg�
i�˵�[މ`�f�G^���}'�(�i+�÷嗴�qc����������L��p��Ͱ葂�m���X2�p���:Nv���s�ZU�3l�j����/�Hn���>��n0��A^�!?�
$�cN��*����ҭ���7wd�AdYC3�aWY�L�w�#��ǉEb�ȿg�4�!�A�����o�c��$�nr�I(��RGV����۠Ƌ6���<C��Qa��!��*ڔ�΂*ڶV�SMߴv/=��Qs��֜٥(��k�(�U5�B	Lw��2�ےs4���gZ���[k�H�; 7S����P�] F����bc���A�:����&�֚M4}�kix E�"b2��ed塧���B�iJR*m�J�lLǌ.�E0�z�Pw�]l(�)���a�V%�*���8����7���m��V75��+Þ��v�xu��r>��`��43NJ�f#�"�ȅ��j��ʒz��U�%�������I~O�kAV���A
{�߫?�K��K��Zr�о۔-G�O��`NǬ\�@"v^�t�p�r���Y3� ־Y�6'����\l�&��Y1%��"���sy��|��QF$5��P=ioKEM�K�2�^&���gI��E3�����U�dC}A\�1v��u���_x�Z�%�~я��"f=�\V`1Q�9����h!qKc��-����z��ݏCS�,��N�m�Q�Si˕g�����E�,�q��N	���>��cA��VV�r��'�,d�h�'�zjL6��h��h���-ީ߽k��ɏw3��7 ���Cvb�M�;���\iW�zF�x?��i����E��'Я6գ��}�R�h�"|hTO.�Z��؁�ȬW.���K�@U	�_�*��\�Êj�3��>2��2I�zZ�,t���+���@adW��%��;\�i���c���3R�9���q e�a�<O���n��:�������]&��֤7_�a�����Bդr���g:Md�%{�������d1�e�ݝ�X�-!C?�o����BE�W5-l����yzK�����Y �q�>�M�	ew�Ҿ�*��x���!�~{����l��"I>����q^�l�Un[~��}7��;��r�
CBzXX���`�2���ʊlNX��i3�J��S�:�ᖞ���dS��D��c�6Z�&*���*�"� ��D�S{�ȳ�������j�����X>��Z��s	Pw�_��,H]�����)�^��t��|:��VR⦰~����7��|��"\w���f�up�~�!�,��yDB�M�Q9�Ơ���M@����L�����XQ�,;L'��-0_�;p,���-M��=~?�)�J�r�f��S�_*����19��Q�k�FO�B����{\3Am�Mnt�qHU�S-�B��|M���C.͘��=R=�f�����ݭ�C*�ek4K��ef��{����M |^�g����0u�}�"�0�	+t!5\@��&��c�L�cux7��k��1E��h���~i[���b�1��塮HwC�h\�m�pk�>j�o������h�qa������O�)�7$�@	R�m^�,We7t�s���7~���������N|^u_t!
��,�bO�����!Ǔ��{d��9"�yI}aAȅi�hZx��T�+�d��X��b�������9��9"s���m��x��mOO��*X�k�k{���h���on����1�F8ؕ��|�q��Ә��(�ԥ�5]�>G���4C�n��͂�����g Qձ����~�c�C,�돓��LkJ��AO�G ���-sb4�8��:�A�� ���P�s�@J���ב�#x:��{��I�<d����؆z�}����Ҥ��5���=���|�6��0�5zM��E_�)gn���������2��_���'!�L�������hLv'�p��Ba颂+ѭM�^��W��s�<T��g�A�
��݌��o6n���s�	g�R��'6���R�̈�w�) �Fe���~{/�X�?���l�����-�I@S�k�OF��	�����Et��!m���
��Ew�{��a[��o-���7�%}�V�]>���ץK# .tT�%�'U�£'���?�p�]%�ص��8��ߜG7{���G>�}�;�����R��� ���el��26q�j��j�BH6p}���r�$i��K�Zز��c�e����.q� �﯏�p��4N P �p��3�(�Hq��l-BX�#�EK���5��j�@0 ӳ�T�ߔ�I�kaz�ʛٜ�%M���	`�����m�:H��'��}�Q����iG[�R�.�B��J�Q���I^��e�1v'���ެ�Y>�%�vQ�Y������9�t���ƀ{Ɩ* ~`Xz�A^�Mc_�1��g�*�ʀڝ�qWDC�Fh�����0D����6L��EÖi�5Y�z�1��J���������(�s{��k��qh�����X�5�1+�����کv�}��4u��`�G�á�.���U�ƞ���
-;B�z�/��}��l;N7��Y�=��M�����p
!��2�gT��R>�%v��1Ĩ/aH�v�%���z��Ka��� ���gv~�\�~���L�^.*i�l��q�o27lb��'F,�5+�� $K��j����H�_XT��"2T�EN��p�C�Fc�A?@a�����1(�s��?�v:�l�}|�W?����i���n��,Tp��߶(hN&�VJ`��.1R(k�#6�M�A�pd-���nA��+uO�93F�Q1啖��E�ͺ�̏�n�%Z����Q��?�	N��@
���jc1���[O����%�@0q�Y8QKF6�-V�PN��TtH��6�&�t @k���D�r�Y����I��y�o>��Hu�X����Vj���+cz���i�W�#!�����A�����:��`wK�o]7��KN�^P�!�-�OH�����/�cD7L���s���M[$˯b�Fn�������N�ۅ��$K]�C�B��4��J�Iߵ%��5�V6K5>Ɵqe7��R� "!�Qh��O�ƾǳ��Oie˟�����c4��pEP�zrR\�@�50��R�k/�Q�=� qI+�l�($�2C_`wo؅M�ݛǟJ���?� 6�$Kҡw3=��������{sĜ�8�m�э$Kj.�K�$e%��"����!Юng�|��:�YlJ]Gh�~��К�9F��`{@!i3�m!cW�V7u���J�}W�!K�.ٷ]��7��M}#���Yq� ���aP�\�wU/N�eo�#�g�h��e=� ����,&�Y;/��*$(�![qK�F���&j�-�,�C�jm�h��E#�T�{_�VJ���g3�\X��0ṻ^��Ŀ?�$E+�s���*�=�J˽���@f��O�Ȼ|I�8S�A��ءy��o�=F����,���H���=�d(=oC���~�\?��C�(��œ�����i�oqV�Is_x��69vsx���@M�@2����,��*ZSWu� �K�##Y�@NT�u��8���c/=�a=��E7�T}�<Y��ꕨ��z?!��{�*5��X���R� �|�c���=����:��@��k����0vǇř#lf�H��0,��Ovf4��~�NR�g-x�}��%uw�sX�����Sq��XRyϞ3���Z�h��*�35������D�bb�����B����82];/��42����p���T�ќ)짆$hܑq-#���t��qk6��[����#i��'2���G����a' ��$�8��Sn'�ԥ����nU�s�#�#�	O�����E$C��^�H��}k='4&]g� }	���&��\J,&����*D5��]�~[�#��#�h+^��=��J��~`��܌�l�s�Y�IU������	����kk.�����s�@��;��%,�%.�AA �u�%��"Nk������ w�m�oD��Y&)�ȝ�d���*�lı��7�KI:��8ի)#�ߐ�-GF�b���<N����ۄ�u�J���� �j�o�,�/:�����L�8���Ȥa����2�)� d�O�� �onf[����s2����9�q�=�)�]�Ă�O��j�,�YI4@~��+�@�T��rv�ͫ��E�%��
�LRҶ�����	��L�� �}��=Qԍt ��3F#)�O�����6�g	ɦ�ߠ�0��[sn�B����.�(g}
�Rn��ˀ=� .6�w��[d�ݳ_Yۍt��7_�>�X���ފ�	���K@^���Q��l���4�4qT�Y͕mH������>�{cI�j4�+4���3b��9<�+ԍp�����N,L����>hQ���ҬK�I���7x��V��$�ӂ��P=�hD�˲��%�C8{��<L"c\J,a�&DA����&j��K�EHx	�IyP7����j�~�;������y��������C��rFP�RXG��{/9�p4R�F���x�EK�mQ=^��H�I�C�}L*J�ǆ2vx;td����k����B	/�c��)�R����ʻ0��d���=+��rD����O���k�UA2��OA��
�V�=��_�ZxP�[8�|�bN��������9W"�Ci�c M�j��<��(Ԫ����� 1[�*�I�����_�p��>b�QD�2�!"�ߎk��C������z[�ڶ�{�@	F��#^N�)0�v� �X�v�5�{Qj��gG8#�Ȇ�LM1P%L��Ll�����㼹�N�δ_}rW�Sh��eł�Y�ywI��1ؒs5�hJ�%E�˧e�0��Jk��6j.6#�_�7�E�EDF�Ry��-�� ��"$3zy���9g۶�E���[����`��`??�i�ʩ{���f���
��|�4����"Q^=�e�qzwŭ�&�� ��=�צ��7	3W^��x��u%Q4Wd��VNV����Q�2�?;��V?�t=+:%���e���+^�x��eZl���坮:c��&��ؾ�O��{~�٣J�TIg} pt~�s�1���*��D��dY�Ҩ��Q�C�1�G�������*.˼R�٣xs��~1	�鉃X��/�m�,#��R�:X�����5�G������5�����{������j���#�
Wi�Ω�kSJ ��zP�#�����ln��a�b=NSrT��FޑZ��W�Ȃ��s�sW��Kv��(�m*.>�=Y�Z���o��j����Z+D0N�ְ0�x�R�b�L��7 �o�Q<��X�5[�d�3;��e�U-�=}e1c㦝@p�b���a3֮���L�i-��L�`�M�[�P������EvQ�N�����%�`�@��3���:T�ʽ�&��b�b�/ڬ�o�v�t���HR ��eN�a&�N���5�f˨�S̍؂w��OLއ}����Sb[�m]��~7��%�u�4������X��,��AD@�J
��Ӎs �&�֏��:���JJv�g�	�9�k��Ε���4�y%���iV�}��V�!݌��=�y E��b-B�?!I�,I�B�<��xC��͸�5���W��q:5�1�я��}����Z׈��ɶ˅#�/!0�U��%�t+�r�qAqz��xVꯚ����m�	O�$��*�B_�RE/�E7���
Ai��R���q�-#���Y^͙���-��x�_2�N���:C�Ng�o�V�C�AwN��5j���2\y�ɾ-�.�����v
{�8\�:K��"Ѭ���<�ej�L�j�>������bT��Ʌ�1������h����I�}'J޾��S�$(����Y�Ƌ��ug�|�B��*�M����
�}A~�}y�p���a͙�X�D]��@�n�-f,�PQ����i?��ئ��o�8̑*90�k�iчUN�aŽ�ڔ�����>U�vۤ�����;�ri	�o2v���վ+�y�n�._��������� A� �Q�[Z�B�a�?��."q�4E)/y�A�B���<VG��wx�
seM!��Ʉ��[���	��:CR[kC8��0!��+�D�I5)b���Z>]�*�N��_�v����� ������7Z���Ƴ:�t���H	�HpsIMX|���䐒����F�1%µ=ڭ�svp�(�j��$7�p튶�z{R+$狹�uп��2,V�DǊ��R�ݼ8�&>�����e�/���	��n�ς87�:��d}����+f�� ��c�� �`����OA5���t<՟�����z��'z�56*���I$�=��[ ��G^jD��� �f�=p�Py�Z�U�cY�"Y�B��`���XitR�W���E5�|�ʃ�j�vP�a�d�a�e�6�s{^��F<c��Ϧ�<G��l��v��U�|*� 7��Y/�0��)c"(-���`�ѵ���3|9��3�)9�a���O|$�7(Q=����db6���!ƌ�� �N��9��7�s�W�1K����}���+!l��6JӠ
2��'fgup<��!��~��S!A�3�b͠��Ψ�S�g!-?���ZYTq �a�,�8!��ip5j���:���		;�X�9�O��'��F��]+h}{�\�f5�f����P}��h�F5��+���!sײy?A��	\A��tڮa�w�Z[9ԀE�F�=����}�,��V�/��/n@�&��eֶ¦�ۅ\��7�B!>ͷ�$KR�wkQ�1�UoX��e�;C�����:	6T�����(��$L޾�"Ǭ�'C;qc	�F�a+�`=�g�ҧX�T�,�k���nZ���j�jd�<CP{��Q:�۝`�Mwޡd��� ���jq��u]��hO��<���跭��!��1R}3}^T��fԥ|(���Y�;j��%H�O���y�{�dV�3�ի�@%A��A����y���]Sd�� �~S �����>�R����p� @�ֱ%��2�P˕��s��C�D�	B�vn�)u�W(�e����>w٦~�1�#�X��&|1����.�/����w�g�xfix�Ek�����@��'�ky�65�f$.ˆ%�B�����wޱ7�g��*�RR`V�Js�7���(1��6R̒6s�_ֺ��/��?����P��|��(���+� �9�����u�s�N�'lԌ�"=���%����E��%�,LNj���&�*캙�2w�8%���	��kJ<�������YT�0���q5 4Y��9ZXi�Z,��J���C��N[u����@��.[���_��ܛ#�����t�>��r�< <�O���g�4�V��`4of�Ȓ�� �n7FP�F��������r�#+J��X�\IJ��|���Y�6u�f^��M��9�ϐ����h�rZ�s��Lc�cN����iB���E"ߊ���'�BA
�Ԓ��Ӗ�v��#w� �P�JT:�O�˗�-�a�2a���}_�l�S
��x)���m��A�d����,���5��n	2AF����� |~�k><���.Ժ�)�r'4�jƏ�n1�|R�>��*�*�b�<r�:0}V[�G̓\"V�=�0<^S��ȯ���.n��i��
(�f�9�Ο������������;t������ı�[M���R(О�pI�
�{�d	�G";Ѥ��F8�+f��q�z���T�fV�z�9`����ѭ�#�k�Q�>�^��Y/�܍	*0��i��������l�q�g��P����r�w�"�6z�候�����қ���%�U)�3�G�j�j�dL1u�`�'�.����b���z�%��K%�?��x��+���X�z,Fg����0��ֳ�ao��Al��<fI&��z�K�M=3�sU�G���!'½�U4rX880�����P��*2�J���w0F�R���.1� ���p N�"�%�7rZǹ���_�2�-�Z�
/�kV��nܷ-x�A�2�i��t�e4_31�V;m{�؍���y��	l.��_�,0bĕ}�Ӄ���3�8��c�OU��;|�g;�gG"Sy6�)��\��˯#J~	��)8�R��c�UL�w� ��
���oOmK�[��s"Mu
��/.��!=����+t}�M��-[""�O@h�p�F�Z�O�=�������"[�S���QI���O9�E�	j)l�D��Pj�M���ҫ�֍s����bLSj��{�5u�zO9�G��]�(���ِ�;�#�e�Xӗ�w�g6ʒ��0�zj�;2T����Y�C��#.���d&y��_�)�ĊR�"`p�/�rO��a'�aZ{V��7��z�Kw�l��ׇyqO�n��n}�~�I�*&�_J�͞u_m�?�7$�W�~��tr���J$�#q��͚=�����|d���ꜚ�N�C�Q����o~�����'5�$`	�f��G1U��t@Y�=�T�rh��ؠ��a��(�?|¬�U���@���x�W~�,Y�/�������ro+���8u�-b�mb�c��ލ>���~�9Y���ي[p�RW_��qͧ(���4�	��75bδ#~��oeaxߎ���6���ҸM��X��k0����������A;�����i�&�J��:�,WL=h��l���|7���?�7ԡ��&�
���M�#�v�4��V�{��<%��|�6�w@�Ow+z\<?�9�)�6����V`�?�����TA�5�mL��<N���CϠ�{T8n��l���A�f�h.,�
�Rl������`\{�Ͽ��}�;N{�Ζk��V\P.lr����F��M�cC�~rw�H��+�������oyԣ �1ʦ p6hOd��d���b�{ wS���E��;K��T	�~�^b��uO;�(+���I��!��yW�4���횮ՙdrZ���P�q}�����8��9���M,�Y���U�'Y�Kg��Z����K_s�ٌ��e�����9�iA��əmq��k�s�C!�X��'�']��j�ͿC���R�!��M0=�C����N��.�y���S������2JdQ��4���g�b)hO(��q���#%�u0e���t�oA��K�$)��.�O�(��~$nY�⮿��I�[ggbd���4G��΀vu��Յ|
��T}'���L/����f cw�3�;�'�{n�9m�Q~�H���#/�ۼ�]�\���m��#�9�i�gs|����S~��b̮a�>��)B����ߣ�B���_+�6j��i�r1:�;�N�ƪ��~GVB8��/rɀܛ��g�q������-�,>�M:�+7�R5g��$�P��2��co�-|H ��u���8��P�&�����Z��B��	�_Q�Ѵ~��\I��Ǒ��E���	8�+�w>p%�p"'I��$
���<_bt�mw�ن��é�2K�ʴ�i%=}|a��e��cX Y{9���_��c	O��.��{H_�lg!K�m�Q�D�.����W�r��D]�g�z6��
�'O���gD��d�_��
�����JP���59�{�)�q��TK+Yaz6;�k��aIf��N^�'��<r�N�+�DL/K^�Z�q�Kn�UmaR,�cWX`,봪m�]�r2���%���/P�QJ�ҷBVC��_3�~8���3����+����}	:na�z���cY��'�uT|�!B�-�k�V�t5_����FӘ��OZ�eQ? ��#��[m��#dI7]Z�&h���{Q�эf�m̓�۽�Tְ�Y��&Mi��i<M�z۵�V�\�&��i+K1�4�r��ş�:���$�`bjU�����b�ֻ��׌�֓%�kQm��uѫ-�}'��� ��̆S��:�Z^�)
��l����^]��� ��Mo�xv��	nQmv�]#ҽRdO��#�ys�u����G�wWT���s����4�T���o���q*�Y��q���H\�Am8kS�c�,��e0�:y4:`���3�b?�b䉖L8[����\3.)���(E���b��P�$".��yAí
)Y�I�N�Cl�26��B�d?�L͡nJ{<W0�r�sG�_�*'d��Mw�.�/���hb��7��S�Bs�C�(��KRj�"�;Jf�Z`��J���hg"�^mU��o=+Kݎ�<�u�
K^Y&ƃ���-T�T
݅��/&T���#��.2���D|�S�lvpB�_Zw��N���ߟ��D+K��VԽt�*q�q�]�`0@ύ���Џ��g��mƇ/�����PyE��j��n&�������u���\����sϽ�ZC/@� �Ц��N�ġ'��!����V�x����u�/�ڱj����Xd͕��L�
�nء�I���E&+;\�l/�
xƲ���LOc��e'N�v�~]�q�&^����Y#�'=re?���ygJ�~d�^f���ˣ_.�"��*��x2*�V�]ZR�M��2�tH��L3l�uV�l�Ug{l����ux���켷ߒ���ayA*N	g�D�s�A�WT.��\K\q52��@h-��"rJ5�۹�	�G�P� `Hv@���Y�LXi �5*]� [_<Y�~�Iq��q�7֩nP� ך�9�@'�,{D�g&���%l��B�H
��hK,�vf���w�S�KB��sNf�g����0�\a;j��j�[(zur�q��Ib6���Y�������b�$��|s׽��Y�dm�9���4��N���G��~�1�z�PQ�Hn�Xts���5�Ȧğ�n��Zd��/���;��U�i�`�*4zdOZ�T6�����k���N�� �*�ł<*����8>����%�f�q��z�SI�5�Vmy_d x~1�n���LK�"��j������%W�\�y%�-���JO�~�	�Sr��)���Њ/!�ւo�!E6O�-(�6�b��ɏ #EE<��v���Ջ�<e����e5�[zG������^���pi���u0(pn>f5�f���k��uǧ�X��v�M]�s�����R��g
r��LO��P����f�N }t�#ήW���A� :L����pS$�vyg�򾧝��
���hn������i��n$�&���� �m�;\�d1��<C���t�iIsX��A��c���`6q�#ǼR�ˆ3��8zZ����_�����;�3�>8���E[&Hl�8�]�Oړ��)c#2��`���<H��n��� EB��B�(xX���2=�yC�dDu���̝��x:�i"�	\����G��M]�M�,�����,��a�S��`k#�X�}]��N�����@��+�q�z��$����b�yt$�����>z�O�!d^y�GQ�X�ޮhh��Z���b�VuDB
����t%�৔��6�9<�
��h>�u�68j�|i LO�qUՒ���݌��w�b*'�c��(lTiE�TY�����F�O,����`��	!�H�"\���T�*=.�ʌ�C�mk��޼XlF�[2O�� D�B��<S1������h��S.�	�lK�GR8�Wv�~���m��1�1al'ˤ�t��E���E"^�'�'��*�,��\�Z���^=�(r�B�CT��Rdʍ��w�@����RP�|�?���<!
���+�l#R�}�ζ�e{P/��=3�������I��O�����c)��s�Smc��&l�b9I��5�KAĞL�`+�SMz)��`O�W��O%'o���]1��L�6D'd�}oD�O�:��>�U���Ȍba��H �r�����f��#!�e����O;��b?{]ct�&|�s$-��!%F�\�M�D�S4<Iq�P{��Ǿj0(���	���*�� ��n����%����-wE+��q�#0-�ߔ�>�j{oWD�P�#bX�I|Ykb,�yƥ�h	<�����Dͱ~+���g��!�x<�,�G(@�Ж���#�;�����C����(�������8����T7��z����l�b-�:��΀Jڍ4X\	�e�lTu�/���K�����9���4},��C*���\��'z\��:���.�u ʺ��%��3rWZi`�<���B�����&&Mm_3��-aOH_�O E�x�Sҫ�^�2N�%�8l�� F�	s�O��'N#�[	�}��2���Zs=�J��Ӽ؆s!58�J�����Qxs��ش����c�tG	�-|I��ҫ����J��ҦJ>��3�y�P���F�8z�n�j~$dod"�í���b�?��B
?4/�)%�@*���\m@���A���8;�=�E���I�L��E�q���t��~ � b��_����#k�p�Cd�ש(��� ��=�6^�T���P��>�~��k�����p9�Ϯ�C�I��N�a��Y�)wh�̗�vp�������/ڟ�`�c�0�)�DWPCu�1��tZ/%��-Ѡ�Jљ"� { ����'�OÀ��!�"f����?�Lɥx�$	-��i<����q����׼�*�?,P;l86'�*h(w�So��}&��`f��`<��壹8���HE�w/5��������p`���GYkKM52�����b pC]Ƕ|�����'T,/Y�Zr���DʢU2^,K����!���IЙy��#�В���j�:��B�P���.���
��O,�ۖd i�s0�M�ͪU���$:=G�������>���_.ߧ��H�O�@�KmOn�^�|�>�0�G������y;%��&��-���A��(B$e�ˏΞ(�� ĥ�����_�axu�l��C�8��=�3YC��kw�.��8�y`8��T;@o)��[�k\�^br��G�%���5��y�GZ9���h'�Ŵ/�ܥ��8t�D��
m'F�[U��;�g��)����c��D��@tK��V��V��'��ir���Ȍg��Pl���G�q��u�SR�LA���.d�[�+�,=�B�;j��&4�}�<�Z�o�P�+>Q��Z*���.lP�D���raa���w�2��Q�+.��F�1�\ t��a�c'�ϕ����@����L �T���X�����'��=
�F��(#[0���!6Mu�, �b�d<].c�:#����-Bo��-$�N�`Pj3�V�$Qs{�@���z9��ٷ�T�ɭ݅�0����7g�2�p%σ��8�� H�z,��@[�B��A�	Q5�ߗu��r?�~E����q�Ϙ%�� ����E!�2��5J�)��&4��R������į`F4��}{	{����ԕW.����Y�I�ݶ���I��-��v�D���o/�(��q7�{p�P
�$iu��	�C�s�NXn�^.7�_^�a&�f����u
�Z(yb6W���ֈAҞ��|2�: ���X4��$���F��G2�h��Qg=0g�+�{�i �Y�(S{����,.�槰�����^��L���a�����K��9���3�k��n�
��G)`���H���?	b�Z�g�u&ϙsuE�R�9z��Y����\���W4�Ŵ� �	U�=]yʄ����+s�J��Ֆ��2t�aV�e���Ҥ��u�!�]���z_EW*��a7����^����"��+o��`���}����]P�vt[�B~�y5��ܵ%u Q�a���Sq��$�p�q�
�Z#{�m�����g�ӧ��@�5:�Ⱦ��Q(^1ߗ�� �xr�(�Z	�u)�G4��XR�W�����+���ӄ"�ͬC�X$o
�J��<L��*=�d�Re�<�b�TD�<D��~�^��(P��i�uvd�]X����*/��
��,s�7n�����k�|d�c+*���i ��m�����Z�+��1����}ʌ?6���-�E�[,�>�+̚j�*Xgo�����=��%�uF�4���d�g�7��5����ʖg�+<�x� ͒��Y%3���lqz��XB�X�����a�%��
���27���� ����55�0ھ��Y��08�b������ʭN�M�,ԣαno�q�a�=��|�����и�p�4I� ��#9����!��Yݘsb<�s�+;؊����9	qs�:���,"-Xp0l�T~4q�Z��n�B���N�����zD��QӺwY����RP���F�9L��p� �I����l��+�XM1��es�~�s�
oĎ9�H�C��$���B�M1x��Y��;�q4k��wE��[�E�?�o��=�+���0����KVJ��<���Cf�C���`��`��V���M�(���Wu}�����_2�!���c���/�P߽�#�p]�\��2��`���[>|�6����P��ȗ[�\Uo;�[�EQ�L�"[��qT�|���z�1�
�t�M��\�(�g�5zCnX�ga>9y&��B���)v*iy�ߎ��{��q���Jc��z�ph��gCM���m�5i���i�ۋ\v"��k����b�j�7��{���K���ދɔ+]�B��Q��h���&Mw��w���
���p>L�~���7���sf�Iǵg?Q�r2!7<ja�[k1Y���q G Y�IN��vꙐ�$���塽מ�IB����Y�|����	�1$vI.�֔��T�;��N�%��&�L~P,W"vـ{�#�Ȉ�<��4�A�e�d���c�[�D�������s[7�OP�f���S��(���.y��asssFe ���A۫(q�]aA5!n�u���/i;m�_�o7ː9�6$���U7c�
蟏W�҄��8,O��?��7XŦvV�FbG��4�!�`�9�z1>$
�r�ːB���k�Bў�5Ф3��5$�}M3�s��o)���b������嗏��.u.5���=s۔�$q���(�b���д�G�cU���&�'TU�U�E���BR��������5ϥ�, �{�i�fkR�
�q>����h�5����C�C�ܟy�*��`�A}?!��a�y}�ڱ ��믌��H 7޿ez�4E��Ϋ��YS#�
X�Ĕ�h�~qh���W�������I�X����JaIȂ�Q2	�s�Pa�>��U�2���C�X���vF%�G�i��[�H"�25.���n�dׄ��pMk:ߴ�F��V�����x{�4�@,���k��v�|_1f��� �P,�+_͡3msGC#el�:��щ���gK�A�� ��J9��(�-��7�C,y���K����)�_�E�R�9��;����)e#Ԩ�9m � �ao��η�˽ h���f��Vi貍��;1mj��SC(���Xt�IJ���T�C�3!8�3�e�]�f��,���wRʶ�4Q�Ek�Q�%ѵAoLw��T<�H���U��Ԧ�@�_�����m�2�1$+m�Fc�7�
.Q�KA+���V�v�S�T�IZ���|�Tr��|_"�q���N�u��N��/�#s���PV3��jkłx��P_s���'��77����#����j�R��y`;N ySG�5��2�kY�Y�'������X��/�srH�{�����x���[ak-m���mi�e��UO����(t��3[*��*��L#���:;Ų��a^-�W08�fZ6��]x�j�Ɣ�n]o�ډw�!G�����S��g�+�*6vi�[	��}ǈL��| ��ї��l��q?�}Yy��h�c.��uɅ��2�3�s`�.�|���6�5��jX#�Qeg�\��סzb��mх��C�<�_������O]�Xv �3g���yc��~��ũQL�%b�+�i�H��4�#{�m�I��1Wv���@��eTO��������'i]ս�
"����2vj�S��Q�Ŏ^t�Yn�K����B�u���X�kg	x�d!QILmcw���N�7f%�MVE�O�L��d�Zs�A¥�Dכg2GFE��=	̙� �!�G�S����\�����} ��`��4M-貜�ң��1�-U{�Q��{m*�-z.�1�5l1ϔ���s=ħ�©�[Cw���A��E�^���B�$f��'�z�P�]8�����BaEqt������k�S@�&��6�̮�k����v	��\Ymdo��"�����w<"��,Ӳҁ�C��>l%)�Z�iw�.�����G3�Y�G��tăy�)����`�t�����	}U��9�&�&�^�|W�2 ���ɮ��e�
��QPH�����V$��a��%���.�:����WE�^$�-�In�v���Ӫ�G5�F
��"�Ն�*_`ˋkyR���讉Rx���������>���Ld?��k�f���T�Z��Gd��:Y�AY�d{�U�-B���K�%�}�
0�j��be�q�1,��gm%��|vx�� �Xz}a��[`�(�	�NА=���V �ԝ?Z��Y�Z#��֝p5�9�P���sy��I��ʉ��^#*4���״e2�#��~����N�q���A�]%Q̄�����>�S<���J%iG���}�w{Ǿ����Q���8N6���P\��~_.g��a!+|I��K9��~̵̃n��y���p���1$Dl�;w?��̉��^�w�іt�V״7��i�e���e��l\���&ś�5�XL �E׫a4�@!�+6�Bsg�56�Ϋ��EJ!%�*�3��Rɹi]����;��%6̕�Oe^��� �!�F��1m�\5��f%�`��gԴ��ݯ�����&� ±�+a�"���>-���f-�Y�� q ���&&,"s�ek*Q�m�v�b��Аg.̩��*��"��롫2�K9T$譄O�!�N���c�'��b��n��׉�}ب���4B@G��B���@��kn�|nӸ�^R&$F�$:�����?wUun(}�T�	w�� }��_��y��J�L�ol���"ׯإHL�mۀx����g8���XտT �W	N�"���<(�k�%u�J�(��i��4��]��ߣ��2������Puq'�X�E��r�M���G��&iw;�7۵I�¬U7M��v�w��0�}U�����YbMa9GFmsJ��d�"!P�uR�X�j��@f��DCn;џ�W��!�[��%Lf�c�MG ��1F�NR �w{u�2��<K'����о3X3�J��֝�wJ�sKBA1��Aߍx����>�4�)x�'��rW�������S����ȓ6aW=w<�;G''�/��x�k{�>�j������헱�����Oj�h��}����1L</���i�`��N���,�j�U�c���E>c�t�aܥ��v}5��ç���F�.��c�)�f��7���x$`�4����H��z�>ε�-[	2YL�:�'��%�i��}�����]��5�l�
�V���H������V�c��93���r��|d ���z1�eun'l\�B>����"�]e�h��g��K��}2�Yj�ז_�6u�8<+�idb�oP����[�k��E�K�</����uK��6�B�A&8ÔQ!��=h�\�W=��2/ �<L8|�po�a1����#�K ��N9&�M7�>/V�3�x��k��&�)KTƘ����K��="L4����%s59�uC�Ym����bS��r�8�Ҧ��<`�]��p1��1f��eK(^��a-&f`��aWd; �^IG'�F6{.���W���gj�����jN��5y
]�Av����mM^ѐI 9��5�š��e�C;��!���]h�qdS�ͻA�1Zο�� ���\�Q�D���9!v�NH�<SB]�_�׸�.�Z}ɒ�,Cg$�u�׿_`(6 z\öDa4��5jX�Y�����b�dPA�Ma!�vQ�jo>��"��6��p}O=`A��ŒV��)�Y�A)6�Qy6L����{�pc�"�@�~:Ř�ț�V����v�A�"4T�=_`޳h�d/x�%Q=Ņ���Df��|a������>�c�4`g���|�[����b��f�{ug1�t����Jn�x�*�_2���?�"�NU3ѱx�U|�ɓA1B@�3������X�O�s��9��4L/�lQzDS����f��?z���2}�
���v��*RS�o)�:�Q��]��}�l|�;�*MD�՟I,�9�P���p~s��T(�*�����hn;��\¦c����D��E)�(cb?:$ ��v�}�s��$�x��2�&������^��6K��en�~�}�(#G��.����>S�B�\���xs4�G]#�=�]_0�P�P�H�/ȻYe�Y�Թ�T�H���z�rVJ�w;���;�ּG(�7�iɋ�Q=�|.Ѥ+Ԅ���]y=����A�mC���B=�i_���Ы�Yp��z��-)dV&����R�&���$�!u6��,<�a�.d��mF��8k����	�o�at��2_��i.�%���S~ژ���"��+��C'G���0(�0�=s+Nt#�GBjH)�����&�~٠�?jf�5���:IEB�m���X���e���mW��0�ɔ�lj+"����x��N?>z�h�u1|PMa�MÃ�;w.L�`oM�Zn�FѶ�hx��oN:W&H�TKH��57m\��������4�*�|keƣ�>m���,�xS��h���N�;������[=��`1}4���4��KY]'�jq8�S��ln0Ɵx��q�t�iUgA���Vh����>
�g��;��?*�̨N�[��;b���9}*c����:�gse��I]-M��<A8w�K�Y�3�S7xJ;�b&â{���1���q�Q^����V ve��4T��k��w]s�l.��*;���I�u�܃±�M��!�h�W� #[�-?~|K�G�p��&� �$*\ߨ�Ke'��f����;�*��0�7N�i4�!#hB�?�3sڱ!v�C���V�7x�
'�8>y��7���s�ۑ����A��X:�y�n~L��uV��A��m�xQ�2+w�{Q�B��łS��0�����uǍSQ}��O���PZ7�s���{f"�9;U���JTl����x$ruӔ`3�sX��iRlJ�Ɏi~(�]�5Oɪ�k&�K�o�au��c�s��9#cJva�����ݲ�d�Z��@|��nKȎB��f��E�D�7��1�S4�C���j��!��+įA���W��y�k?A�>Gͫ��~a(Mt����QƵ�����+=��.R_㧨3`���Z?�4�1V�U���ϓm�[�e�%����%
�Z�+��c�!��-�߲��A�n����}L�lڲ%���{�V�IJju�Z���������smA	�g��[Tn%1���F>x˕+�5P�8��=>����q��:B�̔������c�&O�BѢ�C�3J�T$��&k�����F@�ɟ^Qn�z�欷w`�?+$�9��
�
 ����]���=�w�jZA��-RXC�!�A��{3�wp�$��1�S��9��KbJˇ��4%��4��&��bW7z�E]7� �'�tň��Z"��c��`�*&v�f%�Յ����A�)2N����\��8�Xyn��6)y���˸Yk����{!�Gv��J�"�b�ў�
͐uuq|�' s����^N��*��	����B`r�Yo~(��hN(��eR�J�{��i�M[�Vx	�֧�!����������aVr R>6O�뢯���c����/�@%x�M�`��բ�O�¡��ґ�>haV��+ZS��]\2��`�^qWfS+��^��#�1&p[�@Tq��ϲ��w���x���X^SN��h��&���m�]����`����\��k���[���vo1��U����4�5��[0Zs҂z�*��-�h}��]����_���A���|��0��@^���M�'f��.���
��GX&O��C؋7���눐�>��W�=y�zy���&��G���al���&��TP��!Q�&3�3Dm�*�ݞ/R�vAmα��&\��HF� �*�K��!�>�D��H0@�%�E �`掴���3���2������F=8��?0|����i����L;���<eI:=?Kfxd/Č_��:��hN�2�!ldS;_�	��FYc��=���V!x�9:��.Ў�
�� 4�J4H;}d�$�4:F~�!���\�����4�c0�E��*��v%���ětr*cg�B&�h)=�5/?��f
�׽��W)�#�5�?�g����(�f2j���y���M]���Ns`����-�Y�)�(26�o�Y�9|��H~�PJ�#[\�`�sa�v̵�0�C�QXx �D �d և�]�����_	��B��#|k؇C��-E�$�Eǋ��=�������K�a%
��M�5u72&C���062����NN���;�D0Ρe�4֕���1ޠ@�}u�����R�x�_���ʛ�p~�$uz�{c[=0�}yE�e|�)�OT,�t2FMǼ����VOf_`� �[F��a��;��u���<���p�Ni �����o	Aɩ�HȨ�����	Q�ÁՍ]v�����;��r�I D���Phy�
�����R`�p��M��%�娢��̍���1�H��G�;~�u.��I����E�o�wP���v�ιPP(��3q"A?�Ŷ�t4�s�B&��_c�(� �p���f����	����u"J���C���G��@�V�z����a����04<�"���*�Bk���ۨ���W"�h�)�]0Ӗ��5a�&쁙B��� ;�_�0�C��_�伛�	}<����,��F״���#r�$r�3��~?���lD�}M��S0����P��3����{�Q��O|H�p�����PUR���XM���\.;��irC�'���sH ��_"��4�OM�v����[��q��g���ۖE�U���$����I�zV>�]x�֐��
bq�M���u��3�Vp�� �������h���nF�#m!6i�i��9$����6 ]����>��=lN5nL�����Eb�}斬A^Z�'����|\�v������'��>��}����	~���_�d{�8���x>��.qV '�#��_� ����9��@���II�uHM~e�X��8͂�!�UN�1Gi���:��?c7�Rr����3�Gr~s�y�Q	��xw��vI�Ȁ��xG��.��d�l��]��nVv}y��&����n_�֙��Z�H��ѕю:ݻ�(�x	��\m�k�^����������"j�H��Sz���V����7t�9co�,:���H�M�*0���e����xM�_�ݙ�%�d^H; �OK-g�e���k��pRݰ��I�t����݄Zn3��o`���F]��FA�j^���8�P�i����V�r�;ďr@�O�d{�4+����3P����E)�9]��I,��v����r3g.ݝ4��vi��S��ș=_����˨��Fۂ��;T�54O���V.	�Վ���S��:�� .r�5��D�1K�ݰr�0=���}D�Ư��)������Sҗ�s�quj�Ā���J=�Y�+����<Tk�v˅_U�o�l�Y��;�rcNp����I��l�v�SG2[O��ݘ�9�D���x+t����H~�Q�d�A�iw�Ʈ{����VԔ�9��V�����Ľ�>'��
���9\ �c�?toaOػPF
������Ф�d��mRD�[���l��QA	�v$������7Ò7}���и�A�L 4G�J�����d.��UG���u�?�
T��J�vmR���Ɔ�e�[!5@�+��EXWp!�B�7{�F�J��ju�&WgWRo�?��
l�|=�r�Yt�O����]���Йt���N�-;ei�w#]M/����o!f�yW�AQ�`��-��b���`�r��
���&ԝz4@C�C�n����6���Y���p�_��Sx�T�� O��slƈ��x�L���Ҷ�=�QI�(I�ք�g��6._.�e;<��X���`[�M��Y�{�`��Y�ؖ����Q�����L<<OT���Ff�9]�9m
yl�LV_VÃH��R/p�Z�2hשB)�s�u�6��4�!C�rV?{(7�-	?I��d&kmڻߔ�}�t[�|U�@�U��ϔB��р�B��Z��-��t��G'|��WS\ҵ�����ά��$L��,6Uc���1���ȁ���#�q��1��y�4��J��B.ؿ݂.�k����ј�����+�L^zE����B��p�g݇�, �'Pm��*�vhp����2�+�AA����y��A�Q5���UdR�,�I&(䷌��f��2LG�	ugx�fT���N~����a"�"��a?�Zc����5�q,�����>�I��>��6
�a6΀���t�1j��j	"H�&B� ���`	M(�(F��ϑL�n��b<�f+�u��2>1s6���^��_�YWH��ʖ3�{Q�[¿%�态��O�n�O���eΜׁLm�1�Y���L��q7����D�1�Y1�`�*^�.���1ڟ��@�p���o&�>�s@�
talB,04+O!Wz��v>�����ZcM�
Lh���C���e/���m�O
N޺�oȿ���ާL[�����SRee����"�!�9��8���'ی��#�'l����Ne�Qꘁ���S�Y��;�8 1K?R�p�y���=}�b������r#�SC��:�������E{�����IH_k
�[9L���n"���vvBC����㬽|�������������& A��̟?i�m�l��Z�kT+{#gm�/�▉g(֠@�x4�#u�FF'C�1�,�c�I<18��i=1,qu�o<D��3z^�p�pT�[��m��������7#�"oe(��t�?�!�2�d��s>>Nv��o�ਰ,*���'"G2�X[?��b�ū�7^���69[���ۣai�<k'�3e������I��A�}�C+$�77X룠�x�5lX�����^�6���
�� p��'w�����v�&E�^�<0���$���{��N���Kk�16ST9������ql����Ep�W4�/��+<e�R�ge�k�&Q?�']���0��O�tXc�\֞���+����"�mP��ą�D�@. A�1�!Y��*BO���+?�;�����-K��v�� ��/��0��i]O��=����(h��X
<Q!������B�>�ƼR���]*U����?-�.F+Z���GsjW2�����]��e�$(܊��^�j�STL}Y���)_�T=2=��x��:�%KN@P�`�Ԍ�u�
��$��?*�����j؋�JdU���C��|�mGی�
���j��[��-b��7�w+�R��X�����֓T"�8������\�e�(B�=E�*�t�q��:��_�$v�ʒ�
E��V�#C;�ᤌ�˚d�u���Z�@��<3���"+�OU����k=$��![C|f��3���o5'ڟ&d�&렟�]�HaH�V�b�r�Ҡ�zn�9� ����\�{�Jԑ��m޵ю@xf����d��*��<[��~�^E��+::	6�RE�(���Hۻ��qh��Pt�!��z[����Ծ������Q�h'�cG��9�j{Z,�/:�ģ������'L@�	b����&ڜ}��	�0�qW � �%:'+���->�*�7<��A�WE�j?����e�p~3�O?��B��?n��,o�	���I�8Gh~�Nm�Kd��?mhM�({�V��,��0"���N��Rf�k;�O����p7YJ�v�e&[*�[�ľ�I�r#�~����nBۢ|b�)X���8 p���`��ߵڢ+�p4L9f}�S`\��iQ��{�6\'?2ռ�+�hc9�ǲ�AA=�LxT�r���/D�����QT)3��{����a��A2c�o�]�dV��Z�k�PQ(�l΅5x�#�g�іJ��nb߈���� ��$��o�9�U`v�;�R�bۑ�K`𷗴9���c�(Q�����˖�\;7����{p��Aݷi��?ެO�zW䶦�M�$��hf�7��MϤ
����戡����:M"1Y����`��DP�L�ȿ���v���6��h������f�A�+,)-�n�<�œ}ڴ���v�J�~��j~�׈N'��FU��N�"|�п�G|H�Ht䩄���K����8F�4�q�F7�{i�K:�U�$��!��s'�b9�:�(G�<�����:�\Z�L��`TFs$���aq��K�`���V��B���p/�� Dy|˨�����QFq����'�ΌE�p��s^��4�;�:������x����/w��5<��!�����N��H<@�Aﺴ�|�k�>A= |d�E�	���b>�Z�O)	J{Je� t�=*��<8+!����n��jrpM�j���#�&���p��yaӚT��ْ�Fq�����t�����D������+M*�}+�A?�&!/�F���d�(�+1�����;�������Xzۖ�=ϺF�,�H2�:��1>J�8-�_#���zRN���s� ]7IR�]�|��wѾ} ��
<�5���gV�����6/x��!��+��=��j�'!�	ooHcQӷ�1��s(�i%����w�p �u��Pޖ��b���2��H�uG"�_������UZ�ι3��FE&��M/�rӅU�]_����J(�>�?�G7%�
���v0����yw4�o�Z��v�?ߵV��jW���GÌ���A�J�(�T�{un�nG�pfv��]td���T�YL��%�+�[7y�ͥ�)�`}~0���~NTZ���X� �S������e��������=���1�t��Q'�/>�GЅMo�^��Cz�4�?��e�!���q�ٯ �B����ʹc�9:r��d@/���1u�C��x����̴Dp8�J��፠}�ĕx,�����">n�Mه[����@2�F�rv	jV������������A�d�QA���*�Vd�V�� � )&��i�`V�  2����NU�g��\�)��|n��rC�&x;f�B2��G�%[��ޱ���&�%d�L�v�{� y�ʲ���Y����{*	}�c���:�O6"�r^�I.U�@��I	S=�c���
f�:YZLAt��9�֚Jk�{�|��p��h�Ջ�W����rk���$ߣ	����^���uD�^�\�<��5GJ�q����0�.���/�7���VbVE�~��aLRۥQ��9E4p�<���XQ��9YU��i6+f�I��J�[�z�>�}�9-3d ��{��W����7���$(U��>�3C��R C�R�m��XG�l��[Ԃ��
w��w'�R���e[���e��<�h�B��%p9m峖�I��ՓmgS�i�T���[��\�@e���I��]��=���vf�*��$�P%�t���7�~���+�Џ�V��?ߒ!<�������N!�W�X�3�ؐ�r�OC5�������H/��P�MG��Q}�=�"M�+^ʄ�= �����|��;�	�(�4���F���B��P�6����a�lJ�n G�����׳5���]8�`�/?�a��=.e�*M�d��ـd����0E7?�����^����ඌ��4B��2"])���2�- �����u&|�<2^��i�I�4��ߒ2􄂓t��۫�1w��Cj��_`����[�4�iʍ+�g<�;>,rN�g�{�ih%I�8��ks�?�%��[��J���K�a�����>�أ�7��a���X�$':�qN�ڄZg;y���ި�3�����Tl ���K.\M~Hۨ�,'}��[�f�(�:H�˳�Kk[��ltl��G��NM|B^��ȗ@<j����֣�#���j-�Ļ�,�&7���"�-e8{��k"^?�<�巿7R�+���4Ĭ��A���F�0�vf�_^���m(�5Z$�#�]�r{�	��áC�ԝڂ���s�JX*��5�����pލ�W�#S��
^Ҭ�����<�Ul�l<)f����yN��{O9��y���F��jp���������d`+k'�Ǭ�(h�IG��C*,� �Rz1�h��6�)nw��dZ�4a��!=M3q
�w�������9���t{��7��y�ݹҁ�y�}�H�?���K���t��F@m�uOP��6�7����_�Z�Ũ�U���Z�����+��R��v����P�V���k�s� \pÝ���}�3F1�Czt�?u����E�#�s}�]h� Իwks�}��963C�����(�Lw��{����<�p@�'����J���&���X�	k��A(�)��nm@���W�����]*��ַ̈7��W����S��R�m���ed(Pr�Vkf�,Rqٮ-�Ր\���e�>�;G��F��������3�+Eihj��7E�*R�'CL
��G�"��]���m�;*�J�����{�<\r.ڋ]�q�����\�t[;LI*�9��+x/��=t�Aҙbr������av���9DV9P`Ux�<��Y�s|h�GKZ*A�I����Y�td�g�z~B�5��k"�Z��~��� -���C��k?d���; ^u�ȋ'��ë$�Cmo+����³E_�?���X�����Z��%�c�EF�]W����Ӵ1f*�%p.!��}���XD���m�+l#��V�:s?��1�V��rkNp/�QWT��ӀjV�vNq�a�	�Q�1
Jj��x��K�YLV��{��)��W� d%�.�|z%gS��%v�ډ_g� �]~�\�HZa:���/���G�$�;	e�R�3vQ�78mx�J��"��ȶs��þiw��nG�G��R(Vn�sG@MS��l]�*	ª`�����#���a��`}+�Ua�W1�QhFI<��.�A�V�F�X�4e|P���BSQC�<A�,��W���	���at5��5�d-���������??|@el��@��ScLq�m���R�E��H�_�hO<;/؝v�u6Ҽ��v�<�>���O
�ˡ6�[Q�>�SjL���<d��?��1�)��*.���?�
6q�J�w�,~�`�e�j4����/����fs[`���9$���4�W��0�Y	�ڙ�Y������UE\��[]V3�����Q@B䃅���G
ݳ�VO���d�" ��H��<�"X�1Ia�����'6����^��!+G-��R�$�b�e�0Z��'����0�i����BxlW��Nkt�2M��9o��BvJ��w�)��E�ǉc1��*��Z9]T��0��	�\�Ye��4�==�$�������K4���|2�:ɕ;��v|����U5((��j�Q$�u�����6���#>�I�&z;<�����tÀ\�X�ު/n��}E��0;S�rX<2��t�JOS��y�9Ry�\���2�*�/Y��.Wi�;(x���F��X�E����<Y�A���D?G~�A�r�	�$�S� #++zB���a�}�sԀ��W(7�c���p�3��$c��"f��	�������75)E���r�r�0C�"u[B��B:(���Ω?%)����ur�pr�Ѽ��ko�MU��<+T?
�s_=�źppx���_1�`��s4b�O|�T�b(F+!���V5Ư�[`��&n��V>�����B�Ȑ�.���c��kz�j��-��z#Q������$�u��<���5�ܴϟ3u�G��K�*��f�U:=Y�����O0�XYT�0S�_�/��&m���GM�kH�FH�8�g�E������A]����%��_Ԏ��i' ҫ���{���s_3|��Sn2�b������t�q��`�mg\*� ��*SF�#��e�O�:�ʑ	��?Aa��,::b�nG�%�G�=�i�ܨ�v݀�.~L�B�-�C,�{��^5;��C�y@ҿE��5z������]�_��c��(�+�;����l�0��9�M�^�Gj��q啢��`�{p��0���w���{9	%(@���z^�̿�U9�3��/_�Ϗpb��+8jk����W6RK=�{y�����l
~�����"ĂGw�����xb\eڒZz,T�(�u8�}s�+�� ��G󝭽�(����q��3WO��O� �" M�O�r/����B��q�#�3��#	G/,��d*#��ݹ���P�VMʟ�5���y%�>��{�̹� ��TB���m�7BG$*���Žx7�EG}<�p}6�佩��ߜ�����>���w8J�ܑ�F�=E�r93���L�g��%�Cn|�4�//ј����3.���Jc>ƌ�Wxi�5I�1�ǅq_3O�X;#[����`!�-u�(����>�I�	�c�ZNQ�@��?���ߵ��t�\�`;�� �k�g�i,2���<pb�';,4�S��IM��<Uд�bgjk���DMF;��+"����
�+ޒ��������">�+�(�kn�=[|3o��h��qB���F��C\48�ޅ��=�̭��_�
��ݚ%�O�g���Pƾ�����1}J�ͮ6�<9ܗ�և��'�����޽��?i�7���/˕��V�#��IWP$�~�w���.<8�q�5�+�R� �5)��z�0����aT�����G}�m�&�Wz��K���:�僁��(Y��S��mT�.lR"{ک�T$��c%�>PX�y�P!��"Wf5fs � R_�'[m��L	 ����d3-/?���ϡ�.������%(;>�]�Txm�k?D�1��\�2��4o����!J����|>�����R_+��ݳ����IT ��b�R۱��{�݆Tb�kHkB{
i�\O�0 ����|K�Y%��<q$]�3�z��������l���ϲ���q�\E����Np@#��Ѻ���Ts�)�m��)v<ڿkIA���+���`�X3�wkr���h�`����*`܉��h�(�Dƛ�� n;@��n#����9�i��ꕚH�a��&F�ޘ�iuR�f�s�w�2��@<y;���g��PA8������ҮR�&�oc�DQv�������Qfr�Q`vO�h|�Ќ!�߮Lu2���Pxê�����x��$d!��􁙞b�A����x���c��u���+P�Ll���<�q`�fT�~�l��ZW ���2<<6h�O�%&��3�i���K
�_k_\��A�"��6\�_�a��FK�Q�!e��N̡xUg���b��.:�n�A�Ͽg���i�6Hr��?�T]��Z�,�_ �l�ޢ���W *�7��;6����8���`h��px�s8饓�eX��Ò�q�z	6���d����x�K��xri�=5�g%a��g���c�_7�u��dڠ�5������=�#bo��n ��L]ِ��E����j��7�:�K$��ް/-J4$�3�B=�P܏5`i���^x��1$�o�E`?'���x�A2{��U�8:�09]��2R\��451E��d�M�2�8hM׭��Z�����`o����V:�?��h4yE���-�����U�
�йd%(kf��/��{f(���ft�Pu[d���ig�,.\���^��}'������k��+�SI_�(c���;�-:	�9|��U�l�e� �3��f�A'h�V`L8�պ�- [j<OP3/�k�Vq[^,�pk��	�{�"E�y���2�J�]��5���O�K�$�-R��B��+�}n�Bo�M�q�QB��g7�R\�V=�+��^��]][n�"�G�ժ�����ns����ك��I�uu�|A=��=������������Ά�.����-��s��[��46��&N4�������q��4<�fa|�x1����)Ni.E����-�O�����ʿMK��0����3>"�e�^D�Y��ˌ4�o �A>`�r��Nn�����e����L�6H�t�*A���E��Gc�<�EnA��	)0��*�x.u�|O MU�Pb��Q2�9��wR�Bu�1�˼�գp9���.�Jk8ӊ�r��^�f�I.j�a�(Iz�Q�d�)G ��!	r	-��&**/B�5��Zi �������2 n�IS%��B���y_����`R�:�X��X�7��cBPULo���l�������s����9��_1n�I7"����h�&=| 7�B-�q(:^U��i��`����"܈�9gw������]��[�^�v�HжKI�L��Q��+n��&��OG�k��j|�n)>	˴��%$�W�/�T���j>���74�aֶ��qHG�H��@�S,l E����b�j���)�Y��O޲��w�6��"�x9�|;~{%�L���".艹��Q�S��@�2g;PǱ06 ��m`��GԺ"4&������8�ö��%G}��	*ClZۏ�\̱��s��L�}��e�&TCy7kZ�9�B����A�+��o�	s֩��n�Y)󯝥&'���L*�>�f����}��o��p�輜[i��?rf��pA��xְ���=�;�<�z�lE⌥�L�b_rou��'�-Q����C���Yµ��DK��E�iݷ�=��R�%xaU`o��
]��w���<t?�e]�@��Jax|�l�dt�<.���+,4�Y͇� k��d��ҋ�%�-
��:����ZP�X*#^�,��3LFYԕ���"�^z�*��t����P�}��L��g4 8��vA�hp٭�ZR�ԝ���UhsL@6�<}q��r���#%Ȗ9�51p�p��u,�ϸ!�w
�M�$��	J�qV���mf�X3TiA*���|ƪ$��<G|"m�e�Ɫ�\����rB�|OἭb�y�m�4�XHy��ݬ-pG�I�m�f�*#�����Zv�0��
�gj�W�:��0Q?�ԅp�����E���%���VF�n�:g��e�X<4�N~�D�G�KD��@F��SшG9�'�x������q`�3�g�,c����*��\�_}��3z�p��f�P�56���>�N0���<����g�_>Z��$�W�L��j}=s7EmQ���d����g򢂃�}��*�꿁1�.�.1��s��x;Fl�:��uo��&���o�a����<~��l��fE玨�e�lӴ�G������i-f�|�/w-�u����|�B�~��!�b�zP�CsxX��4Z��ѵN�[X`�8�&���[���E�O�P=�2ׅ����5S�� �J�Z�����@�,9Y��z������R�h�`���jD'͆�0�Vq�{�EC��_J9���� /!V�*�|q�hS��酘�d��q�@<xV�6b�B�o������㵲��?�V��G�k�utT5���шƋ3\���И�����	�>V��ঊI�wޥ�_�{s��G��=j }@�3w�<��QA2\Q{1�

AQb�x�o�^bK�ݫ2�L\>�==@A�0�����B� %����q���Uˡs[l9���V�ϡH���A���rl/,IP�_e�ζ����aBШ�C��sc޵��9�ɆG�G�t%Dͭ��J:kf���t TdY��R]_���C�d:u|>�*F�wu\#�oS6^lկMde��D��r��/!\/0�,ޙk�t+���H�Qaگ�ϟ�o3���1���K3�V��|e��yli7��cY|D����0��4������N�i9<g�nK�LW�X�yo$�X�r�T���=!������^9�C�HU�����]���BW4�Z����˩ۄ7�Ej������x#U��eF��:�(�S3%���44(��{�:���!���3u><��C�'��|���[�@������1|nW0�H�S�<k�����5�f��=��ǭѮP�Y�Z�)���E4� YE-~E7 ;�aM\��3�{gg�^�`����W�������#2�p;&�� ��!m�B?�i=���3�¶r�»��(E+݊�T/z���q�X�j��~�_ww��ݫ<�����y��{;��弊(4=�
N��q�Z�˟@k����u�ࢨ���d��|�T�^S��%S�
Hhw�"�
���V��f���gr��/HZ����q�]��͉��e���Qꠥ��#��f�?t�ͷ��ӵ�Ѥ�,��?�^������a����h��R�]�v�e����6}���V����9a�(E2�~������x�
��u���&�7W��)�ʌ��O �D	�T�JG�������Ù�wD��Mt�ڦ���:X��II�]X�Ö��S�Z9�9�~�-��ά	j��O����Q��	�ōQ4Q6:ssi|��H�pO�ʽ�O�߹�i-7�˙={z���_k:��H-Y�t��ӌ\��"!Ϩ������#�`�	3���K�� ��$�cq!�zc&P+>.�dk���P@��^#v��5ϧ�V�q�$]O{�З��*^ȶr�,�e����~}�!ݬ`�5L])��쑎TO��%'�5���a+�|kzJ
�&ӹ#�-&&&���	��gl�f�Ev��L!�!o���1wJ��ĺ��pLt�q�<6��샮׌�^*=܉�������XR���#���ҳ��6u-�i�<!����zW�
O�D��?��.����q@�,Į����Y�u��/�J=�	xa�8���SЊ��=J,	�*�gƩ�5A�m_|f������K�»!U���_)��j���E v�������'��`k)��P���D���m(N�7բ�Ul�ű�ۈ(<5�*M�y=*�����[H�i N����G��"	�/�Ae1�!Rϔv�����0��x�H��r��"g<+����ݩ4�0�\����^13�߉��V���G���Y��2��M!K_��ɢ<�n�����ronR}��ހ���'ZVMc�ڎ�8����E��!�ch{c��=g�v�&�!�+�e(`qeԝ�;��>. [���&ޥ>������l9ПЯ�V���e4^�f`>֫�2Z�1��*��� O��cG٢=.L���
,���jW�?h02�EmI��l*�&�+�/���H��!X���xz������z���RR6׺����{ƣ�b�V]kֿ�X��/ׅ���l�FE�E΂��}�{9Kv�]:��q��z&�\�<T�)y�`�&;X�"�ߜ�����)z��2��w�	�����T }�����x9p�~)0�1sb#O5���F��L3b������~�p��؍�̹�}%�P�v��Q1�r�z�0��$��ӼO�TG�UY�7����k�e+�ջoqE\��}�@t�w$���=fA�w����Ldj�V���~�	�eA~��5b�Λ�X}��M9v�2O�1�+�W�5������V��@4m��n~O����vA���������d�2��=Ȥk��8i(^Yį�y����4S��PB�Cj���YlO�d=I����۞I����Gx��,��_�X3� %xB^���2��
/!>$l�d񹯟 ��B����W3O�l�[��ژ��9���I�v)~��co����G,*�������iۄ�o���H�S���f���v�l� #�d��М[Ǹ�o�U��;������� dŐ�}=��E�,!Mi
��9v��N���l�IÄ�U��'����E%�=Q�.�]�L���RQ�OƸК�A:������*o����Ϳ.�|Ϡ��N�M��̺I���V�@�n��d�^�L�,��y���2�n��5���ͦL���D�F�D����7��O6	��������=�N|�T���65��Uq��R=m�<�w)�� "�4���j=f���Ũ��6��߹�}	��7V7�zWp�w���2;�-O�g������r�n�)�
�w���Q�))ę�w04k+)L���~X�����L}"�~�e���^wd�+����|�	��ƅЫ��Z�N���e�7��(��k�mw�[���햧>:�{�t��I��KkYP��j�������Cv�v�N�C��̯Hz���%�"��1��!��b��\��/Oc�_c��q�tNc\\�s���8���ݠEh���
jr�H5a�;<Fڒ-Y�i��f�v�l{��ڍ�ʭ��P��%�a1���ZǠF��m��RMP�V�]Ѱ��QXb��x�C��
?�-��sb�o�Kt�����լ���g����������j�{t���|������X�> ����ֆ� ]w��qc��(��iC"��=?\�m-�$ہ�iV?K����K�X�y�������9C�f��P� �/��������Ha��Q$RW�MA8���H��4����Y����` ^��eCҊ�-�'�<����տ���`pb��+�'�'�P�B-W�b��t?U�d3�7n�|�9�����M�V F�pP�jV}ۢkW���Ǯ���X�B<�S�Z{5&� �k �Y�\�}A�Wc���#/TQ6��fU���'CiPnEs�^�������Z�`}�wA���:�Z�E,�f�	�)����Y� w���iX��1��՟��;s���~#2j�~p�����S.�sQ����е%�P��-�?P<�x�	���"��EJ	�h�oY�e}���O�e�n��sPWN��uw���J/��Z���
���f����m8k���8��������'��X��&�I���|�0J8���nǧ�����}�j���}ة�
��Ҍ�6-_T��R���D1���a,l(B3����<رBW�	yH)�t�D)�4�Ոh:m,���џO��n��:*��1aq6�+�S�"�Dg�/���YN2��oб=��z���l�̻�.���
�����9�26R����(�AAͶ���=�j�r�d��Y�`%f�>�V�i� ���^�Yߪ����0垕��#���է��եOZ�r� ��x:�u�����0���V3#@�j�^��� 4 W���r�!�rW ٺ��z� xIW��h"CY�������?jJ6v����
]\�d�>pֲ���'`ڱ�u�B*h,�\��2"Z� s�k1?|r���Fފq��h��U�*^:�3���+�3�^Zx@1���:^0&�IǇ���79�_׬��/�՗i{�[��g1;p�¹�%�~�ˠ��ݮ3ǿ��O�w��;<�
�nw �w�:��^���R����D��2K����Bv���^cD֌ ɛ���Y~�'n�|ar����|�^�ԛ��2�>	'�= m	� %޶0=!A�?�����.Z�W�t��q�<҇�J��~�X�c��#�.n_A�}o7
$���R�^��.��v��PFl5��'񻱯Q����+����ѧ�qV&O��_/���}=(Ӝ��#�����A�H�V���M�����>�l��/�� �1��q�R1����Y����ڄ�7*�b�:�ҡ�|rIu
¦���Æa���J|��f;|���Wi��{�7p�U���0��J#\�Ѓzbm��!����zQ j6� �0m���H*����,����MVQ��|"ѩ�8y��"�O�h��َn9�TF1����c��{B���j��K;sdk���*I1��KŜ��t*�����X6=�N��|��$�80��[=��Q �4*V1Ŭ�o��o��m����٢h䬟��0L����sޏi�����p%��9��ZBJ
�`K��gWi̦�^}��D��lH]\�kb��Z��FO�>)��.���Z�?�C�f�>��k���1���>x�$TW���$Uj:0����)d�|D�4�d��P}�5����������#k�T����¯ӑN�lj.�2k^O�mu�G�D�������q�0�-���0W(�"'�J<�䵾���|�>�5�y�Frj~���K�%j�c���Κ\���YйP�I��& R��rqz�R��d��8����O��dVH�[��gKW����|Cg+G�cp��P2�l.�-�E��ج]������Y撽�WWv��zU�E��9VT���j�^��N�0f��a��[�CT~��;��_k�s�Ҭ[����4V��w�l��.&T�v-�}JS�}�!�G�S��,�h.�y����V�A���R����m���#BX���H!�;lQl��Kp��	�՘�?����9�/u[��z0��Լ���Q�k����\�p�ZxEJ??,��s�t����_�c�)D��" ���.B5�J�V��JX�$��Gӆ���C`q^_��w�N?PTpk�?����E̻b}���.��`��?PU�f` b����!�wZ9��!ѿ������	���rđ�w����1%�X���`��Y�]���?�"1 ��W\>�k�Y;Z\A�"ѽ\$>�oZ:)���%A�6�G�W�娑�YN�g��n o�"�;$"Ι�r�����%��Uh.�r@��tD�qe��/ߘ<��6[��\ �����|�1U} �r�_���K����dUb�KQxZ['b��qb������c�?��lj!�C3UO[P�uMe�:pB����6�RN���	7�����%��1Ի���>�w�t��>��u #�E[�bƆ�GW�;l?��&�-��l���AE�g��	)硷\涩�|�Ħ�j/qvW�=N�b�|�Erc���Ԥ��mb]�_��s^V�?�����"/�#N�a�����V���_HvI�?b�l�S�ε�*��'�w��Ū��>^7Iߔq?��/��8d�Ҵ�lڒ�$�D�2Y瘿,���،���u�EӲҖ�2I�y����"�)A�$1��\HH�(tk$��P�',7W4��_! 8���2��ȟ~�Q ������Ջ��B/�)� I{ݤ4���i
l����а��5��)�������;�9���_����C�;��4�KT͗q�lJd��K`:;�Ul��3=�����h��q��ө�eP�.�9$��+�fN��3A��.��O�.e���uJ���U�}w�0+4��.�h:l���3?����SH'W����R�����744����Wd�Ej�݀�1=G���l����}�$Mf���:=�𖧐��Es�:�iWp�s�2�����Y�Q��6��y��m}O@��{ �r���4�.��4�fo���������,�����.A^ ���v;��p�}���)<�T4_S�ђdg\ڨ�n���\:�\���C�&�p�BأzHW�GW����� 
\�f2B�7C�J��������[)�8Sx�T�"S�(�k#�����'[5�E�@}H��(���ٷe��N/$�x�������r�"O�?�cܘ��L{��aK��* ���䎉S��Fa���18�a���eZ��4*k�b��,����)�ju�ˊ�5�Ipc0����%�S�)N���P_Ñi�1�T����?�a"�0`�U[���Ŭ��X���]qX�.r΃��G`�t�ݫ`$Imٰ�ǁ�M���-Dc]��:�wUk�� D���L�����+�Lu�߽�S�[G���6
F�̽����}�v�LFo�E��$�>�|��m�#LBP,�?H����1}���k�*�b~���0�^_�8�ݘMY��q.�l2̈�rъ� ����^UY�8���##V�-\�y
k.c��ӽ:�)̋-j�D��,�YY֑[���P�I8�Hx�7���<]�l����>������M�:�o�t�ā�%Ә�		�0�0.����	+;/�Sz�[w�4V��K��]���ǃ�a����?�Y%2'����� ޕ� |��#�C���|�S��)��\�>+�����x�k�+ ���ϙ�q����c�
�ܔx�z�uv9�{�=��Z�~% �M�=N����3�7�>$��K��x�2���M lf�esI�{��jp��\�ak����D�n~�?��3o�o��G��X�0!�H�Z���	Q����[��=T_���RPI�����6e]Ժg#�&|�l��5%�b45{x��A)7)[�֦��*8�����!�zMԟ��[����BՖ,介O`g������Qy�T�t��u7�q���S��$@f���D�v�;��f@���U�xl.�� �C��;`�C��!B��Gl��QHA���K��a�C6�א!�!Q�X}�p�!<�������:R����0v�ܧ�ьm�3�L�ϛgk4��:I��J�H�2������������ivk[�G/E����ݩ|Nv�������C1����'W�S�uNȪ�m��P�Jz7��W]��]��S��p���شRm'��B��0�c��M��U"�@�3{�lr�l�͔�8����;ᱪM�.��������0��Bǯ�:�Ɏe�@��
�r�T/�R��ߋ6P�z�H@,)$?�zOԩ�!R��{U�ƃ{�w&bs������o�#B�,0�iJ	�r-��}�Vq��G�2�C5n�͠��0�b�[TB�[Ǹ�\�,il�oCu����W �C��0�'c�K�	�5� �� �m8ZW+�aD�HR	8z8���uw<{��(�z=��\?���!�ŧ����	j��W�^q��c[.Ih)�̌6W�2�e|�m��k�T�څ�5����t��*���k�o��rI��a��ەU�I/�H���%���m��M�3��'\�ddV*�d,Q�Q��]V��t3^A���tՄ ��b<}�QH0�^Β]3�����e:�.ַ�[�O���8���+NY�s/��ȶ���+��S@!W��>�3�`�\�q���� �~�Mv��ㅛ��4��G)�i�.ȅ6O���PQ��봙�i��)�C�=!0��������u��«J'&�6�Y`Dbd��ء1(�!ڜ����Yh�� �	l ��l���{�Tnŀ��#Z�7�K�'Q_U/���C#�=���>��tS1fV��"����.�����&_n�C%^]P?�H���݄S,�� =���P��
�6`��|�*`DjV��;|�c����9P����SvE #���b@��k��_�B^yC���|"�� ������$�Ų��ލݷ&��S�1�`٠map��Y��\_�%�����YZ����!�.z�e����3��D�4�ԓ��`��r���ۜsCs+�X��Y�R��Ї>�&����V6�L�'����j�KV�czp�=���F5J�����Gg��$���M-�Lw)���o��z8G�n0��ߖ���.LS�(�d�'�I�Б���PQ�/��}��8�5@,l%��4�$ɜ�{���n�1v�U�T`����� +~������Lr����y!'nJ��D$2Ȩ )�ɳ<]�ʧ8��ʊѱ��6��C��rO���l���0Y߿��Q��N��y�d3ʙ�i�6?���W-��V��K#�v�tDL���v�����>2	�K|`hN�w�/�k}�nP�<y�=�v�������}���>��	Ca2�RB]�+��c�� 0�5n(�w�w��y^���h��"�#��0 >3�p��E���l�:s3:���.���9%Oi���a%�Cq�����[HNY<٥�@V�������8�ȡ��@�,�G*dG�	-\ �t�G���@fɚ����z"!��D��+#�3�A�5e�w_��^���1n7I��=�V~5h�77-�k�r�n,�c�_���%�#IZ#d����[27�m��3/A�G4x@G���g�<�9dn/���)a p\8�}iuZ0�@�rXD���j����}�O�/1���k�C���y�d��=�g�Ӣd[W�����3�7�_Z�G��Vehmk���zvn8�a�_����\V��B*-�Փ>�0B��-C��(���6�݊t3�Vr<�!�ϭ����UN���eR�|%�q�����n�qqU�h���rVU��6�ً�դZ�$��y��ST�� �T���>����hQ��k�v�Z$�`�k+��D��1�}&�8�tw}����;rQ��:&5�L�>��aJf	���Y�>���zy��2��Ƣ�!e����μ�Y��P+�6�3�Wy��V�
 �'	L	�é�p�&�#e�R���6g�!.YY�%��/L���O����T�eSIO(1�V
����5�7%��1�c���7/v;�I�:�֕�Hj���:/ưnL0�<(֦���{��&�i0���p�Y�,���4�_Eh������ā3IĐ�!��:HV�p��Mi�ם�/2����n����݊�7�'GN] t3@��
l�R�X�������`mm�@��I��PF:=�+��JE����|�Z����i�N��G�9�(��U!�\���Z/��V$�N���f�a�5o;xt�E�$!�5���\ Ր�0���$资�#h0�L�����%Ӗc��' �i�n�����ؐI���p�3K�ߧ��E������@2�3��|5��r�`��J�(�_`���>/�ʔ{Ϫ}�>2��{穅Ft�t��1E�BZ��=��& vtj'�����W*�A����*[�,������7��*���j�{��f  J����rB]@@7
���a6k���<-��wsver�����&�� ̠�G�Q?u�q�j�S�����x���A�ඣq�>Ǌj�8WC;�G��*2�Kls�U�\�k���ge�
@
�&��p3;a:�>YA��h�d|�����M�/T��I�~���c�V��ر*D_�q������nV㲖�y�.rX�;#�ԥ�9mt2��#f��fz'�3�OY�C9ڴkFP>J����`쾩x����M�&ͶL���$�@���Ƀ�ʗbz���cv��es���\��vI���`�{�zm��]���C��|�i�ޔ~�c���SW�}|�U���]��In�͋���ߒ��O��Z2�5�(�o�Qӟ뀃���ۓG�{��F�:��c��&[M|1�m7��UcPA��m��Al߽J�$�b�*@��X��O�V`Yٷ��CB���a ��5%����(d��<n��8��k�R�q���wt��� c�j�@S�j^�d���B�t�n��HP�r���W�yw`��b�z�h�굇8�7�+�'il�&d���k,%9�8lyW���v��TP��S�I��Tu[UܫXy��p*�Y�k_�#75��=G��X��=�;ݳ�0U��
���@?	�oK���B?��Zw-#�܃��a�^��_:
y�\d0�h����iF�gj���s��t�)�C���K!q>M���<�S���". �P����4iW166�`��$�z�	%� ��ԕGߢ�h}8A����i�]�ʗ��j�<ɶ�+h;m�A��߾ȝ5�R��kzW�j���o���F���8���4He�	��숻���&?=�P�ǚ���'V�imJ)Z�!j\a"eB��#P�[�<%:_�uI�q2u���*_�����b_E��L���L�J��c�O�u/}�<^�R$�s�RY�(Yn��&[o�(�� �K8.2���V�>���%hv���@�˻}��7�����IMca�$�����]���F���ceE��6i>�eJ>(�98�XI:U\���Z�0n���QnQ�{t@�#���!���2�?� �P���;�$͸��UR1�+�I/K��{���O�Ͻ���<l�".bY�q�Z�}<?ٱ��Gy*)G��j��i��X(�hPz��n�ja�����#�����iO��8��O�L�g����i#��0��5�QC���̻r/J�>�{cV�]|jzu��w��^���u����/�T'- ���d�$���q>`��9>���C��|�s����:x��v�N޿�i#&�B���:�dQ�������{D�x�e4��_�L#$�e�e�q�O�lO3���͹��ҩ'Y�ѝ��$�P{f����R�����ɰ3������'���]@�K ���O��T�m�J7¢���K��α�J��sJ�����4{�gYJ%b�[�:�����/d.��X-m	�l�w�
(a���`�\�ؠFO0���)U�qD��rE~��յԵ�29��'��<�=7Qb_�V@}��؍����<j����#BGL�"�\$sZ}�+}Q�>`d�at���^%�veK��Y˘�'��q�A����!���S�D%��(�� =�e��Ƃ�q����
����Q�9|*EkT�̚���XKk��ۯ4�Õ����0�[
����Ѐ��vfÛ7=�+JO���ci��e�Ƽޙ4[�wG��Ti��~O2��v��t}���cI�Fi��ەu�ʼۤI�A���c��s��!�4X3�v��}��/U�������8q��Y���_�����`��PA�"��5�~��P�[�}؁�\3ه�Q���w$�vF(��Q�|f�-�{�h�5N(��O�E���M��N����n�w�L�O�C�@�����cd89&ⓗ�G��wCV��pK���壗��"�PE% H�
T���R���S	�r���:>���ź�|.�e���TI0T�.�%)�3�#,�H�d���Q&��_����d��nqUQ�L��~�(��7lr0fR�y}aZ���$�����4�_r�b#�&|sR�F;��[Cfq���ncI
F��Y����d7�2�Fn����n���#4M�Ux��E��3��)U*G�&�>>{�X:��Y�җ#���F���t�E�E�Xb������8�T�nZ��j^��<<�H��~9�#Ra� O��{)�~@d�2�p��1\}b��9f�|U*ԑ�W��-��/|��k�À�����ʞ�R8ވ2]O����.?=�]���  ˧�sX�O^g�2����]yF]6����	�����h)� ����s\j	`������ݣoU��Ѻ�+S�YX������4�O��(˳��D/�;Q9[�����kױ.pݿI��6<��R�?��7� ��}-����(n��%u
�E�I��Q�<'�:��=��3%	_��i1��z��\��b��n�|��73��B�ꗣ'{�s��e:�"�D�q\�`�-8��x��#x��v�V�8�!x٥���o����|QW�	��<��y^�2�o��X�v�K���ffAk�B�
�͢9Q��l���h�����$VaI�1���A1쨰3�u�_��Lܙ�+�ʟ u���XI^���^VR';k#J>��q=e�����]�2X珦M����ھ?N�@���+�2�8e�a8	[)Ǆ���C�W��@��E�m��w�\�B����3c��1�˗[-(�Vi�N���F��?ϖ��*(Ky'v���>�Z���<[P(��ʐ� s�6r��i�I�r��k+�ql�A
�BQX��]�)��n�$�W-�^��8��oԨ%�P�!���OWj�!R������Czg�[��/�.�}�6;]<��~j�S�����^_��H[S���H �&��Ө�xceQ7�!�I)N?��p�sֵg)m�A�Z[;��9Xp�G�(� �f�s�,�
�k5/�|"��C|z-W4��$�G����e�c'�>&��h����oHʙ��*�lPƿ�_�f펣��&a���P�/�����G8Ñb����dv��-��l'ޕ!x���j���c��n�φ��<�͐3]H�IZ�5���SP�V�<�c@�פR������IF3�Y�٩ě�3���~�k�Zt�L�������kXan����'�J�co�ʌ�����6;$��yGpJ��f��|����|r>Q��1Z�?���Tj�ȁ��4�N+��!�Guo���T��1M_׾���:ާڛ��,���y���Ͻڭ�Ƃ��Vb[����HǺ��ٓ���g��f��}��k�C:�E��q�"7�ΘaB����3�YU6H-4Q���S(�!U����-<���]�a[~JfD�+^_R�׏OWP/���Q�3��v��+`�����V�F�<��U�nx-Ŀmv�ҫ��$೏u�)`6U��1"���Ȟw��-�����ey4�h6�$���*�r���a�S�w/��5���)b����ٝ��bc���l�X�pa���wI�w���Ԍ�8=D���cu��h���+w��8����1�`{��vl%Wi��Z���!��q@�E��g���#w�U�㛛w���E}0\DTZ��n
��� ��rG��ϻki�W7���
��� 1�]+|9�=Qyr�/�ZP���~�Uk�R�0P�����R29�P����fhT�C�o�����&g���c�}J��+��8�� ���5�v9TA�����&��C^�{�#9F,�q�Vӓ��s���R��D�IQ*�&˯�����l#�c��[�A�ʴ]�ҏ��<6V�Mg2[e�x��d���v���&Ʊ�����YR�|�f�:5��Na+�ts:��ג|�Z��p�`9+�Od�W��{�I��b9t�fWg�ѳ���o��k�L�p��=T��D[�a3�J�q��b�Fq��)�GK}N�8e��}���$tۍ����;�*��r���
�$��\J���U�����m�R��K�
�����<@ˡ��#�Ȏ��4NVK�h{���Kf�
�$�E��k?��P����CtpQ�����:����O1W�f�Թػӊ��>��3x�ꢞ�R���Ix�ř?
-�����r���s��Lt���!�H�O�hM�e ������/� ��o"�(�ݍYC����R�v�&��bz,*��k��v�����j���e�ф�XQ
�;�
�oq��O������� w�8��5�/HrxQ͔��R"�Kdum9��	�������}�Gz�V��m�E�.5����-p��^	W�6���8�>�ii��S6���e-̆�{'��El=N��e!�V#C,� �ϟ�m�Z��7����S#GT��]�o��5^�oƹ���(��7M����}����?���kn����?_�m�2��q�l�v��{^���$k2[�����5$�Q�G�h�l����K��(����~���qAd~#[kH:;h�DxE��96$HM��%dBXߍ�T��3�1�z���`	2�B�!1�N����8(Z�~��Ƚj�Eu��^��km+��,bOO^Rk�)��9�J:�'V�u�O+5��J�|�,���.W�C�OB�_��-�Y1� ka���t���h����꺣�s���T-?Kv�m-oe?c��<��%��b��͛�j��ȭ�f�i�h,��Ϧ��~�b�- �w�h�~
|@�{���B��W���6�2؛�ߒ���3������@��*ݽ���/�e�dR���rP�ȁd��,3�����H�v%_�ۄI��礆&�J�gU!eu�\F7#�e霦\Bx��J�hJ�Rf����_v*]*-0��3�����d��t78M6�C#�l�ыYɓ :�Ӓ^�E�?���A@�b���P�F�2���â��PC���!�v�с�R�<�&[�b�KRݯ\��(o��T[W����ډc���%g�E�\���tK';�/a�筌��*Ҡ£Krƴ��잩����mr�lqy�ej�����}K�����c ���i2NUW�us>�jy��k͓�5j�x>��VV����K��=W��m�]���Ѐ���!��]��������Ow@.��1�Ci�A�1P^C�v@��ћ2��2�g�86�TQ}���Πep@�7��gG)MdT"芥� ���(4�XB��{���6s��I����}����0���d�J��%L�B�V�p�.��x�,%��3�Gk�����|�?T��G�/�㸅6v\ca!���I�P,9���H��� �?'>�#���+��P�*��D-�F6q�)j�v<��gP�yc��M���&~d��B,�gn��Ci���qEiW�����7c��w�j,���#��ʒL��6��G���,B�S2��`p���r8	��c��鈺���ľ����#*~X6p-�e|��>] MHl�?��;�_�r�ØC@�?�6~�3�~��SF���gs�a�
"�� @����_�F�:�l~�=����^;����4u�TdjHm����{�|0��n�֧��epANA���/Lv��ҫ�b���МOAt�����P/��O�LR�YC�����:�NHy7���1�?ڰ=>�U�t-?�;l��P��T�'�=�%@,���M����6W3�2�sθ��^��7���4@��������{��6�a�^���}����g��p���[��^I��F:F�6�z��;uk+<x^R�Gn�j��!7�0j���N9���;!ce �"����ء�\���������]���a�
<퓶oEIr?4�J��������v
);:�~{���ea?;���c��J�ȏ扥;��=�Φ�0�Q�H�`�^��HY=WDt��'X]x?>�Ěe�G�W�j.�����ƅ\ggV_1�)�n��|=���s �gDMn�H����/�ֱ��%q/�!b����.fP���9�I~ͼӭ�X?�k_W$�6sq��o�G^>:�)M�?��bC�� [Wҁn��h`.���}r{�KŒ=�kA�# -%�]a�x6Z�6+�}!
i����r�!x��P1'Ro��\�3�~Dߩ�>�oG(�D{t��6�8�؟���Ŀ���s�K��UYP��u1�M�@X�^dhd7B����΢���xY򜆦�����_.��!��n�o�5��c�6D�R��XK�����A�'�_@R���X��j�G�i��qm:qx�WUSqM!�A)&˾��T�!�(���@Ld�jKh��`67����a����ew�5��F�g(&�[��ɰ����8�y��N����67�aB�7B��ԗ:�����<}�M�`6O���O����G��@�0"�}��a���;����c�~s1��
�Oϩ:(�|��/��_�S�K�����Ԣ���P�g�<�5	�)T8A��2K�g����'Ui�{�>R��]��7\�	��W�\R����ǻ(�,��g ��.��sm�D4�O䉸�>j.G�v�F����sb�����<�[�1և�̃��k-���yʒ({}����x�#�4�e�u3��;�sq?����_:�$F>f$��x�1�3^����J�jm��U��\c�=rR�<
Ї��#�	�
SD��N~]�-y�����+�Mx��Z|s^ k�Bb��E��QuW�)�_�:a@4��J�J��Gm�N��3`;i��{!d��m����g���OG�>�@@k�cq�d���ƶ�S6dk�}B
#�p�1�~:6��`�y��Xy6��'G�D��U�^݆�`m�ӛ��t7�6&�գ�@�vH��$�ͺh��Sx���K@�DD�{�/N|��&��cCV�`�Y��Q�W�C��LI�O)�\SqS--J��As!+���U�َr���Ci��D��`�����_��ދ���6 K��q��v�"���6^H{B��d�F�����
��d�g�^�Q�Ǉ�mc �������H<t:�;g-�+��j,���;؊&�̬��n��p�L��d��вr2����c�h�bj����ֵZ�����X��Ӣ��,���ޜ�h�Q5�
�f>z�b��X�����T�,5����зeA�aaZ�h���L�g�ao7�~|��QCo�
�;9'����u��FT���'s�Z�Lj#�jve�1�����m�i`E�)������7�C��\�E��������6�g�C^)к�e`	�^΢�3���#��c�Ąu���s�?9�ď��iH��\��A!rb��6���ɽe)����?$��w堔�%�ώ����1���Q����3h�� 7�
�2���㫰�@}��,�dm�V)?ɾ����o���N,���(���f��dSI�oȽm�g���q{w���i^#t9 oYI��^�KZ��6�!��i���ڒ�6�,�gr�?��i�'z9�T��}h�a�gN
�g�s��[.�b�j�.>Q6�zc3����3�ܰ"���L�Ӥm&"9�.�ƿ�g/(ܔ�9#��czW�$<��0~b�f��׃o��@��{˺��v5�Tʽ3�р�'�@�!!-�doL�s^ۥ&�V�5�� � Ï�ws��q�kn�T��ռ���J���p�O�_4��h�F� ����+2�2�U���de�
�K�G[i屫(J�ڑq���'�I��kq�M�O&��� ���'�6q����{��;s��Z������` b��*�ɻ���*�,��ɰD����/�v����YZZ�C`�V�!��Z���쳖�c�,(�R=O]C��c���yR8���<�����_�=;�M�13��] !����Ay��K�����|ܢ/��/� ��U�� � خ.,��I:��r�2��~j#1}GmԖc�h��'s�ѳI-� �B+.E�9(�h#̣Q'#����$�<%�p���oGl�9��W�O2B�%�$������5]Bǩ`\�z	�{�����h���{��Q6*����xz����p�=qO�b���D��I`g7�=��{s<�8�qn�����i���0,Pc���;�p�����ݕ�9�Vhd$-5P��emO���т����Lgo��@ڢ`%X�e���A��6�m���C��<X$�b��:��	�PM�`;2#�9A		���y�$�Ф����e�̩�#>�r�!��Q�i5¤xA������'��58�9��;p�hj�]>�i��!ו|��m;#�H�X�ٌ�L7Z%"٫y�Z��֦	#!RǡlWݐʆe]�G3zE{/�mU�<���MI�����X'8Qz�lj��Z܃���$9��}7�Z�H`#e�dN]G���W�:�J��V�@����u�H�]v:���ڒ+����o�l���H�l�z�!L�G�f�p@'P�]C�M�S�=�:f��|��(�~���?v��Mˎn`@��/�	�/Ȼw�"���x�G
�[9e��]��tP�A���[4�.�W����^/Cܶڊ.�~��B���
��d�v\[��%��}��T�n�1K�ז�&�<M���@>7�y��*8�:$��L݌\�S�&$Dݶ�w`5۶��-�=�	4�i`��s��(��L���inp��L}���1���JŘEI	�:�dc�._=�2�\��͉�>}	�;խ�`��x����n8a��e|'�x�⯠�7$�l	N�~\P�Y� j=�з��e:�/q�_��g���sV��k��Vy�cv\���K',N�� �0<':aR�Q�k-K�V:�p&����ٔy Rgs��B���h��үK	&Jʔ�q>rA�w�"aHT�g٢�)P���~��� c}�f׌������Qz�E�Ah!��ڪ�jM[S�7:���6�d ��|pű�D�MR�&Œ��������0%09�v��	�j�۝���h&��榵h����_�ב������6j����FjbV��6��+NO����3ą��m�6@SD�T�vC�"5����͵�>"�	�+-3-qḊ_i�����]U1�o���*��6�na߮�
^-X��xiƕ�[/�5�:��;��ꖻrm/S��O����?Ǌ7}4
��\x2��n]Կ"J4$�,�/�`�a��C��F��ĺ��~vPN3S%_�^��� *
�f�
|�f�{�ꀕ��7J��������I���1�-��}�[�cqk蘋�O�Yc��[k�\æ�OA�k�/�f����lR�B���'-�����{���{3���-�dnS��i�,��M�@cG��
lzH>�e����9II�ȿ$�����t��IC�Gb�������[��`_'0l;B�� {��W)�ܻ<٣�>�H�j�rͩѲP�Yl���"U�e5��^�����5YR_�w������k���/(}��I=8�WkW��?x��]�~�"PsYuXU�}]P��M�\$3�(���W�X��kJ�U�&Ŝiz��ŐiG���Yb���'tO�+�5=���i#�5�[��W�ꈱ�a Y��?+�M�Tׄ����tZ,�`�8;-�'xne�O��э؆���Z���ԅTj�����`�2Bh�A�s^�m�����Ґ�D#�vij^��<�f��������d��?P�������D�9�?�܇v�!s��j�����!��%+4�6��G?qڛ�ܝ�4 �)'Np���׃A��9����aM���|���L� ,�"�3����V�P��s��ݦ�m&/\�ʩ��A�MC�[�4>�L]���5�D�����_��7����&��A)�P��3���ʔ�/�X� #�U�!��"����f0�a�曖i����m���T��=��9�'�<�7Y��Dz`;�{��jD��['e1��Y�7=4jr���Ip���b�I�Ay���䤘OC�?���%z���ZO�66([�D�b�J~��6���sեN�0�8y�y"S��JS_ĉ+q�Y�b�M�Ɍ�f0����0X]2��4s1�fS�ņt���װ��Z�+�h-o��'`�]ͫ�q/���<],5� �4u#Q"bD�U��q"��b�!��� z٦ްC�����eD�G�Uͼ��l;d��դ�BD3M�o���?�=�<��-}��J7���E|A߃�;�2r@�0�D���i�̈��J��.Jp\
h��>��2"�Nw"�S�Q(�{Iǈ�
~��2E�S	�A}��e(�ڙH�8�&x"�L����b�Π=J�Ϻ�)����s������Ϝ�9� ��@Pp3��h�ȃ���k+�b `l�r7<�	f��9��}$��RjL�1�Qj�ƀH������Ȭf�?�u��S�e��E)��Z�>1���8.�D��1�Z�Fs���)f3�«��� ��K�����f��yˊh@�3�B��1!�y/�"���}����k�=�ZF�p�Y���킗{U�c1�Y��$�v/�4�q�:6����@Um �������HDH_���xa_w����%!��bi:n@=���O��p��9"��XV��/`R�:�Dϕ�Ȫ��7���sW�I��=�O��^E��t�D��Hf3�؃I�1�y�;��$m,}=�#O}O���=�+�GWÙ��#���J��
� "���1�'ʿ{~�ͼ�F͡-(��_����Ķ��)�T���[���ojt��NL��z|�����
Η��6��X�H����2��	9�Cz@V�s�����KR݆"��3v3������5e�8���s�6�2��Wsus"z��Cw����'�)E*��v���e����%�3���2p	�=���&��9�^�;������x��{�۶���z��MV�4��y��;x����"�R��C��� ��i�h�ń=j�7�c�RX
eJ�5�kY�ߤ:(����|��e�B|�:��R�{q��H@-�t���VJ`����X�}6��n<C;n�if�ر�U���t��H��>�
��*(dJO!-����Y!�p?����X�|/�p�|�X��Qͱ����Fr|6
�(%D�����M�����fP�a���������5-������ǮF ��0�.V���i`ƅ~V�U��w1T���P2$S>ߩ;������f���:pF7P���vHv�k�H�<����MРRP�ER9�����^�{�ל1�3cd����W$>�A�o�ة���JM�����������	f>�iM\4N�
�Z<*�I���$t� ���{�᎘�ܭ�'�c��|����lw�G���b;�t����c����i���1�DD����;�!�����xӖI�$3�+V({�gܓ�}{a�Q׷�1FL�$��qs��z�$h5�Q�^;U�����;�L9`~�����q��[�si�@��m�X�X�R�nQy�U�cҖ�$2�rϏ�����5Mt�����i��{�N@�ѵ��Y<�N��Q�H���/)F�4N�p#O�l�_��b���u(�P2�_��o��ű}�&m�r���N55�ao�0|�{{�e�ޗH�.��B@l�k��Z�N�H6�Ys���@�&B��������Oy0y�W׏�K�p��ۗNփ�ڊ���Tlqc����%���m,Tw�T65f0�ݡ�N{A�h�h}���@�*�0�H��.��d�KfU�1؜R��[l�uqI��7r�mm��p�br=pڶ�$�}{��|�f�ͫ�d�0�u���ڰ+���X߁��l�ض��]��sS��������OL@��8k7�	�!�i�AlX�c���R�D�ĮsB5Ԩ���6��Tx�g���s��F$�YN_�7gf��>l�)�ݼ�"�M՟�
lzXT1xP�xjL�������I�1��k��b�;p��Ҭ���y�QO���v|Q!��2�[�/�,����K�n�P��zUQ"ON�b8����kΧ,@˞����i
-;qͱg�ُ��xU�WL�mI�ܡ�Io�|��7�ț�Ts�h�+:�9�1 W�,�˟����E��$�����S�[O��a}Z�C��l>cN�Ko�il�?�L�!B��]��{��g��q(�x����\�����;�EE��V	덼J�kڷ�˹N�8�����V,�����=v��8IB�oZ�oV��!M ��A�Jy�p� "��0���C��N.���7v�\�7f�#�����!��+����,��7n�r"hx�KB0���T���y.]�<�
S�e>��O�Z����M��F�x��!ɷ���i�Jp3m�v����j��sߗw:g���eQ$WEF���G g��-�*+)�V�R�����u��M�6�J7=
�1pu��I��d�}�-�׷	���)�
0���DI���/2��ʮz}�D鬆h�~.�zf�rk�͍�B�xI���	A�ʮr?�0�	������
-e4��佛�d�~
2��QYA�ұ3�48X �0�0u
���@��Nݣ��FK�P�����o�?�p8ے�~L^������K�P<��b�h̳�+mt��0��@��P�e�n:Aya�z`I@���.Ј̵���[��:oe�z���0��-"�����n_N�(�gq��0}D|��~n?���(�9��v}��$,���] FP�ڍmKo�+H�eԇ`�M�7��Zز}9��f�݇�Xz}|�70�������I|}Bᨛ�y���7��tq�n�i�> �!��~Ug�3ugIX3�ėf��x]��&�AqK�;p^?��
��N�;�oD�SW8�����UT]soS�����0}@j�fh&����y��Xy:���s��D�$���n[[���V��2+dO�w�W���֙'"c�c6䴡au�1��[�T�D�F�X��6�h5��~ߞ��$H�����H"��Ď���ܡ&?�D۬����0PnA��i��[�P\�ŗ�͘A���M5�y3��0����^����^��f�f?�u<�UL(�N=����$\�RXV1[	�Jw�����T�%�Ю8�TU�K�?���X�6��>f^#6�Ñ����`T&l/�bMramD1�ۉ�,?��')����V�p^�М�n������7{���xh ���� V��-���,�b�� &�U�H�t�7N	�xJ��T�'z�%�
)����xG;��D�N ��#W�di��A��|��}QPH��O]�ud1p�Ḯw2�y���= �W?+�oܱF�Or�?n��#w���k-|��s���h��7��o�6�Q����~r���}�2Σ$�DZR���-̧6�N�X]pМ�^���ڈ.H�jK���S�v[�y���?��2�;uR�;��F�Rz������xm��=;�<�'$?�鑐�I:R���Y*�Ƿ�OC�[ȵv���˟
�q�\�Ώf�7|~���:��ue��)�GB���<˷w�T��"��9!;-L�ɠv�22�R�����&������b�\5�g_�o����������O?n�Q�諔+��?�,R1 �%K��;P�0���k��%b��6��K�7�z�=��[������"˥p��ou��� ;�ҩ�u��[^څ���l7��+ș�5�j�=�w	�(wԟ�d��M�X�M���C˳Ky��l���lv�Q����X߰�gx��x����8��*L��B����V>x��L7��/{��U��縬�S]�M���h%����XB���}M&�'T?#��L5�p���tMZ:�zs��E2�EN='�K=NdZ˼�D!�n�]AR\
��R����+�	�����ʤN5���C	��PW��D%z�v����5��K'|��{s0$�Qm��Ђ����s�鵡����D�4{?ʯvԘF)�~�̖��o��ZR$�7��U�(�R�U
��FD|W��&M��o<u@K�S�=����󺫑R��#�.��b�7��?�t�S�"k���n2."!�K,WC�HQ�e���=�o�RA��P���@��G
i�}t��3us��|�	N�70����I�8�y���:�{�5m��T'r|b\t/ǌ���a	c��c���\$y��l�Kb���펛#{�XXS?Y�>��?5!�T�3�<ޥ�3j�5� A�OU7;�F��V� K0U�r�^�C�K��������R��(}ɰ�SyamE���5ojʪ�������I�Br��?�E<ֻ��}����nFλ��B��g
�v�!.ӲQ��9��Ԃ�%n���J/@u�@
�n)��l����v~m� }�~+3b�{�܈����]��Dr�[�Z8�w�x��J�V8Q1�R��p>���6��{o=��5�K��֢s����5(�%rh�Z���:��c�K'I/�mY�Q1���!MƱ�?*$���n�G���{���QŚCB�`uK�7p	�?[zF�+#�*�\�!Ϯf�����ω��vq`���Rxr���᭼�q(9P���Rij�r�J�H��Ax駘�Z�ZJK�<�VԍY!�C��f{�H�rV�%8�{6�&B,���ƃ���f?���&�!�³w��*��y ��
ɞ�6BVvV$���̧̐����	�$�B􍏛�,4&�P��1ϻ=o��w�y��p1��C��zI����VҺ��
��d��-+$�:�}�z�RUMU*?r�9��'�T��"#�ǌw�����x/��6v��:O�0��d���Ge��bKc	�{KE��{;3��5p:ߓ�G>�=��@��3g�"Ky��P� d�V��IO:�)̬u��`���P,�X�q.�{�fa�jbSpZ���BKp�X��[���?۳U�?��T'	�Ǒ"�����Ȯ�)#i�˧H�N���`�-��)��c{|Q=�A��u�ˌ�/�Q݋댓!%y&����N��ť��x��ۂw*Ù�A���.��Ů/G�w�ի �@����d�6�y�N)�>�p';cx�!�]`��$a���c#�ж[�n�T�/5@)a�*ȩȏ+	O�j���+/����E9��&i�����+��Z�,��#m,%�K�cX"�"@�f�����ao#-u�k������ra�h4!��]%!�U���~��K�l"qf�>�����<SZ),�dD������^Ea�W���=��jJ��)r��t�n:�S���y���y)��ê��ɯY��6�s�jic���r;f!);�G/�FY4��d�
֠Z+�-�����I�J-��� �����Ӑwq��������݅rb')���;��p���T�򕈙�'�7������1��Ͽa*���n��쐞��P+k�gK��#��0��мW�g'-�X�Dc&��# �,���i���qה��X�,��ۗ�H�%�|�dw�MiyiF�GU~E��m�uXv�y�y`0�@#��1.����[I���ћ���6gN�g*�ّB�SQ�=^�k��m�d��:����j��Wy8�LL�3iA��ɜ����j��õO7ie>�o��R<c���8'��\^�t]��i����0g��K��S��@�K�F������k���a�)�1n'�>*�J�Tj?�BI&1J8���*�Mw�_ͬ��X�����~j�����M��k,�&�b#�O
,lt[]� �Z4�짺���^�0M�G�%��3�7�s�m0�X{��aɀ�ud�������c1�~�U4+pa��G��5���YSa��s�b6n�!+���YyZ��Gp�(�3W%+/�FX D�QӁ�~O��K�!pP�IE��#t����_�G��*:�u j<�@+�seɼ��҇覇z2�*��;��MD�J?�O��V�ֆ���Ĕ��?[��K�n�_�h|��!��k��DL$I*Q�H��S��>=[K�8�
������~G?�&.C�k�.�W�ry��H3�(9I~���k����,�%�����	J��g�����Ù4CE�� :T߽ݖq4��CD�
�O%J�zʪ5�szr�]�����oH�S�u*�rf����5>Mz�7�K;�G��ϑ���5�bەY��Dt���LݢE��&2$ 䀎��l�	���ap�X"�ұ+[s9d�<x�P��?HQ���>0V����2�3�W�UYY�Xv�%��9��֠a`Ή�ļߙg�P�L2����Y�1Љ���jRݙ�(òߍ;�DW�]fg6 �RT2Ϭ-�K��u%�L���5{����:{��g�!wV������?�H�H�tj��mİnzX+����K:ѭ�n軩���i*sAe{��@��w��l�*�5�%��b�ό�)�����v��O�b:����X�.��a&�|��g�/E�G*�%���#>��r�zT�����Z���Q�kQS]�2��4p �k��@h��]Cl�C������4�&��^��=<ؽxR�_ސpX���{� _�z���3�8A<45���f|��<,����6��?�Ң��P!�M���1�ihF�v@B�~�ƨ��۾�q�u(9����.�q*�w�p6S�i��[�.�5UPd�@"���W}C����JO"�"M�%f�{��ζ�ɢ�eq6��,(:��ճ�R��.c��/ӍY\e�I�퉃�Fv�m���?Z�B��c1ܘ��y�J8u�=��a��[����WZ���9�S�tMrXD%�g�F-��FK�
4��G� %��O�Qi�l�l�����m,�,�x���F���%����9um(�5�'�ֵ8��b���H|�.�	�!���R���A���*8��!��O�I!��CV�m�����w���/��T��B����~�v�����	��:h�����չE V�cԷ�2�;�Ό��$�{r/W�t]�f���đ����x1\�	�&}����Ef��p�԰�e�uA�r���4�͞��0�����h�^�t�\���[�Ҿ�x�Q�����8n.<�l�2�˧�c;U?0�C����Zo$fS�����{�D��C�~@��ݮEKV3�Y�E�|�����=q>v�Vׅ���y�	b��.��)��E�e:�f���i�ƛ�lTP��D>����|���0�%�q����%d/���ҖP5xw��sBˤT`�f8^��=N�B���;x�m�i)�.6���UV��0P8)L���CL��8s�δ$��M�G���Wdo�Jr4dr��x:�q��3b��[�ᣉ���lc���xY_�2R���,�u� R�������h�
�  �j�%�J�RK�$`�Pp��H�i|#R�`��*��p���c����?}m�٬q+V�N�$CR�G�%�Ť�?���ui f���,4�j�ܟ������lP&(���Q����~�Ja�c{�޽~��&Ӛ�/��$u�9�˫��vA��� kS����p�?�3�OПG~ ~=��� � �,^�z��|�\��q��[J�>��`(S��#�Q�R
���M+���_�] ����Y�}���Z�/:�b5����0��hL���()��4*H<�S4�G�[�UɅ����s*���k�~֗�ǹS_i\�����C��kGKIY�L� έufSS񷒋F��y���Rt�jMA:(��i�Y�g��K��Om�K���_��_J���b�)��;��@s�×�U[���-��!�����P�Oo�/"u"z.��C������P6s�9	��QY&@�
�9���5w���۴(�}Ă��V�́�5�����pM!�����*	��,q��n0e�4�*v��\M�I??������`��l��.z�\�� p7�^�L�JeŋG��|�m���I(�c��?�h��>W����j/��nzy����/Ѳ.���S���'X��}<��B$��6봨�eb�����l��6�����[F��*���Y��臘�[e��˝��?{[�0� �#�Z!�թ�V �	���t@w%K���Y23*nv��z�������Ɠ,esR��?#)�}�&Bm@������sC��\�`NՓ������z��d>�U�]O{��9^	s=����m���?��;�¥�l��--�'��=�����E���$�``Z�~�솀A٫�K0ȥ'��[5N��^Uh���2,��Z]H���&���(��-� �����s����:��'N��ʜ'��]���� �%�Tqw��ɞ��E�%�Q�����F�] ��8������pH[z2�Xc��N:D2R_ƺR�i�S�ʾ�a����`߈���a M������|˺��)0cLI���|�E�|�#��i�i����m
��Ւ�[�п`���6u7; QLĨeהF�θ�a��Ho2M��Q&��%�*~e�*4^,��ĖZ#~���
z|��E|9"I��`�{X���yP`S=�#A�ncN2T�I���w�g�/�;`@@�^OԐ�Wnk������7�S�K@����+5K��!����o����3ez�ͪ\k�*�Nv^�QO�f/tP���nB����d�����1�2;�����o�=�Ә�.0�8�X�d�l�q _�\��;b�b��i"�|���eV�^�y};��6p�({��ht	�wi�� e�ͣ�@}'���D��]���5����roJ�tp@\>ُ���D�C;D7��`/�b��0F,���&� q�{4R��HA۟J\�
��lQ��_�˃�7ഺ�hV坯�I�If�s���Y��B��=$�/6�3b}6c?=�`ҙ�&�W���@ċ�0>{�*���%�_�Q&���S���j�jI����6�S	�\-�.v�!��&�$�-ș�"79��@RC��)�A�܃���F�
lfe��B�S*�o:"�|dFm��W!jI�9Ô]2���/�Ez�fD������Z����uk�����5�b"�45-���y=�a6�J���ArF��[��74�|,$�gݖ��xj�낪�e�����P^�1�2�f4~���'7��ݬWo���,[�������������c� �|'�$��:�w��nr��q���}� I*���~ļ���l��"�)��k��L�q�?����V>���.Bi_��0j-��Y�Z*��}G���=W�|!"��CW�E��݀'\��.�H��x\��eG$���
~�ђ�n�*p襵: Ӏv�����4�r�R�^jY����wP6Z���$����k���>﹫��.�����ٕ��>��K�׃K8�Hm��j��q�!n�o1Q�@1A���'4Z�2p�)��W��ݐ �Tx1�=��> JHG�*����3鰕��5�05Gvv��h8�
�}�jS[/�#y�д���k=�����OBW�xpF�rl6�����c���\��g5(q:݉��2�X��m�lI~�h�s֞U> �;��唓>B#����9��Y#�@c�v�=��g�}�^�/Q���m[�@�P��?�m�������ќ|qB�,QV:e� �H9@*ޖ���r��i�]���Bު��EK�K����[�
��v���|�Q`#��-�Lrplj������O���a�u�AO�nI1lW��{o8I�uRlFD(]g+��mc<B�j��T�È��%�Y:���%��'��D���X�[����*_P0�X}qbo���Ԏ���V
�y/��F�w���|�Ψ��k7�u֚	���9��Q�'��������Ϋ���_�,N�0]�Z~��S�?k-�{7j-[�ΜlLR6�����]��Vh6�x?�+��j�PW[���1���+�Ի�P�
�Xɞ��fP:�As}�.:FW�2:F�T�����*;�4&�Gޗ��Ы��Rm�֩r�	Ĺ�j_PL��{ԯ���?���I]U10�w^ YjPף)
�l5���`5-5��w�(�[����7�� O��DCD��������
�����Y�CM� K��w�s_o&.e��c
٣�{v�rwM����٩M7Rk��L�����&F�{�<Y��D�|\>���J6���i6  ll��Lh.֋����D����t_��\��-'\��L����qu�V��1��y��vWNDb��1'ѷH����Yhĳ�J�]���asX�9��{ ��_��| 1��i����E ^��.*�<��u��8"O��S�g��FgRX0eÃWLc龆�4S��xw|��J�W��J��.RP�>�:l�|��U���0|j�%����&��5�墟��V_�
WU�q]AA�����u�˰�����S˚���j��5s������E�H��v��|�|"�kW�����hӗ��]_1�ȫx�X�}Ģ3�jnJ�&\�9ab�"�L��6I�\�S�a �Og�j6�����3:���͍t7� Z���fJ����-���9���?`���35�/ĝ����}ݢ*����R����w���d�j^�7nSC=W�������x�l��7�:��+c|,!�t��c���|6 �[<@��=�N��
�������T-�	��h-;\��}O��ߋ����N�U@q���|̋D�\'�̀A�|.̱I��Jx�$��q*�J��z(�� .f|�{�ם�_�]٭��&Nչ49e�l*/������O?�IX��1HT[	Z3�R�Ρ�j͕X��^U�c�SHkL���i��v!��/z{����`*����]9���7;G*�ˈ���p��vV�*�'����G+_+��,�O�F�6��[y���1��DR �	��p6kYq0y�~ �#�����fA�Q��QC������!BdR��s��'���/y
�"
&Q�ZP�7�BdPJ�-nW�:V${/j���_��ޜ~��xK�����h�淾��}\7�c	��ͱ�w^�ӷ��:G_�S`�>�4?�C�4k`��9������P1@�S��pdK�ٻ�i�yH���u�827���-�h���^��ecZ
�>&x� %��̀�ENk�����ʣN���75�v
���M@S%��Aq���[�W��+250BP�Ux��!�����W�>��}������b�� hs-�Ě�$E:R���� Z��O����ibu0rAdD5U��=m�f����Y< �D<$���)�&���`ٴB�Q�)M�5~�ٍ	6��D�:0�L|!6,�䀾,X�m\�8\�Zj��/&:u�p�ձ��wbĻ�{�v���c[Q)������Sꚞ5�d�퓷gv�%�Ԗf�����LShڟ�YW����?%����1�)l	�8 ��뺟S��8�!��OZ���a������g)�T���Ey��7�GY�o��dS����m�Ov�#���s=�󿱡��0Āi�We��՚U�c`��D���9�٢BZ���~8�$"��-��i����r�]b�x�_��q���^p�a�����%��q8��:V���������<�.�4t0^U�"��%��S�NϚ"y�LS����V�{̆T�\�ft�K�=�T�o���pav���3��[VbF��4L%�Ca�S�r�3��4�[!F�a u�Q��ߵL���>>���9������qHAq=\A�Tm#�Ʀ�eQ'�5��4PB��B��ܝY"
7�\�����ĞI�5�F��~@Yhe?��	X�a,��l�D��<����-�-�����k#BB�W��x
�B��H���@R���3kжѴ]�ي�ޖ���{��}�5���o�S�A&�p�0�,�5^c�6�������h�p�+u��+j�t��$���B��cC�EqGy�>��L+��^HL���&��׺�_�$�d4���.o��D��u�Gф O��v�e��t��夅���Z=� %I|[бp�d9���8��N�/v'm��?<�(�Р���iL��7#�K�ǵFZR��V"�]t2�R���½k����'q7�
��ΏGV���! "��(��Eo����(��jDkeZC�P�5񇵻��\pƎ4%)�U�~��C8h��r�e[|^�ə%7��n2ڷ�t\���\Pa��kS<����uW��~8��p�u���������	��*�,]C�V]�O��u��s/[0x�Q����{��ӽ����<������n3m�~�  AU�ᬝi�b`�D�BƤd
��t�p���[��4^1�%ZiR@ǝeyf`�4ѻ,`%!(�%��C�b�����Y�5�-a��J��mۓg��~�=�7�I<����7�����y�Ͻ�(�j�ag��t���g^�*_a���Atr��������i��*����]��W���-<B�~�B�R�7��}z1ͅ��H�zi��g�M�X�4�W wkec@��ud���T�r�#x����,�)5O4ڇ2É^�n<��m�!"#��P0'�;�4�����
gMh��I#�>�N�w&�z,T�3�C9������q��jq�[�$į�)�^��%9	�5SB:K�c˕�{i�k�=�I���B��	=C�%��?�v���94�O}��t��X?�D>0�"=�T	c��+�w��CZ"�J�@&�6��GDB�����4�^��^���q�p���w /nҘ�%j\�C䢹D$#�Y�&e�����Y�����^�3���Әp��G�'��:y�)���坖��L�8�3�����d���`S�}m����L���))�^@=��)�~���셪bw�'@��R(O�C��X Vzb�3��d�}�2�:�2d�糂�z8�;�V��}�f�8l�⼎��vOIQ4��)"��;�)ʶ�����%�ĳm�0}�AHwA�vu5��2
���>M��6z���A�?�K�Nɒ6 �Ѳ_�<�+ӘS��FW_̠D?_�l�hl݇���g.;R3���%(�q��&��崛5�����ꅃ�rd������-�S:�;��PP/Q�*ïA�����=w��J��ێW�j<Y4��ϻ����>L�!�O�� ��P�RzW9�=pX���M� >O�SƼ\% �\;�����E�K^��2	Q*�v�Y�b�(SL�����s���sc64g6��m�:(�����`�-���r�)@n�㭊:6��c;�N��G�����XpfB�u_���L��@�"L�|f�:�o�C(������vX1����3#��)�j={��B�n��Zh��1�hWG.�0]Eu?l����*F{>lA�]��
>�O�`����(�r[ʁ�֫����A�1w ��<�ܵ#�D���:�ڄ��cZ�#��\����Tc��q�{��m|�%��<o���M�8g��Ea�Θd��N��N������zK�8�?��p��E�t����`(!�[ٞ�g ��hX�*yz�Yb+�~}['�eW8��P�O�o@��N�B5gbR�W��4����2��ޠ���۰��բ>��������n.���Y��z�}3�e��Ja?[3 %�vB�n���H�}����[���N�ivn_�Љ��Q�w�T;Y�sP�N�����Q
vp��r�ߒ%0�us!1	����B~�e��	��nW���t�/��1�Ř-z��=�?9!�g��/�!�2���QKaD���k7��Zb�@�[k3�N߀��DĲ8r�����-Ys�s[}�k�BneZ����qCPڣ�.�`�BVR�b�#��P�9y�H�3"Ä��SF���>���j�<��$��O,�*� sz`����㫸�W��(�g\��+��:�gG�����޾T��!�S�sب���& �� ����a�|����{� ZU�!ѱZ�����;����Cٞ&��P��/M���ŕ�I���F!��{K[G�����Z�Q~�m@�����ye#q���#�˵��\�d�:����?ѯ�,�?�7��Ȑ/Tf��8N���f�e|qx�% #+��w**��n<�M�pe4/�����Xn�c�Ų��͜yF ���T4~��(Y�_ƅ6y���
d:�?;ľ��0�2�B�Z���O�Y۸���_�b��U��"���Fs�V��ﹺ�k��ƕL�j��\���}>?o�xq��S 6�|o���|�:���
����RH�Wޅ��,ӫ"�Lc㖑��-ʢ�q�b�r*wҰtoc=<������A��Ne>D��3�	@���9ܨ6+	A`���ۅ�9���v�su�Y,L#X��J�1�Y�Zf~��c���j>��i�=�Z�~�C��A!n�N����`��鶕>LeH��K����qe�)�U�4-
��hߊ��p�Yߊ"#lD�-�L�4in���U�K���e���}܁\��#����`���4�S�C����kő�D�����Y)���V�vP��(��r�������(�����iwk��ܷPXD�k띕����]�����V�b]d�mӡu���o�;��h��K[�n)q����(��T�\}�n�0U%
�\�{�[E8<t�	���2��c�O��yw<¦I<� 3�Kq������*�w�����
�i>>�����%��s*�uE�d&�U�e:�;��"��nY5����(ۉf�8���pSS�
R+��;�����{�y��	�u�~�w�ꎡ�ޮack�����)��';lLX�*��63�+jr���}��{��t��w~F���Hf<,W7K�Ȟ����B�u�/�wfS3���HQ����Q8��f�0�c?�Z�����-�:�GFO��4=2jd(���A�QPtR쵛��?��(}
�l}�`	�X���̐p<��&4=�gjӐ��{����  u)���F��V��]7�0��.h���h���.�sn�@�K��Tþ�� ����m���/:�I���֫Wﺍ̍��P��u�����Ր����S����_Zt�*h�[��Wz��=��.=j~	��iS�<b�f8��N�Ye��x��;�
�����1���T-h+a9��ϛJ��{��F@'�}���9#6��
�R���߭q�t���+�#_��.s�ING��Ye3�G�o��j���[�3���ޮDr�0>��V�r91�� �:0�=n�J�Y��/�5A�I߾�~��»�$GV�j$js)N	¨%�)�`ס�q�V3Qh}4�[����uQD6�ǵ`�C�7�5�)Q0_���R��\Q��$��]W�b�b�m�7Oxf�����t�xȸ����p�5�m6����*Jg��¹1EVg4n���7r�ޯn3�̵
@6=��5#���@�a�!����2����  �XN����C���i��ڵ�2݌I�*A0;��]�D�Nk�3����wz9�C	���7���9T($��;�U<G�˒>�QH�|io)�8����M�7���Ix_��cKdy�7�Use�٤�}�v�*O�s��_ΐs�?���O��"
��RBRaW��0�r����p�<p��a��Kk
7ғ���q��h6�L��S���"�TlTƿg�w}N�$�$���`ǳ���{��xk����w$��`�t���[� �"Jgs�.@D�@N�w��>$�&���6��^j\ɋ�E�+�k�q5��9I��ʂK���/�O���(���� ��q}zs�'Xࢡآ2�Ŀ���fk�5,
�rd��C�`~�N��`8C�k��D������3��� �z�'{��V�i'!�Ib�.�z�g<�k��J@s�����c��[DJU�����m����`"�ޖ�>W��r�޵:|���.�C8����T��<^�^v����;�@�����]*�VɷNp=��^�w}��ɈN�~#��8$c��!OC����q���|�v�6T{֙//��ŀ��A��Z�K��i�AQ�������Լ�ΑJ-Y��\w����]�8V�A��onr|'��
��W$�X3>P�p���E)ҿ��V�A1��:8èsS��GN��6�H*�
��gx8�*�:��_���u�R�еX�$�5��VԚ�R��xV���N�3Ƒa!(���b��8���݉�U����:UO�g��`m��I� *��I�]�2��O�E��Z�(Ȩ�c����c�
�Kͽ�U�X��3����FE6����&){�N�k�Ӱ�?��-�1�N��'��pK.	U`��H*3��$u^Gj4�u:�D���&���Ʊ���SQ�z`U���c�AfbQ��� j�͔K�� )�.�v�F�L-��^��U�f/�Iv��kuJ���-u�l�����c�^���2x�:��?|�k�q�ok�\��u�д	��&NtС��6��� �`�W[�
<����$�s�躵gb�u(�u*\gK?-�os�iJP~�&7��s?�;V������F�!��m��c����|+Wa�p/���w�jv�m���H�a���w�C��]�i�Q���UbE-�8�k���B��ڤN)a��u��F��_M����A��j��{�j�0T�`Χ��j0��d�%#�kj4��̔ǩ�s��h��=vA�?]�%*�Y��D���t�����<�Bb�lu��Y���:Ǔ�_Pu�O7�~�f�Q�ꦏ���.�\�ߟ������X���~����z�h�\�,.���.U�ۤ�0�؎���60F�����ɩ�zN�y+�����鋦~�m:ue5���C�|p��<ؔ0���۱���{�_����x��������o���Q,&��Ua�Zѥ��]ߤdZ���r����!������_;;���Xgn^V�'�|$\��K�-��z��� Lk�%�\�%[��\������8� !]��7�T�]�39Z�)��@�/B��!��4����Xj��`�0$-Txe+/��/f�G�[���s~�]�c���9WYo��ֆO��{(T	>m�	9+ߺ:zˠ4>�Z]Na�r1S��e)�C���]#���./��%p�z��t�B.2ꅰ�3$w��<����DEDx��G��&>6��ڲ��y�h�(���b��߳3�	q57�D�T�%��2�PCM�O˗�_=4;��Ɏ��^�?�}�54�h��'�� 0b�\���+�ל��S�B�vze�0��A�c�O>�M��2�IP���]X��(�(��T��v��3���w�8%�P�D����LE�Ā�':VgN|����M�хL=D��XJ[u �vYs{���!�::LS8t����g|�.KŽ��\��Qwd�zY-��<U��@�+�b�K�:E����A�Z�U#�/�%"�G����1�q�s����(T,t�$���Z�}.
�y�M0'��Dcc�x�墸'F��MS��2�,>Y��,A��؝Mm��C�<� ig��V��fD Os���K�P�g�W���N[hn��
���8��ڷ��%��������`���]�D�����`�(Î#�	96���Fh�7� ZA��*Y(݅/$1޵�5i��T��[nB�72�P���v�T���r��c�V�鎱�"��x�j�DL���ՙ��T����ز�xj���ϟa7q���z�75U#�f���v9�{Q䵾�������-�û���� ���b��tz	�ǿHV������� 5][����r���W��:d���~��D4�qN�e4*f����0�y��q}�Sa�
j���"�zI�(�i�7�����ʬ�գP$��-�Z�8�<V�7�]X��"�Y�\zzɵ���o�V���M�퇤�����%|�-�AV�?�J}J!KwWhE?W�H���!�R��'�#s�I��������]��.T%f��q	�0= ���0Z��G:���9��?\������l�d�BT��Eܴd)�f�W3M��m#١Pvq��3�m�F[F������,ddDxu('h������B���d��H�Օ���]�c��.�W�K�;{�,�LV�J��S�˸�/y��߷��4��p\.�[��q�ʯ�E���e ��e��)�mʹ˞PX���tA$��p��Ӟ� w��FS��p�b�fl��|@S��eй$�_J3_��;r�k�����5L̅|���{=	0䟪~��2/���̬�����@nB`�C���;%�ƥ�0��{[?>���\Jǚ��p��ᡚu��:�~�c�6��C1W����`_HA�S�QѨ&��<�0:�rkR��Sx6gDL��ޢp��u�3�먳a~���k�����^�]~T3ZO�*�0�X��둠���I�]}��Y|7��v���DȆ�W-��1uC(�z'Mj �dA�'�.�H��)H݂���9fh$ў QAgF�c�2#P�AH��Ǹd��i�D��%�I�����U��Z�f$�D�K����Ȝ����q����"�c�m4̙	����jQ~>���Ӫh���eC��Oe�d��{،yh�m��vKp�5�����mIäVXfr�A��.�_\%$^�w���V{���j�>P[�15g�5��c73"��
�ǭ>ٙP��ק�Y�vH��Kx��>g&z5��=�8� ��~���G��̄���պ�l��؏���o�^��͹�1uC%h2�����d�;���H��W�L+|�k�� |,�:%�3���i����_��C��]x��e)�i��g�Pj����qO*�k��R+���t�}-\Ա7�.x#�@5{p��������T��ڽ~��)C��-Bc�1lh!)|�n�HYK_�ŉh���Z�Ti��>38���3gF��#��5�bXv���D���Ѫ��叧�qn�Qem,ߗX'���q�r�_)���C�b��|s��.�bL�Du��>�w��kZ$���֟<3x�P��+��7q�&ݴRʼF�h�Ș�Ve��p��!�/��s����B=P0'_}��M���3!9L�N����T׌��}�o;.�'�@$_$6�*�v�֔	�R�꬞�G���(jF�a�_��K��1`Fk৫�)�� �3i��'��9��E�ۂ\�S���Y��/c�E AT�ֵ�g�Ev#qB����`d �J��5�pD&�j�Q���sI� fwj\-�w���8����G��sͲ[��44��s٪x���i�q0Ռ�y�jZ�����I���Ȯ�}�ϴoE���U�����j��˰�Yxy�r![T��(5�~������b�/9^������[C����z��u<��$)�2&wt��M�a{e>��L��Y�E4ǃ��ֻ��"��ۇ�藅�$���x�j�i�2ʑ�uQ���6t;�p�RŶ��^��cy�dU5VΏ�`����փRk�s�1*��XḸ��\��0<5�������"�]�ꔳ?���/����P�,�_�juu�(��q�Wiw��ӹko�Ape.
�t	�PK�|���Q����b���k��r���D{���[��Zp\��L�:���^	N��H��q�B;�ׇ�EWڑW�ĩa�����*郀9@I���~I���G�P� w� �k\�mQ,ew[��;�)��i����p#���m���&��@]R�E1eViUV�
#�3��n����o@R[��S�n��j����.	0��ώ�9>�Dú�@<Z*(�Т����B���'�V�$N>VO�#�5#xw6�h� ���l�f�+�@���-�<�Ü��VSp�NH�f��T4��:�r�@���|i�g�9s�X��%ѳ���,��V��O���T�S�`�a|V�A���y��L�PH��z���	;X�$b��S4v�(),����_V�s��!Y��d�S��h���q��c����h��b��$C0��x���lD�re}��Τӛ*-?2���Rj3�����g�g���3n\�yrc	��Zŕ�s�o/UtP=����CK�b0*v�S̜?zP�h���.��ϸ�/R�y�[��� ��/D�m���Ozv��&��ѫI�h.��/��,��d��[&��Ѝ�Gs��2�&�w���[��/���v�[p�j|����S����0�[�AA�����K�t�w��Zb�7���~j�
���ʪ'WU��ަ��Ngx��LxB�7�	�}x��V��K������Ш��݌�m��P���KK�0�V���ZV�G%8�0佌�u-�&��L�7��1YG�l 
�Ȣ��A�~tv0?>+�>��N]_��7�"����������X�d�`[~���������ɒ��]�j�ON�c��k�n"YKQ,�r��=��b����ZN��::�b[Z�����ܽ��ц�0�@CTa��8���*�ۆw��|#��y�c�/���$,`���: �|��4����Xy�����a؎ ��ͷ��޷����e�E%��h�8E`n��l�\$o���^�G�-�E�;��첑���J�o�P����i��tV�t�0�
���B`j6���Dm�J!픿#1$ִV[E\�A��/�z^�
ځm?�	�i�����x�}Z��Sw��1��"f;Ә۽F�jY����>Ն
H��)�ehF�"[����N]���S6�G4���]��sލo�}-�TG�j��0X������g����t�><	�����6T����5�	�2�������BS'���d°!�5�?����[���'.ݠ��W����Y��7AU���%����\�1�V�C�e���T�g���
~�D��� �+���%i��c��{�Uf���$�6h�?m��jP�dy�}�k5I�Ӯa���C�:O3�n}��Q�� �<*TXU�5��ܜ�ur=ru�:X���J�&I�P���t'�}Z�g4��Y쨍#I�Ѯ�Ю��Ap"[�N1�	|��C~����Oxu���J�N�@�����>��}�:�I�+ܚ�wJ��m2��1�i�"��h���=T6I�w��6�X������M�b�$e08�.9K��� UHi��T0�>U=�_Lqy]�T`[g�SV�Q5�=.f����?�#��?�����ġ��k`\��|&εq�����	���kaO �l���D���ea��y��y���Q�X�B{I�?�)A��[Zb8��t�/�aOl��S���}�=lc�;o���ߑ�g"�=�dg�cې��dQ�C��7��S]J��hhFӨ��F)��[A�)�|l_��u�˕D���I�`�f��R-E]_���n�m/����bܛ���s�����8W��͹=j<m����nk����Qv� �E�w����.ʄ_d����)k�v^T�3��h3\�]��ȓ�&�����CA��"�d~%)>ؖw�0�� �+D2��ZSŋjF��'��|���M��pք��.#rI�S���~��e�BQQ� ��5|�o#fi�YLdqŻ��J{�u��v�ĥ��>`J'6ڶ�{� ����Di��Q��T��tF<�Fнx��)o���#�.�}u�d'�<p�@�15*�1��Yo�[m�N��.XRU�����BT�u�b�#[��z�(9��M<�w�Z�}�����Իn�TKl����M�
���I#�a�m�V��%��A��P鿾n��f�D_89�шi���H���z�E������@R����Hk�VG3[L�1Q��Yy)%<M�Rg0@��.)��i�eg�y6u,���%�=�l���[f���_��k�~�V<����<f ��S��������Q��W��dL�v�S�������$�)B� $���D)��~�L��r�@"�	>���ѻ����N�M���o��XaTn��~��@�
'�j�O��е�3H��G1mF���;3�`�*�)Y#�~����)0�9˦q��N�j��:s�?^�#�~���gwS'���1���8'��sB!�����~B�R�S��:l^�d�Z�2�(P�����K����;[:�6G���խ����`����^ƶ���x.��iUT ��ފ֘�%6BE�I9*���r�ߋR�s䅤?��^b���]a�jU*�Z��*�-H����P��t�V���(��P�R� 
ߍ�{���ARE��3��ӧ���<�bBW�p O����s�(��t�?�_�:��+Z�Im^�^�j�#!Wi隉�掅E�z:V0�r2'Zb%Z�'vzy�1d�>�o���V�4��v*ܸTKB\ƕ����!J����$M�U��TCy�s�>J�E�����UJ�X�B�S��|H�u����iU�_ �	�٣����|̽`�Z ˒�:q@;0l��+m���n�3�j葿̀Eǜƅ�:kYY<{2aޞ����F)���ڛ�7A���Q��{wk�8:d���[�0(�&�dIʱ��9@*Ѵ\!IJ�g���j�c�yC�[]��G�(/��C��TE���A���P'�z��s��vl�j�A���N�;A�q	 |�P/{��u���q�Ma[KKj/���XJ%�<Ӄ�����VZ��`zg�1�hL7y�g�I�ű>F��o������H� ��KEd#<������ց�:EN�����=�)�����_w`3�σ*^�0\�<��Qb�(آ��E�S�.:@��4�<���Lw��\��vxу8~8��1WF�]d��!�����V����`���������&�(��Up��Չ����Q�s�t��E�ѳ�7[���|�K�~�
���&G���	�#�z��Ĵ �j�DtY��8)��>�#�� �TӡU$�OMdt�$�f�`��;�	Ya2���Q�(]IS������@l(~��T%'�9�]�i�Y�`�oɜ��p|�BM7�HU�R�d^�s!��1���3o��E�����Ah���R��w@'=QYۆ�ޥs1t�����F��y��K�w_x��4ީ-˹��$�����;Ƀ��DT����()o��v�u�QO��J�L����@0��7����-i�Q��ʗ�N��,{ �|��iH��+�J�b�Dr� =5V�R�?�6I��?��e'��?d�b�W-LS,1ND�[��߀G�W�i��<�._u�j~e�c��L��p��y�S�,>d/�W���+s5����%�4K�]��r���F�U8�.�S�H���Wщ�oh�'r��j`���S�����Q����p��Q9RF�8�U��JOd�P�8U�\h:�;w��)�H@�z���,�Y���������߱�����ٶ�B��T%yҒl�6�=���'�c���̐�v�K^��_
�巇)`t���LhJ���ZT8��8'����r#�9%�;�'�-Eԫ� p[�Z�B��nP���V��a�Zc�X��4a�b�"hX�	u���!�^M:Q%"���#�s�-�X0��j�"Xn3���)*T���8֍\��g�%~�޳xM��h���148��Q�I��*�ZH�7�4��0�+��ٷӝ҅d+��ũT���{y� g,�S���.f{�6�[�p!O>�H�PL4ZJY�5~�./���ϝ�g��ֽ萿��@�@L^7;�A�����#�Yg�Ģ̋c3��V,3�0_�Т���p��e�� �X�U('����8��N���]�d�[�~=$�=��\*u��$�4���x0�B5�ɼWt�y�c~��:~�V��c�~E�YX���7�J#����8�WA�+sjr�D���]��C��%���Yϋ�z �%5�&����!�rD�R'���rR��*Z���˟��w�]�Cnu;�sa��������wt)U��4��ӋE.���������>_��`m�B����1/�=B�88=�k[1��3��n�:��}��1�p����Iі*0�%D&�PvU�C0_+W�=5�Ϝ���J���2�<i �N�U
�;�hI�,%ۡ���=�:<8�4���kS03h���P�
?��n�R��p�i`߽rx&���[adfv�U�aS;�S�J@�Ѻ^��)F1X�%�`0$O�(�*!� �[Ӣ3�q�4*]��G��U���ޒ�R#b��y��a�^�!W��"�;�?X�:z �F��!���!�c:\�1B����*c>�n�Hm�T��z���c:W����%��������f�v�Qh�b-G��y*���D����/��3���3j��7��[:晹�In--m��ŗ���:�L��	/�7���������)PW�8u2*q��dS�i��eX���s�h����w�����$l���i>z��ӑ>��ig��a8�4�M���fZ�m9F4]�i݂]��t�P�l ��1��ts��p����W_u��TDҰ[��J9�_|�{.�Gf��^A�^������g����eɘ!N�D��@B`J�|3Z	?��,W~z��1�oN��{08I��;��8�a�,op����\o8�9�yޓ�KQ�����9�����X�S�I8�:����3����y�p9��z�]�K�䭎/���Kۦ��7�n��!�`�wDc(W�)&��}&�CC�c����`7 
�O=�&���kƁ�vOv��װ�u���F�Uj�q�����P�D���I����ShG��4؍FÐ�w�mK�cci��}��1�v@�*������j���O�=�`N��M9���l�vpwM{�c`"[p�/r���m���v$�(�xpYO�����ɵ#Y�`	��-��y]\���`�f�$�f���8GaG}l�1!Pڹ�҈��f�i�W���o��#wʾwbRK����tn�u�)��?�@���3�d���hߣ�����m����"�2L[����3��I�ޔ�)=S�#"� }��J�Js�w��d8����m��	��V�U|�*]&��"X5u��)�F�Y%�D�q�\*N�O�#B1 @ط.�#�.��L�H�ye�Hc
܉Kc����Q"A��ԾA���.� ��i�3��8���Pb�^�b�5=���x��W�ܕ�^�kD�R�������#~���Z]�����?����s��y�JW�97!/P��0�i�p�hZ�i[�Ό�S6������WFă/`��O��߮��W2af�,�H	\ȵ�����-FB�v�iG����&U�j��$��/UmPՄ�_��V��T7l��d1%�L�V��{�f�p�iAB��l4��0�^�!��1k�0�ґ�Nɻ��K�6D�9#�{j?U8�e�����"��*�UNY�H��\�u5�/���� o�_@��X�O�aUÿ/݄�7^��r��O�v�� *2�C��c�9���H�8Z��og�eF��&0���M��\�U����7vez�z�\�,Ã�^�)��.۔�~߳G�^o�Fm~@�K������HL��#h�m$w�a�xTQ�B+�s=���P�V��־�� ��Q��Ut4z�e�-(�l�
߶:�>SR�]C�'�V�V�~{ɑ]=Y��H�Y�)6�%�3�3��Eb�x_8(�H`�*��~�'���Xg���xʱkwW`Z)���n>�_�A븊1-\���Ͳڤ�Eg�B�8�u�M�Ze�(F�0{�˹Xt4H�����"4��ȸ�*��05+B��Z�Gdʥ�U���h�`<�v|{���n�����&wst4�sM��f�w�,��z��	�����q�Ga��v�D^oK��=�ㅕ�Y�?D*���`��)��4�G��
�R��UK�#� 8쬱/��/���:�#>~��`��!���i.Q4x'\�0���x4ߗ:�>F(E�� =��5�����E:G$�b���J�hg���h��
�,T>%�@<�����{�61��%�X�Z��^�&130��X["[s����?��VPkm��ґw�Yat@���r�}���a-���b֨2�n�<:��,�
q�)���d�Lr�A�i3��]c���H�	j3^�{�Q��`ޫM��Gt��ȅK�]Ѯ��o�#�r'y!b�"YG3�zT��`���Q�*�q����@Wq9t4޼����	6����.?��C�y"��͕��b�+{E��/h(����B�_'C�yQ$�ϯ��5\�Vv�i��Mcd<��T:1z.s���#ƓeZe2lc�"���S�5��WZ�n��?�U�����l�Y���rj!Ϣh���$�,�g�+(�r�j4��+.Y��
�4����20�i�Q._��0ߟ��ϛ뛜���5��t��^�n�h'G�~��{=#t�4���Ykv5��
�b^	�$�]��1��@=�&��9Jd5
ܣ�a��@��l\i���ܕ�T�T.~��ecp����̾�3�r��Q}�a�6����KLӷg
����̮�9�r��}!�D�6����w�1���௉pW4=Ic]l�+M9�侄�lzh�y>��P�a��%M+2zߟKPk�;j�k���pܙ�FT��ߓ�ee��5��a���&��d'������Qh�a���鴮/�zH����C�r�Ċ����|��<�@Ʉ}�������+>�����:4����a6���{���W�H\�S��\����[ 2Wb�ԗ�y���}�Vgц��c��D�.��:�'T�ł�t9��7J�v���Z?y�(�k{�Ԇ�mG2"�B~A�G���4��޹�o8W|G���N:<9���oF�w���B+i	�M�ކ���K_��f�aꎇ���|�~)�w��@�)�v��ۺp��o^ /W��^a�n|�y���/*}w��5/������$�X���Mp��tJ�ۤze*]���e���ڦO��2���Ⱦx��n�L�]���ʰb肚�5���06�c�[��fq�c�Ya�W�c�6��6ut}��6������p��g}ԭ�|]�=��q�u���~0J��;Y�JBJ��%���[4A����*��1+GU ?_���D�XP��lܵ)� �Td�g|9J����+/�����TK��ϐ���C�����[ɜ�H�g��h��B!tu�ɨ�$>�QkGLW@��P$�R��&4��^��L�\�=�J+�)���t�vǸ}�s�n�8Fаη�S�s<,��pL�M�HQ����|�1U�
4DW�џ�dH��o�I���v����Z[��I3��U��>H�6��M�4|g�i�|�N�Lh\�鈴!�f^��ӉR�sL�����b���k��-�D�=0	� �6&�~m
���`�of,I曝.�e��&��l/�����5S2�k�!%nͼ3�\�x��jB�	���ƹE�}wAN$�q���Q}���S��~	��`����g��&8>�8�bt�3_�)D�������.�u��Uu� g�F�0�do��+���b F�|�1���):��`�(j��ʻ��mWWJ�r�v�r��<w���:��ߔ���+?��uiWt�������G�p�$�ܾ�''�f�Cb$���mx3����hӶ�o���w�ONtk�_�6�s�E���M��x�Q�� ����y���T��/������[;>����Ќr3��ů٪�8�3�9h�Z�w�opS�ARy�ڰ�&EJz߇p�W�/�:��~'&�J��H����}N��s�0O۝#�ZщR�^�Xw���-b���'�$���ʹ;�tNs�n�p��|�&"���lX��e	i��-S�����a���-��!��ٓ�K�O�o��t�ɢ�0]����S�&�|�-��6&��n[���aB� #�MwtZ)�I��n=�d�'*��i�	QC�x'
s��f�yl/��t���i�����&�4⺽��8��Yy�BF��7=w@s_?T����~�#�UP˞G����lǠN��t+��K�}����t
=ko��Խ�����ҥg����n�F�UK�q>��+�\D�R1$XFӖ��-�}�i�<S�����z�:��|\p?����o�C�g�fG!�Yh��?>&% �G�ᙤ^A=Q���oQ��k��z��O���U"tg^�����>l8te�bPԙ}�4��Zs=�^f�օtH�/�K~%��;z�.�M��Uʇ���"OG/��t�Wn�;�Ɉ�̘��˄Fhı�\��+'�T"�%t��D#���|or^��ArfA�6A�5`՝`��zOs��w,������n�.�Z��xg��l|1���s�)��ֱ��u	�JE�x�ek˄�W�����%�5��� ����V-�=�Eo��熰��L����E㈅ܡ� N��W��_Y�|h|H������f}1�-�Ə��k��g�UO���܀�!��$�CA�P?�X�R�z5�L�f��*J��cZ���ۋ���C|��\�/'R;��z�p�*0Y)�iy�I�Ǒ�/���4�(?ؿ�tk��|yx�N��:!p�38�WQ���KK���*��������VX���F��u.����F��H��]���/�p���xi]*�����$�Jл�����$��84\������lS}�u�� >��?`s�[���"�Q���_ʆ�e�f��.����C�c��^�;�����"� �G����Y�������w��#�J	 ����}���	]��6�d��6"Ĝ� ��ꫪ7� ���/ss�a��Сߺ1�"��( �a��K�y�x���n�e$��B�x�+*A����䚧�!{�^Ny>�Z[�
�H��q�G&v�*�P�� �1/Y�h�LJ�Q���{�Y<��ߝ(�.__�� q��7��>�9�4��$�<��Jr�U�D�t�tؿ�O�eڴ��|��|。e%Շ��W,L��*5L="t�}B��Y#T,�<9����)�x"'�@g�)��Gwǀ5�S��x�?�o�ЩH�Z4�ocw��r7���|��tqf^󤠹��{"�`nv��/���W	�eg����P��t�Ɛ'��9���ʊ��v��3;H,�h7/����	o�L�Вׄظ����,���c^W$=�Ta��M�������T�>�!��&��:�2k����r�=�I�b�{�<P��/ɦ��������.�>T|���5��P҅s[?�9����q�|-��� �q�a���c����yl��?[G��|��]m��JB�� �в����lo+��|K�[M���Y$h�5���"�]�P�4d�6��fCL���h@�s|��z��X�����
qSau�kR��
��/�t(oŔ�g:�����������I� d�9E�ď+:���yW�	��j�DDv���YT�D�����,�!VZ�hk�yZ3[�v���0q�:gf>KN���P��:"= �璩��w@�`ٹ����V�Z�Y؆Sp|r��OO�^�����/Ȅ�;�[���?-_���~�FSỦİ�8��z	P���$A�N^>ee)��02���^��|D�=tm�-rC�k���6����<F�,��lϱ�ہe�K��]�KX�z�e�#���HQ�D��}��y�5�G�>~_�R�,���E�Eb�,���<�F���ę(YZ��
za��(P]=����'�$ v��掫E�sJ�h�J�Z+�k5'm2��O��"f��'f�*miU�^�b�qpE����8 ��+ 1���T?��� ��
�*(a��/��^���"�/�%s#a���TJR�׬��:�6}���.�ߊ�Ch��9)��S�ݞ@7���r$W�$7;4��6u�����‮p�M^��L��0�#��P�Y�����u3���/]ҲR���Ƀ��$守�����6�5�4�����E��l��5,�v�f�iSt�e�*l�3�8���O���N6NA��c�W՞�_���iO�@B���U���F�{��Sm�Ҁ����/�\\l��l_�Ŗv�V�j����?�4�T�}�aQ� *{=��1 �j�E*��<��"�;�	��6�.
.L.��W,�)\���AX� �8��o6.���I�8m��*]��9��������>�@%VOY��RJOy�͂/���U����#͗?a{~��Ω�����`r�����;�Y�Z]M�c��&
�9�Ê���eK�	k.�k��KF���I�'���mn�Xs�$���с0}*�*Q�)�����������?�QBX8!L��nj��6X�Է�������<A�6���ڪ����+�0$� �Y�*׀����{��Fi�+�~/��gФ�v+��]�9�
��8
�H�~�=�4+A�aʂ���L߱�i0��*�f�jq�&Q@��(5��m��ґ��t)4�M�X�i�?���k�%����7DH�l� �Լ�.Ԍ�����Qa<�9�3��h#�_.5>�GD�8h���h8�

�5iO��B\J�O��W�Ch�Wnu� �����!&L�����ԏ��z���6a��b��u�7�� ��ƇxS�8����}������p�ff	eohwm��� b3��g��� ��Ո]�P�����"yo|�Z/0�^����&x�sM��hh����6��>zһ�{K�l�qY���@�o�l�K	U�v���E� �$�����I���,g6��J�G�&-��<�'���7�덏	R��
q��^��#<'����Q1� �=��2�0W�JV���;�֍c�ا��ϟ�>�x�e�(~�er
ݣ/�)��TҲkܴ���{C%1#�AWӭ�7�9
���`p��s��զbX3�h�f�޾ı��g�M�ҥk07�6ܢ:����p@^2"� �r��f��bp!����� �����D���~L���8i�hC3�"g���#m\,���:^�=h�ғ�]� j��e���%�T[��@�4�NY0�����7�X�A��?�nb�
��έk,��ve58��1�b�.A���h�p�""6�Bt	=H����Ğ�P��x�.�X�q�ѐO���4ݓٟ��?��*n`�<}�7�^������� F�"ײs�������@�9����kޱ�a��z��j�,.oii`جw���ҦO�����0p�����tzߎ��_�4�1z�嬫�mXb|D��҉��y�S߂��9���} �-C`S�:��p���9��Dք��Sy����k�t�,!A�?q��+6��n.�*�แt�)���pi�!K{[BG+?ʠm���$�f�tcR�\r뷼�M�"C5�wߙ����`o�H6Z��yIz?\g������7,����$�Y�%
TQ��-A����b-v��nMm�����4�����&D�*���F���Æ��E��(|N������}�3�2���|��S�O*6��y�*�qB�?R)>X���k��>�H�q~�(�aHT�"�Sk�BNs{j{�X7�da�p ���ڃ �m�בK�XG��FT�kx�t^�A������#�~��,t&�}�
�����jK�����`�����W�ҷ�/#0�6�§ڬ ����ȝ��u�����ߪ����V*����RH��	 �L ��(a*����F!��u�N�0����5��E4�B���ɭ�[VE�<x�rS�,��v�(BG���4��)%͹��"���V ��#��Dm��
�'{:_9E
�&�<ߜ��mP�0��Tף�՚��"������MY����V�	s"����P)�;P~�1�-r�җ��?�`���Q^�g��?]�ı�QؒD�'�;;�c�C��l&2rQ�
�Ŗ4�tu�b
���n2�F��n��~�j�y(Н����˄v��B������nZy.֭q)΄#��p��-���H@����߂I9�h�Uf�Z[�o%�%��B���1h�`%8"l�?����M�'�Ԑ��9 O'��ov0���'P�Vt�O��F^�>ϟ�>�2��9�~����:ר�J�W��F������|ʃWQ�(��$��{�[ߌ/�]�#���WmE���U�9��Q �j.��/#��`Pn�$l�+%��C���Zn��o3��aW�11 A,��A7 ���	ٙ�.0JD�a�3����۝���~q,�R}R~T䒁��hP�w6��l����FR�������*�Y�}8�f�g����=��8��u���C���39����"�:��9��:>���T�-��!��X-#�R2l��Lp5Һ���ԡ
���;�?�p�Q�[J��J���v�@�lG�y����{�T9��G��G>��h�o�e��:�1{)1/Կ���@r��Z�b����3��NG����ĨM�Sp����t'�H��IM�z���IA���U�|�6n���1��bJ2�u��1���?Ů4��K�0���}�L��F�vAM�,�V��.�B�a
�T�j��T��kğvr�`<�-��v�cg2���/������D�~�o.��p��|d��T��9mc ��9}]o�W|H���c���o	��裍�UW"��>���5�}��i/`_���U���ђ�Q�Q�?���R
@�Ӑ���v�ʂF�L�C���Z��a/��C�����\ɍm�Qr�'(ggBe��R�h)IN?'�O����7wgQZ̫
��7�Hl���c�ؚ��&���j��^���9�Ǳ���hi5��)"����S n{͠�sr���ڪ7X�6���p��f6�����Ba��7�@h�m� A���>�T�7���>��55�*��'�;?3S�ж��!{�d
`I���R�LͶ���}�q�(��~�B�g�-�0� ��mw��k ��;��ľ}��x0��*]:�A��*�W�U�l��ؤ��?&L��5��� �k�|�>O���Zc6a?�o�������P�pO���D���!�N��,//�@mARU�K����Bh
�������
�d>�U��/;_�y'ы���A6�e\�s]��6��~�����5U�)���9M��2�4��[I���,Y"�.���>�4�����(,��R��;}r��&��F��\�c<h����{!Z*��ò�an�U3k�yL�	�hm�������mE&a�tgVЛ\���L$�ے>�4h�'��������.�?�X��R1g�[�Q+ה��=���u¢a���0B����H��j{,<�/��ۇ�� ��jU�:�͵"!!2�IW�XϢO���������?�������?͠m[��f-���	2!�!$��#�ot���0�6<���%����H��%�W�g�D�[Ƞ�d�ϓ^�[�C��Ģ���r�q�s�LE���0�!�u����N���n�F��ǒ��~�T���QQ�9pE�O>}h�C�#tW�Ԗ~#�bL'�'����."���p�{���Fw���z8�&� ��9uwW��I�A�+��4�"1(	wJ6y���̄�C�R�����6|�y���Lv~<�%��o����	?��G)d�V��b��@��+�J�bV�tQ7@/]A.�@1���>�TkoPow�~i��`$��T�,���&S��_[q#1�T��﩮�,n�SWtd��D������1�ҁ5�RU7������Shm�����{C�-v�x>n'u(�h��b�1�W��9�Q���/���H�ks//D�3x�j|�� 둈}��.~l&�5:O��b(��i!r�O��D�%59��VwS�,F&<���=T�T/&���OR�8Z0��kG�?��N���0$�}��h�{�UE �"t���~$��	��|�-8�]�<} ��v{+� b���Ze�]�����<��;�*(�:��������v�Wc�q�Y]J_�Yb��bya���)��h��f�{�������M�
'w��@�U
r��\~8�kH���N �j��M{͐��J5��\�0�*N,k|���)d�n�\;`���P����Y��:DƁ�Ʈ7xKi�=�Y-��-�A�����0b���j�@�����Ց=�2�[���&����؈��*Ջkĳ���``� =��R�T8�}|�B�ڰj�j��:���¢�נ ً�`|�h�ZG�{P�l_"�����!�
��څ$���ê�)/����`�]QW�?�ZH'(�C�}<A��{�}���Ȼ w�f.%�ى�����J�RG]��	j��o"Do��`�_�G�:�]�b�Vラ���K���|f"�=���Cޮ���J�p�K���m����K�Z�U�� �ͷ���_~֮ݹx�u|�5J�a��X�I2A���Rx���BP\.}��yv���Ѡ`��k�ߊ3�4&������=N�3���D;�O��+�߸��S��R�ػd�6��ap�ؕ�Y:!:�]�Q�{��l)E������%{]%*��r���
,>�|��2)TF�j�o#VY��O*չ��E5���.�"R��d>��43=H)��d��JD�}�2	^R���>/n'A���p2�`v[2o�^����y���ew#�ӏV�-��_��Q�����ic,(OA0hDA�R���|g�ί	�0lb��_� �@<1� H���<TFZ�F��n���O���ý���	�J���CUS[K��^�aCz�jL�	~V����k�
�y� �%-������R��£2����N��9��K �1���x k3P�C2�eZ&e�Yr=zʔ|`�p�� W�63>잔�,sh�ꡦ�A�ȍ6���h�D#jN�ܦ�r��������������Pa���� V~����^@�'qa5��҄~<�Ʊ��-��������$���Q60�aK�2���X;�P��w��G��p/³u��,ޭuh��Ǘ0ބ�L�Z�YȟXp~#�Ǝ�Al�b��|�>Y�@W=N�a�>WT�$>k��I���E��i������	����i:qYVk�j밊6~={b�����Xq�$�S�!��0A���k�]��F�$�_���� -iIv ~���0����a�ZCJU^k?�p�ei�d\�f�)׌y��x5���ȩ鹓e�q��
�{�����������I�t�6�]+�qO�39�< �9�2"�h�,I-,����{��-��ܻ�1���y��1���(���k4�t&0X��'�$4�e��k��#���aJ�_x)�)5���؜�,d�4b�[��7J�z�)�f^C�׶.�/@��L�؟S�� gVɟ|�5���Z���&���S.^捏c�J�UKY#Ѭg��(v��O��(X��&)���X�z_�W�Ǌ��:�B3e!/�Yw���J%�M"HԺ~Gv�f"L2�^�7.b	�����������bG�0ɫ�͑���/t��S�F?I��駬
�w��h���یb.�zB�	�A�c��q h����Z�������l͌���'���R��G��k�6)-�����%,^�d�WX�jj�}Bs�M)H�4������s����\3<3g���6��uU�6��ecc�Z�[uZ�ћ��G�!e�`�]~wn�)��7��W,�藿��R�??��%���8&�/}���\��?v{]��_�ӎ�1~N: ��nm2�orVZ���Ckѽ��t��|��ZvONp=w>I!�u�
���X����RU������c�d�T]g��d��yl1υ��
f�9�n�A|i�h*��tq����ԝ�Y�0!���|V䘶�naȳצ�d��e|o��cU!37�;�Y���Z��(�%7l�}V��ә5��F@�.�������CnH�|���-��B�խҝOn=k��`��ϯǸڛ��hn!�l���Q�,[!4�
1�*����e�m�l�+�-Q@N7���q/#����u�?-Ϋ��7՟���g��ru���N�u]�P�`��$� zfk"���!���"��i5L�����kڱ�}+��E;��x�x܏�����s��\�C-6-FD���e@J2Us�4'�1�Yc��[A��zb�aG9�+�Ȉ���W�
�h�ܟc��g�}�"<tx��a���~zu�c+�6���l�w-4J's�	`�8�KP���5A%���;�A���<���/�`K^#Ͱ��T$%�>�嶲щ���X����
$a�d9����6�a�w��Ǧ��ɠ�I��w���f�o�g|o�#���}2������¬���D�KĨ�e��y; )]>�s�4=Y�怌w�e��H0g���zH}�,��	31D����8�suÙ��\�9o�q
��C��I�&=w��]2��[8� W4@A�?{mj�)%O7 �����e��nu���R�f@�@`�zv��$�هԯ��fv���ҧ���Z)9l<�� ��r�������>����V"��f��V43��|.�GdqЖ#Q��zr���(+����a�B�9,�$�|,N�M��}�@�t:��g��T3� y̏�^ceVL�N��g:拵�ՓI���PQd�9��q�ٸ^g��&��nw�Ai�V=��Mʜ���Y�ܜ?�����re�.��4����;!�Z���>��A���2����_���~bl@h�#
-�O<�e�#���IO`�z��$��-Dw0q%#�,#����<� <WQ�W��Ç������T����7d���a�u&o��ho0b ګ��p���6������� jt/��`㞛nkD�����*�b8��a7du���n���r&7_nCX���
����5�jd�(��7�(+*FIW`w��a�'$��cSYpe<�o�ѝ�(!��Y{��R�ڄ���8�Y��^��Hu/��o��!���?�|M�C������^f��xS��g]��z�����R/�0R>�o���)d$����nxc�[&J-���F��w�1�}B�{i���_�@N�+�����O�z��h����ON�+;յ�"����`݈��O{܎��!��O0g~a�_f	<	�L&���-���c��`��P!Ii������xJ��5����ʼ|p	���zBe})^�݃�;���`?��ٰ(ۏWm:GR���KA�M���d�`��W�4��Gq�%iѠ�_���:�X��}�TL������E���P* ��%���+q<�F H)�	:��F��� �WI���̯?�4�>�:6�����C��V76��4�LZ#���L�ψS�)���z�ʝ���@����*�U����`		>�+�9�%C�_F�W�ݍd�[t!"��e�P���>e���Y��K�x�c'�����叅�D���J:s1���=f�� j�ճS 70�(��o�,n�o�z\��8a#��ׯt��?�a�h�w�4�o����l�KwQl��m�����*RCӑHX�������C�� 2�K����	6��@<߯KNe�^��{���^�^耴y�
��$�$h{�]�����o#-��Ӕ�>r:����Z���	{{!��;��!��s{%ƶ�]nv�&�����������|����Fr3�:�[k,�,��*�R�.e_���QP*��YS��ZZm����)`wnw`�� 2ʨ�5^ա��F��;c���	O�\C���	���2f��>��Λ͗t���K3���8���6Mޑ]�~�]�]I���M�>LN���2r�d�`������}l��f�K�}�vFW͏�C�8�����;_O�υ�?�^�i��ҳm~�3�ݶ	�8�3��y���~F�9�a%d�Uj�ƹ%D@KG���7
v��Vb��U�U�;-�5+�G]�ta�9�옉��Ƞj��/��$���݅�c#�̰�?�͒=/HN�ط�D-�M� �a�+0����D64�$����m�b��Q8.��W�*ݛ䭒�e�^a���Ӷ<9J|�XmЄak(2�\0�-�e��I��]	���Q���.an��J�n�z;��
���>u ��X��W
���o%�9+y���o�H�NJ�J���F-�v&p��4F5TZ�9��1���T��te��o<Iz_@����T�D%��_=+Ֆ��}�9��N�����H�7�ل�Lx�Gb~�R�
�l?�?W�6�>7.}^d�C��*^1��0Ā�iY�0}|Z�#�&���o��M����\	^(�4��õ��m$��(Q(I@��Dy$�,J6��
?�(�(Cᰫ3%�]A*��A�7�x��|�n�}=d��b�ov��`=j\����ϒ�>�� h����a^`��DCP��A�:�XU���i��t�"�G���o��t���Z,	����_���w�����C#Z��u�
�s�U�g �4a~T�t���^��M���<t����g��	N[����m.���9�f�70<	��(K'��4����Q(*�k�e��0�a��0 ����R���R���Y���g^��Z"Q[�g�#��w_�Հ���ogo��_��2�&���Ϭ��{��ž���J&w��ᄄ�W��u�6Y.����H%��g{f�J���\�w6�3����4�o�޻o^8S1����Yj�|�dx�"�q�$\�
�H�I�M�%��<X�*H7U�Zrx�
x�_��T�iğ뼓��v���kY>Ys(;���r0&�G�?v�+����K�N��>a�fœ$�Kl.� G)�m�vاD8W>USi�X=@����o)0����@Y�j%�nL��yv%6����"C��?Ơ�f�fՑt�ʤUxZ�ĝJB�50\��� #(-P�F���/���Ua��.=��;�F�D[:��7�1I��,���i�I��ܱ��ؕ{����$�0�0�Ӌ��}��_����g�3�Qš�O�IѮV	�v`�0���jk��`�vͩ����n�l}���s'j��?��O��"Y����Y��65E�}l����I.��!n�	�&<�гxϑ�V��W�a��-
:�C�sh
�*�;u��A��O��8_�b�v�	p�j�j-���'T��|����.*iI�c̈́��~-|������\���ڞ}��_���g24c���&��!§�9Oz. ��ȉ�E���z�RA�o`���|��-Q�dsy{�����4ɏ�p[t<rh�6[��PX�¥�|i@��4�_F��&N=U���E����_^�����=\Vo���Jl?��侁0�hh&�l��מ`+Ӆ(2�^h�@�ߋ2��˲�?i�8�^��ӣ�<4�=2)�n�0,�>��f�&�܇�Hh_�~�^@_�N`곸d%l��a�Nڟ��')A��2��T��RÒ,rw&(2�<Q!`m��&>E��k��v���G\>@_s쬅���wC'��;�H/��iEb[��Ui� ?�͙�|���Vϕi�����������A�dR�D$�!��I>0�5�H;tr\��������@�C(0�<�%ƒC�|�X�魀�H�:W�lNHCľ�6w�z1�j6��_bP�6uG�⮑�`tf>��4M��{z~�������wO뙽ye��4��g�,���B�`��H���Yz.l���RXin|@V�X8�,S˦d�R�1�it�g����=��@U1
CZ6��� �7p@�t0��?"~S��'vv���f���66I��c��2J&�(3�Pa�*�Q��,˗����5�Rv.7�*�HqY��AT���'����c����fv�?/ڜ
�"�guƘL�s���p'N����������N���@��+��T�2�^����p)+��e�d���v]��2�NU���7C��U�3U�;~蓷Jn�x��\��Q��u�5��!� \��U�ߌ�Q�$;D�O�²@j�Ԣ�+C����i�PS,l�o E"@i�xV�F)���Bľh�F����X��QH��|�A娫Д�Y�}�3�e|�є#�*ٺ����[�~sK��%�u�W����h�@����� �p3�@�)�I������A\���B�9����-��2��&�F�`D
�D J��_mђ��o.�8ۖ�ƫF��I�HGV�"z*u�v�<a��O9Ѱ
K)`_l�|DF?+��nG����*�������9qW^Xf�P6���	��ߒ��$����IE�Y���`ύ�ǝR���]�R�s�V �R`��ROo�^�M�)�� J��j�[[^ʲ;�Kj���������Z�?�Eaq�����xf��E�
,���J:�]΂ ��M 2�X@��/�e?9��p�̤�Lc��D��#�Q�t�2F�������\��R��;5or�n�]�� 1 I,	�������ֽ�dA�p�?�x��$t��#�za�$_��W����x���y>��¢�P�Y��*!e��1?��"�G;׌ݕ���-U��}ը���� �`�G���#*�E "&����sF�����C��QS��飧R�[jM�drfk���eܪ*�arU4k��m�ZEE�E�߹���H���s����}�a!�Yg$n����
�FҔ�ʚ8�q��:7`j>��:�;Bw�`���7������OР�����O��l=�$m�	0�G�G�	�P,�7`�6��jR׭�ͽ�Zd>�����
 ߃s¹�>�/��	K���xnQ{�C�z�I�������PZ�Г�V>��l��b��R_���ه��HQPd^x^�jsc![|J�8����֭�NHU��0�^!�!��Q�lX<�����edf��ri_� �m�ɏKdQ\���KӔ8Dx}*���ʨ��+���XRЙ�=�c�'���9Ӑ:�B��]����i"�q�0?W@����B!�E|~ 5Tu,,�Tqh�W�N�mͫ��YrkP�.iy��+m�6<U��^�� �s�T�Ӛ���D��D.b5��u�@e�=�8D�رM���`¢��,�û{%3d3uk��^�@q��ㆾA;�&�@��G�^�$�1�p����>���$��#��
�+��� �!�F�nzǉ�|�_tZI5���\�YL#2S�z���CS�����&�a��Hg2s�Z�)��|�i��:�b�G�곣Am�Nfq�Q��|�8����P�)�pD�l������ug�bOw�0q��	xD���?�'��N��F�g��C�����u8Y�}��$ϭY1��۪�͞w(���FH�G�f7��=`�ܞ\2���Pb?���<�M���o�%�|�gBM
�-���1�F�t��x.
�y�?���ߪ�<��'3vХo��<��{!Y�j��k�:�j��^iJ׵���op��ΰ4���µ	%�����@B�i�)�}�Q�j�쎙3��=��%��f�)Y�v8���IZr�H�)g|6�4��* ]�L �|1�Nt.����Q��C�h��hi[��&�]��S��"����X��{���uww���tWo/�V'�j��*��I~ьye3a�K&���̇t�+��M�NW8H��E���pw4XVp�*tnm~>����Qfׄ
����z�W�p�����?Lv%$	 12:��A��yT7&�M!=`�g���l��l]m`��Z)j�\���)�9�*�&a���C�I�Xz�����|�.F�eh? P�K�EO=�����-d#w��>ǉ��M��tIU��Q�b��S�C-��H8�x*�4�ڬ�E�����X�!�I��;��ڠ.�jC����x�Kb��7B{�iMƯ,�����NB���;b���w�E�b�[N��fzRR�'%[�w��ᖚؠ�0��Iٻ�gO	�\a�ު���z6�dL�Ut�Q�|6��0X7h�E�l����YKVt�̈́o$b<M�ښ$_���|�FV���Ơ��پ�뼹Mj�҉n�hԝ�PHK2���[ł�I�8aP��2kO;��q
���0NP|V�-"�e�u��C��^�T�{�ĭ�VJ����_&��@(�5���C��9�Al}��s��4�{���-���Cߜ9���$�sQ��t� Q9'@y��c��8�l�����N����I��7�y���t�?rp9r�ՄY����^2��6������A��G�n�,ƌ ��<nVmf�V�@����l��YU♻�r6ķ���@��ɉ_A2宏x߄�w�}(~7�&Of��`�WDHc��R�[fyª�2m��ȻA��5�Ig{@�׼0�^I��'�2j����}>Rl�1$���oOG���/G~��L���4���O>�"�Ue:�^�����'�}Q�יdW�p<�����9�O���X|��}Zr
���3d�P�@�RC���P���"�	���H_y	��Ĝ�� �XHi��R�ɥu��;��P���FT�3���ᐆ|�_��A�qΖ�!�(�>�P�w�uǽ�����Z��-%�-��O8I/��[c��B׵G��51B���h0�$5칏Ŋ+c���Kim<����T�БZ�����U����/f��P��`��+X���)�&����� ՜ֺ�� r��D0�	p�y5����F�����WjC.�7�'U%�O���]��/lz d@��_��%Gqg2�)4@���R��&_���f�����B'�4�0x>��f��D@�W_T�c��T�^��Djz�jI�4W����X�|��u�CS������,�n��D~���D�VJ|�yg��
�}�R�b.�[ȗj�Ѵ�4���]Z�~�֐���Mt�C��d�����x:p��I����p�S�|1\DN%���H���-Y�K��a�E�kg��H�ſ?��!�y��Ь��xeX<�@¹�����Tؚ$��(!φ�e�nVW�D���6a�3�֗�AR�hO��p6ue�֌�Sr,6T�1I��_h0��0nb#��I�/���C�+)v�t��yC��ncSR�"ˠ�e��[t���� t5��1�)����+�k%#���2��Hi���D������)e������a�v�c�O2S^}�aJ�� (c���8��Y���I�s��<k�k�&�(�A�q���������Ku ]��H����%�o-?�v��U�y)g�8�o��V{'@�{����Y�U_�9�� �]3��IB*�s�� I�ӷ�+�2F��bjz�,5�GP�o��'����U/�mzt�6�4$ƥ-�%�^����?�O|���h�Z�tm�}�I���I��B�����rcg���脀дk�L\�x;;ڔ���A{d� �T�ȧ�,��VԆ{Z�
�����%���d�ZhK�D|Q,	���qn,�FH�V����=�O��:�L�9���_�E�����J�^�U;
�d�	���W,;�������|�lo�?�8��R��/"4��?F	�e@�6R1�L�rs;��!�;H��E}��Y�_�������*D����ҋ ��qꖶ� ��jgy�P�h��LL|��+��/�̙���$	D�.�	�.'ǣֽ�"W`�i�n��	�
I���3pf�&�pY;�N�m��}o1'-r� �Oc����8L��h2�1�8�0-s��z�OB�O��H�;bqJ�Oz�������I.b�e��,"���%�.nq'dr����~&���0�c�۝�<}�C��ӽRjʕ�D Ks5�3�1L�
G,w-��2�vu��m>o�a���%f;*[ � ��NW����(|s@P,�M�-�!i����}`���$�а�*�,AëǍ�u��lc�^����KХ9;",����?$ߨ7��#��=��O$y�vvHF]�D���^N��I��+\�F���Uf�I�����[r9Z�2iѫ:�) ��C̰3w��=<u$��ϱ5�o]�Ϝ7�� m}�:lU���t�nW���~����%N#w8�7���WKZ���U"Ȝx���s ��@K��\�
���ۣ���
������K���A�_���p�����*�e��b��dcT��D|^��|j��'g�q��֜��"%,W7��.]����4y�:�~����Y�]~_m�n��(�s�w,Hcĕ����g-��1~`��ڞqJ;�wn��J����zO<F�Gs��1�'���{9d;��ʝ=0徥&���C1����Ƴ��š��/�+�Dy~�Ϯ�.H� ���o/ϸ��>�k)���\�*�[�5�\���pBl���f��ڹ�~6��o�����l�7$���2RU����&{�޽�@��^�1V|��U��,,�\*�ZޞAq(�0X�o���Rw�q[N�e�QtvF�O�:Z�]�3��LK�Ѧ�&��#���,CO/��#m5�U��/�z���ۨ�����w���ke5$4��6j$�����4���LV�ua-�=��C�����L�"���Q��G���^��Ёq0�N�ډr��;�7��~
:>������|���Q��������OOE�[�Gg��R�ma���
{�4׽9�x	��O��|ʺX�����ac�٨��5QQ��e���v�C&R���𥣻J�A)k$[/$`x>��_�o�)Ώ)����^Bd���标b �y�������KdI�(����o�VGWr��J���O_ڭCY�u:{�7�}S�����s;�?�p\�t!X	/�koS1��R����\��2�p"��@�Z��r������iL_���RE��9}qT*[���老�0�zG���ԼF��3ꄁ�,��L�#f�'��a¢5�f�_O88�*O,P�z���MB΅�GO�%���Ɋ�C3 t��{t}f0�ut�\���7�v$׹	{$K;��c4��3�İ-����J����U�c	��z��͎�rU���0`�6���'0Ζ�˷���(�q�������JW;�ka�ܿ�'��ڌZ�K��
0v�<?���#������@�|z�gu���E<�"�d4��P.=)�oun�F�ӊB�!ڃ�R͌5���^�uV�z=��,��M�������,�qv��_�4�S�7�4���������:T1q�tMP"Q�D�C���&���_�4_�o�y)�N j�����L�5�R�&�����%���7�=5ͮ�]��{GY��l�Π���*KX�z�# �WƵ'�#e"����պ]
���&m�r����Hj㹚��R�;Ȭ!��4����YH��M@� �t{#�m^�YMT-��Q3�5���j�lS	ѯ��g@>����Z�\)y�䈡F�{�υ~c�.l�뎳A�Դ䕙,o�1� �S��A�z�.���֑i�79A���}��� `�V� �]��`��,�k\����t�PGm7^<۝r���	X�����S: ��"ݹ��~w���"`�-�3��N��>2������
�0���;-F��}fWP�M/���57���Z�a�Io���):��!�A�An��xz3�{0}P�o�IxS�gNs����ox����B�U�\���@����k�ϊ�'#$	3B���'	�:s�˺G���X'����1�j\�&n�!��ry����)<� �+u�K3ϡ�d�Gu���y���Ft�D�]u�DΑ�pp��(�����ں��9:w�V��9=��>�H�ô�g�>�e�T�ŕ����P���?��8a��nY����).��?P��n��(>���w )OYY7U\~Ai�H|���C���V���b��H|C�:�4c;Fߔ���uKcȗN�g�����pe2�M��<�ɇ�L:u��\��%^�^U��Y��݂��OJ[!s�W#č`�z{F�u~)}}i���<����0mJ#���Fw��!r� �a+�ys{��W��t�g+z]�	)x[=��"����������.1����w�4�5��X/���uW�@�TF�V�б!��տ���\$�x��TL�r>���պե�ǜ�e_�E���#���3ƍ!8ל�2ng�fU,(������V���"jX���l?/K��>ST��m���;����u�-�Q�)x����-#d�w�Yk/���n߁N�_��������mXi:*�Ped��������'d�Z!��YB�#%1��������x�m��n��ճ�n�$��[)i��&S�W����J�}i�/��0���ޖ�P�-�75(.ȶ�Ձ���/�p����r��X�v���OEԬ��� �}��^�BᄊiJ ��0R��R���m��<*)�'�Y��q���lf<����8�������ٻN��=X��G�C��P7r?���ə��R��?�����s�	ْ��Q��i����H��2$�C.��O��
RqRU���I�W�i)Ԟ� H%��-���d��VAOkFX�7{������]C,k��Hm��=����O�η��hM'�����D7p޷r����pc/��(yo]���>�����kH($_%ϰ9��+��l~�l����U�Z�z�(�Hr����x̐Y�-U2�5�ϣ��C�M�<��`�t��Q�{�SI�a�{�"��YD��v�=:��{D�FI�γ�
"�p,!*�</��)Iz�R��fw�A~jĬ�+^�%�{k�/Bx�{aҏQ�]\G8�V�':�c>Eݻ�J�$��$�+
������� �g�gC!A�q��>�z�W	Z�</�qKy�D�yXC�~f�YK*%�i�p�Ϊ���eK�;며��m���?p�ڋ����vH$�v� ��>x����@��>��|��c����?�jZ�2�^��z��o��b�N��JE��l6â�Aݟ�b�P�rfB��PJ+�{`�k�ڨS䔍�D�r�f�:�s8��8�u�͚��+���{������d}H�'l����)�i��x�G<�]�N(�e�_���r)/1{aW|�#ш���ي�f*�	��_ �i��Y��/��mYdT����d �H�cI��6f�����%���wzjd�3��]��_Y ���pXd|�_�`�
��W�}J7H�o|n��f��i���nS��4ض����ngAC�w4�o*4-9`!��C��FT�*�b��Y��gt������M�95��yY�P}���*RH�!ZI���n�p�_mU?��)�$����j0�o���
er�w5A@��[01gR%�F@3�4��U���>��!&��]p���s�Dݣ����1ߩ��I▋b��R��=pk�%q�h}��켃�$�!�>��g`���\�d�-�,T�s����З?��V�|>r´;݉M�?��\���#�v���f��kkkjn$BQ��o��H��Ow�u��xd�]~!�܏�F,Y�º��앩� GB�ev�֜̋+u��rn���Q���h;��q͙�TWM��>����Z⛶F.�OX񲙌�{�FG�Yg�Tv��?vd=�O>h��kG�4�AX�� ͈�aU�>�H��3��㇀ۘ-�g�(-��/�{G �fA�����~E�mMb�t�=��a'�c���
��/t���@~�i���;[uF#N�b�j�E��,�\@ϴ�[EΛ�Edf���Lw�!��+y��[{v$fw�>PY[�/�6]&�%�8���9���7�T���D�(eAu�US�nEl�w�x�CU�W	�;��@�>���}n�A��q�{����b(�Ȩ9�x��e}l8���d��g�D��B) �1��)�@��Qb"�L?ݽ�L��|���K�m�l��#
�A���+U�5�:>Ձb��al(��ѱ���#����\����N��%P��q��(;�����2.ȝ�=�M,1�X��v$��S�0R���&N�MM �� }k��ǃ���(��s���L��>�s�:O�`7�GA&w���d	��ELg �Z����b��F4��6��Q�*�r7ԎG��+�&)�^��X�W�.�fX���\u�&e�j?1��a	��{ay�%�I)1$!ƨ�2�Ȍ'L�=L�E����:���K�p�t��e�E{{��v<�iº��7�h�C\
��ge�7��W3���z
Fs'5p5�xl�_{BJOw���lt=���]���LY$�x�f�6Zè.F��Y��p��L׮�T/�U<n�/�^!�3nQ؄Iy���1��Q����[�}�T7m�����O���`4�(z��;������$��3@a�W>�^O���4:�R'2G��L��i8�1˃S���`�cֆKw�L/5į�ƨ0�K�����Y�j��_"��rAwO�#	�,�>�)2��QX�9���&e������"��g^r�)\�,~q_B}+鹚��ڦ��*��&�J-'���A0=�3/�6J��k��絴���nӕ��y��g:�Y���`���h��C���6�z��E=<�JSΑ�9A*�&v!�%�����*��Z���|ص��݇E�x���w�b��:�1�����(�����#�@���|�/a�m0f2U�"�����s��z^��~ "��͌71�%`�H|K�u�^Nz���&�š���G[%im���V�A�t�M!@wdH����}[�m��^��_��9�g+�rؓ�+��Eh���h��H�ˁ�û�l�nR��[�X��)/R���!�CP'��NK*�X���\[���i���+'g�����ӝ�]��ir�����CR� n��a��u�CK�J���ع�T-����Y@�+�\��Gw�sļV��`%�9_��L 	��p���dz��p ������5`�z�~��Q��R3��,�f�|ѕ_�#��h���*O����	S�rᓏ���߻��c�g)fi����C��ij%}�����V,���9��6$)�<lm��Ò��W�`�7;��oӥa̔��(�)t�N6Ko�	���\M3�p
�����X�	WF�ӟ�V�#Y�--m]��0�Ln��:�0Ц^�a�I9��R� ɩ|���B�-='7�����nL�O�6X#$�L��!+`�����y׺ d�+�jk_�0��h� �������#�̮��Vb�`���J��~aQ��G������io\���!}40+�E,*].J��c�`�3���a^���nCW9n��G ?�ƛ;O��+�B^�e�}����4.�{�r�=��N�,�J316�2��A߇�S5�?|��iۻ��-jɿM&γF�z	
�.�qk�Ft��I΍�5��M7�b�~����=c�n�΀��y��\��J,Z���\f�5(��.*|U4�%f�
�nG�c��6��cv%��_u\�1��h�D��aE 
w�5�@v��,]E#�����e�[J,*>�y��ʠ�E����~/AT������"�)��/�&>@�_b)eK>ns&p,�(b�����h?�+Yg����9��� �U<����D6dG���1���Q�	E£�姖'�^�J/�{xb�B�
��긧I�$a�eg]�f3�~���'X*���`�c�NS1����1�Sg%�U��m�O�<�d�l�(�yf��s{� �~
�"c��v}�e`vI4��A蔸����Q����_��_��l�|j� ��f$��5ڪ��&gd�l
V�������ڞ��x�ې:�1޹�Zm)�&�l��ʠ�ް��U���^�<�7`̖��*���U6���
ڽo�9�����.������Z�8���3����8��9��o,d����HV�I�3b�.Q[��⢛����vv�B�b\����Y0Jڠ�op����88��g&D|:���w6<~���� �K��>�_����� ^d�]F�'�;w��&�/Y�w����n/���d)S��Kd��;3~���Gh���o��-9�\���d�������j�Ts�_R�ۡe~�/1�`ƥ�3i�`�8.L�%�ٽ+��p�r���̦��k�R�	?'"���wi8�h�k����?��$���y8���3�U��La|�6�1�X�Nv��8��Sd0���F��D�T���l�����f���5bǪ���U��ALXpm(�ݑ�����*�jo��g��_ﺒ;�+���!NT�W7�KbqG�C���#$]8���NU:���v;�~��`�Нq�r^͢��0���.�g錁�%�#��|��W�8?�<-��$�I�+��7W�6_�Jx��y�*��r�ֹ1zNU��+�հ�Y�ۀ��Q'��[f4A�]ڤZ\���q
C�*hA��.c?�m�U'Ͱ�}�H���q�&V�����ˮ��r+V�s#�eW;�/�9�l2��F.7�#�7���5�Epq�yDr�~EO��$����ei�/�*�D��}C#O7���g�bI���ͿX$!� �5��d���O��1uc���y�H$A"�Yt�_r�N��h{��l�.��ދ����������f(�fAG��ŧ9���P���26.?�hg�k��b)���	�?��PzQq���<�cRV���(�����_���V:�/��v@5%���=,�u�0j�����7�0�x�I ��j������9͒�)_��K�޾�r�Gؙɳ+~��ߙ����΄���ל͏���+�y��V��!�,����_��f�+�LC&�Ӽ�{X��k�V�{s�sm��|��D�S2�ժ�p$T��E���쩩v�v�Y�R�'ʊ��݃U$�h(p'���a��'�Ao���g�Z��ٺ[ӛ�����q7�0������S���d��-s3��d��l|�6*��";�Ճm��2/Q�G1��d5�M�2֭O�SXQY�-42�,��c氪�0!;cw\X�}��Lh�.�]��a���z�w�:P�&���ٖ��H��=�@؀ݿ����XI��T�@��n�J�������40���ž�΍�7�R�]Y^_� \7�)0�SV����:���=pk8��N�x�<�\��~Ͼe�IPH	�r�nΒE2��T��%����v��p��R��É`�YnQ'X��B��VEs8�8ܫ��6�z�Ϻ�������w�+�7|����ڔVɟn�3�Cl��1�{#��tg1@%Õ���I�m|��6����6`?�Li:�6h�a�[�y���Ԙ�����A�Φ��cv�MQnA�ۃ���Opv�����Np���=�LGr�D���R��ܴ��vI\D��(�h�/*�1�t�NL��+8���މI�"���9sx�N����9�	=杈4��&����J��T!y�so����L�~3獗y_�X
�7�.�Ԙ�h1���ȟ /��,��i��0l��m�b `z���n�{M�{t�);��� ydF�47�����~D~�d��[��Q�{zR��9�\߹��J�
�� o��:6巣�!z!�³i^輲�{��roe��q#]X=>┽sTw|�+Z�����#�����n�Z|��(}�![خZ�|�>�~Q�mo�w�;��Ȳ�5�X�a^)[0���pO�-cYQ��xCzCRx���`z��.ʣ�`��ɲ#�Q�,�0���,.����x������q���Xc�y��4��oP�Kmj�CpI*i�iǵ}��,W*�BL�����s��)ݞ�-�S��~��Ⱥ3��ϸ�6�=:�b�y�>K�|�����?lMc�ǥ�{]O�߬��{+�?��=�?�y���C�m�>r������2k&�O�hG+�]jJ53�e��
v��8�@����o�>P��z"���%��|�Fw��J[}���睨��b�X���/Cǰ�Y�
(�V �lp:
&��;#WQ� �_�e���w��� ��g(���N�	�}�8&*�i����?��u\|�DB��S��k �;|��N����"rj��R@���kΛ��OG͌4��`�_�*(�쇽h3��_xԕÌ��K� v��v&��`<�$I�Ηᎀ�g��S_hޣ�o-A�sqh���
Y�eyzjD�iJ3�S���N�rŸ�	�r/�j�8F\" �P%R�u���L�B�/�
���_��!$�~s�7c����>������5�t'����>�ua�,s��b�3H�M���S∱��ߋ7���#��o�5�zOD�I�|�xE��NN��3���Y��Ce��ݺn6�9�I�ǅԖ{)���H���p�Hb��v��K�{Q�f��K}Y�=V��������h��k3rK��,�6�p�b���7Q�(�y(eO�A�P[�S�7�5a���'(���]��I���[�X3pE������5d�г_ /;���;�}�5��rnA���P�Y�ېy�(��}R�қm}��o� h�X{�HڶZ�5��T:I6�%�-�+�P��W�������:s�[�R�O��V��?�'�}�Y]��ἷ�a�;Yw��L�G��iW\�C����F�p*��г���U�x#�H���-[��neڬ��\h��"�sdǴ�m����� ��rr��i����=�I�w�ի\^�i�HZ1�G(#r�r�g��Ȩ릩��Y���c�w�ۈ��u��T�j������@	{׷A�!�3Me�^+Y�Z��*���#����R���c�z]d�UL�bf�Yzy�ys�q=�zH�o0��ρ�HŒf	�$ລ�5ê���b���SH��A1��D�m��aW�6W&U
��Tp�`;����ʁ������.�fz�/�b!a@�����TPO��K���3��p�.�1�[Y'km5MK7��Ƥ��Vr�����C�����S(�cVJ�Y�!
�y<�"�)&�e�	�
��0�`|B���u8�i���+:b�ƶhJ*c��ew�ᣋ{��'WH��%��o��آ�T�5���{/z�G�~'��J�`�a�e=,M1X{�+�Tu�A=�Prޞ�W#�(3&hU��K�:m����}(�y{��c���j��S'ϓ��丝^aj����v��'�'�r��A�����S ����Ȅu�B��	$��c���2y��-�Qِ]i�-�6g�,gḛpyH�Z~Ƞ��q���ņ�Q���GHb/�K�2�]����S�9ڕ�Ʌ�5�ƭ
c��+ܭ�zG*��M�Ch�.Jx���s�=��#�p�x����޳��-w'��-�r��(E� ��D;���"�^tyl�as�lu��YU�b߈,�EX�^�W�ߜ����q�%f��8�,9��c�-�I¶ѓա6KrE�8�/��B�����Z+�:�1�k6���B`�!���������l-�Ad�6Y��o���tڹ� ���&�\P���1E����RE��:���O�'N��z�j%����3d�=�C�ې9ģ^��-BV��iP\�]�j��l���d7��1�L�a����B�bl%�T����n�ߦ��~������-�:�ٍ�^$���뼦�/	����D4TDhgy����g�#eDY���|Wm;�<�m�4rU����x}kL����cO�R�U��Q�������l�<e���*�;\R�J������'�u_�6Z���KKw!�th�����]�ߞ��|~ߺ8�U�Z�Zw��7ҟZq�YC���wL���L�g���iۥ�NU��}t���iW�.�7���[dvW8v):��s������#�.���#dc�I}�6���5������xn����=�Ó���%�U�Sm��E����kl��XI�[gߑ�Om���o��#ᓹ�8bw��*�䜯y֌�v�0�r�m<�5����A�{�$��d�e{��kz"�D!ݲ
f՜V���\ћ҃@�.���b�N!�1ޠ\�V������iz3Fѷ��s9G�}���We�:��U�G*���'���u]��k��v�6��m�L��c�wC��,z�|_�fz����FL�[�ꅷ�@�v�'��!��U>r�\�vzf�^�p���|f�k��m�0ÿ�'^���-�0���1���(����G��	£�'in��	�eN��9AjG�:1�����oc��.ڳ����MKĂ�>ch�}�{��ƒ��g��!�f�Ql~
�^s+�j�Y����0~�o����D����l��@&|!r�����jF�-�D�	M���.�KW��j::8X�.��z��!�jF��y��W�s�4ϵ���.��Ľ ��?�Lw�Fy֛9y\�嚂E��h �@���\��Y���u��{���]�����0�=�򴤧���=Jf=�J�r�*dP�H�$��J�4�7�\i�wN����� tCC�ox�詅�hd
�(Md���B]P����s �c��4�!
�l�N뮅~ڱ��#��Ȑx6ra��1"c	�Dd�#(3��_�\EK�Yj �f�z��3�����d�}��N�)�#D���KFv`��S���3ZBeq��E���o 软*=�#�J��ްfh�r�D���ˀދ���g��9�`w�5<HJRd���˵��$��gYj�|̈́��<��{|�����'���==��NҬ�`���u�BT�>��D0%!��a��1��^�z?(V�H��DH�+ɵ'v-��x����vF_VLq ��i.�|�Bt�v������X�����é�|�_�;����Pm��׭�8�7=�5���Fs1`(�
k ��~� J6��P]ƶ�2�P�T+H�F�W8I.KE�W~���Jj��I?" eW�
�����S��y%=�m�H2L�̺��1�iUI�v�";C�7MPL��8�w��
xM�z̳}**�'�- F��]����l���ݕ����w�q���="=:�aث�G�`���� ��zm����)�>�����h�q�L�Ќ,���p�u{�%ǰ��m���&��\l��k�pݪ�Z�����"����1�%ޛ~	�g73,|ʻk5�p~~�[����D
H�p�j�gV��o*N|�,I�~�@ �D��X��R�]���Jr��:�vEȐ{sm�JI�ކ�8.{e�jf>�Td�m�}����Z]O��2�J����l<́�&5^��<rf���T���d�bA��Ɨ3��G �z�t� �bU�b�v��QF([�݃�Z��fT
��_�K���������.@ ��{5�l��j�x�)R�ɹ/����:'�Xi�Pu�����9\y�/�8��Y��D�s�����n��j�+���ͻ��ΐ$.�`&fg��Q��9�� zn�U�F��Z�A52��;a+�i*,�yA�u�x��6Ř`���.�d=<2���^��A�5�Q�n�?��M�c.�]d��fPzQ�ƣT��k?��h�=�Y�����JI��0p(&BN��}&�lu�q�zq �cY'B� M`ٻ�:�;Ё�w�ez�D�U���E�icLY��I��X�)���Il]Gx/�R��$K�ծ����S�J%�����4:��~C%���親�Z��o��@�D@TK-}�vO�M��}����n"3���+�YV��1=0Y�(�������- ��,�� n���+�e���IW6�u���%3����P�l�Sf�,a��<=@H;�W��T�V�x&5'2Yki�م�p�c����zz~��y���0��'��=�������?b@=N�|LVY�&�;����˓uJ[LȌȀ�R��}��_�n1�E�����n��|�!���gH4��b.�om�ݍw�~�S��L��߇�ib� ����n����%�Y�B�s��E�U6΍l��`����$��M��(�>��Z�A�wӡb�-[&�ch�X`�i��!�=�%�	bO)X�7������Z�Ûr�Ey�V� O'4<���⌸�Ih��, e��+V�r�g�`'��v3S}1f�5�ov1����ra���A��*�j���
�E��oGdz��`��DQC���uBq����>1�跲��6����ݩ]�M�̔f�O�3��y���,�lF�4+���R�Y}c��������[�?/&DrAe����˝mB6�7Q�#A����2�̒��W���4�}zOrnj80:���}����u�#3�L��E$������ُ������N�w G�k����Gl�
���B�:y���A��fޤ:#zղ�C�g�S9gu���G�&�̑�� �~�-姄��٠���0�M�sD"L�$>��Ԡ�^�#-fZ~����\pe������1�����k��������D����v���y,Nf��'������k?HY���i�뭗6�t��n�T�����+�PN�i�e��GyŢ[l:����}p`���M��u(�
�䔵F��C���x�&%�P�#7�WQ0C{"��W�o�`� [<U�
  �P�gD��e��I���)X�8(�!�%0�9�S6�];B��l�9z��9�KR�N
l��-ա(�
��Ƿ-r
���4e��7�����m�r� ݇ej80��LΠ=w^����T�j�� \
~^�����Q�7N	��]!܎�M��մl��sҽJ�c�'���M<@�8j[K@@�@�b~���-ԃ�EEP>Mtjg�/(�BcC�4� �#%��+�{����3�3�C �!)N�(�01�}������%ͧ(W�nIf��+��O�BK�m�it�.6�w�U<��ZC�mWGGb��AQ���M�-Q�����'_�.��l��G����w�-��~���9u]��:]�����y�|U������{3���`�25�JT��f�����������Wߞz�Jh��ߺ��)���e�Xz��`U��蕩%��!M�q5IJ��&>�����ʒ����QG�։D@�����D��(9Xl�V�!z>�����1VE}��kD�K^��i��z�v=~���Z0��8�t 	�w9���0&�/�P#������ND�S�������Ъ̼Az7�U�T�z��B��ʂW����T����i��hD��GJ���}�j�p�I�
,�5~Q��#p2Rn�S���DF�	O��Յ�&�\KEtRٕTwĭP����S�����ChZæ��d��x"K'$���ɖH�� �V�Ȑ�����v��e�﹭��<Ղ����{��De�<|��b)2�:����zD��1p>�EX��j�K"c��^���'1�f8>}��f��E�`�=�����(���K��*�lً��ɘ�3Ӌ)ʛ���kpZ�6'ׂ�Ԣ%*p���pz���q��_�YAl� ���\������[p�Q�+�;�D�\U�uREt?zEFփ�oȩn@�8 �F_#W�\�[?&��'����E���3>�R����X�)]�5F�E����鸎�X��~�(Y���>զ�P�冞tށ�Ͽ&Lk�X?aB��+A���l���Ģ@��[B�)��]���4�R ُ��64��v�łL'��͵���0@GI��!ہP	�d��)qP�O]��	�e�meM^�!����dl,l�Xo/C%�|}},�K��h|��@���g��̟�N��-��~:'�;$q��WRnQpp �k�V�e+C��pƚ�A3��S�'���/s��ރ�#8E���	����=��֠5K�fiu�Z��g��[��P�UU�L���A��l�eB�wV��@��Bɤ�8<%�D�`�-�$8�S�&Mj�nv����Ὥ�)a�Ǘ.K)kj,�(�~�O�QO.לe�;S%��,�h���c4�� Tr�zp��d(,T0��0�X���/8��?���3��!V��81آ4�©��W��[�QC�V"���ǬxxVh�(�b�]��,n	��W�*� �c0;�H:"0Pn�bO�ٲ��m�$�"�a��Eʢ����]���cP(E�+%K��[�d:�v���/6!KJ<^�{���\�R$���
S�q�-�oOq�6&�ÈB�x �޳ O
�cK<�w|#�;w_�G�-�8̿� �aC��@w�k4z������U%��e���^{�(�j�_��T�Qe{��u+��%�&BLn��P��~W�6�����*\�٘��� Hw��I�>��G@p�i-(8q��s����V~A#�j`s�+�9���̆�8����A�oW��q�h�&U���������5��_�}gK�`���g*#�)�ei�!�HJʳ�Ƨyb���T�]@#���Q���j�v�x�R���s	5
�%�*8�3�m�?iO�H��ˡ����/�V��9���*4Qԑog��3�Fm�|�9;�_�d���k���Mؼ�+�zv��d(��8�� �Z�����x��;
|���+˃#�C�E������-�A%P0/C|�f@�d%���7	4Ȓp^E�ȉ��4h5S_b��fa=�"$wm����T�ZЅ�6)��[�>"�vE��W���YJ/�I�_��q������N�o��N��'���k����JN1z���/�Ę�#1�&´�-��3�&�=�eW�EC^�����?ȗ&���#$OoJO�x�'g���̊S���A��*���j�e8�\8�K�Z77��T����֠�!�ـ2�#˩.]�U��o$�g�t-`�8"�閲�e���F�B��O�_`ڕc{���Cv������;�y�\�N�Z��˼1��\sސz�\��5y#ͣ^�ȗ�O�G�d���ύ�7Q_/�w2H��;�ʏC^C��g�NSIe߻�| ��o��(�Q�H����3�+#��&b�d�|�1��3�ߢ��/י�[�[�N�b��Ֆ:-g'��Ъ&����l2�i��&-�:R3Sa$ ,�2ۙ7�0��u)�l��9�Xn�R� ?�.��/���Wd&8)]�[�Y���.c]5]�mE+�Zy�6،��^m�HV�����}d!Z�^e�SM��o���?!�M.�i��+��+0Ǯ�&�A��>qٸ)������n8#�II�E�95��KS�vpF��]-͞�Tq�v�Y<�~�J&��9'�-7��`ژpa�U������B�^�'#HQV��<Y�6��T<��#B�����vڿ*@P�����j��LS����s���x���;�b�vg%����[�p��ڷ&x�	�\�@{�bۈ�hK�U����5��G?:��SC�Zt� ��?����������d��=�Uؿ������U`{���ew:}N�J��zhQ����m9{�'hA|���َa6���P��U��{�0[�y\�6�+i����A#��n�9WO�(��屟����S$~��Z��U=»�f��0�e!�@��k�
zJ��ސ:�P��uU�m����v!�-כ����&"X� dA�i�y�}���?�����W�M����J %f~b$N�!<�Zs��]��;�c+%��*�8�|�w���̤�o�8p�˨�m��9矿S��M�T��3�I'�z����r���da��o�4������ز�m7�JK�[� �2G)�І,Vд�E�%�|n늳8�f�>�UMB�Ԭ�Ib{^@��2�d�z�#G!��,I���t�"�-\>�#N�0�9n��6���]��V�S'�Q�V���E�b9�7�jB�V�Ț^��U�5���h�,��@kðt�S�@���ȧa�:<��yEO��,��X�
m���h[��㸋��wS&�X_V������0c����
Z9*��c��9���)�<\��4b�6����ZR�K��z�m��c�ZS�쌕/&$ihu�U|:��b5`�[&��oΊ:�F�FlF���*c����".|r�A;r
]�n��eј���_gT�'��c�~����KGx�;��=�8���������KG���An�Ѱ�bj���\�:�؎[������;<��7�Og�NC����f g&!Da�ލ�CT�n>v5���t����6=:�l0��'��8�����1��d�#��AUΘ�D�����>�wѐ��IPV&��®]�g������M��#j��wJ�k"ɯA�=>q������!�OmF�\!,�r�#�+�3����%c�z`��qDժ�.�-p�V{�z!uK���[�T�Z�H��D��H�6�������i����Y���`S����;�������b�uaU1���c���QiU���'og��� =Ny9G�9�C<���̡�%n�Tm�����?;�߮CJsO*���EHiX�;J'�4�����X�9�5���S����#ih�j�o�H]"W`��lF>������'�F��3,��q�C	�k�c&��A�)�@�Ew������$O�gG{A703�}���A]:<���5�#������$�g����ˊ,�4kP��$>ߞl��K��j��-Bq�W��<�j��k`n��L������Κ����?	�t��+T�j�9����|Y�Wl��}&�*�o~�
 Ȳ
�oX�1�bˆ�����ZCזR��l�����SΑ[!+YR��6'����ytlqZh@}��hU�=y�	Y}���|�����W��������E��=�R�&1N�]�&��;�̈́��J[�����.kJ�:hn4-4>k�+���[�O�^���ol'`����)�y���[R T�fk��)�ָ� @����/Z�j��#�܅�y��T=b��}�c!Z>�ey���@t�Is���<���"��V�P^|V�I:�ܰ���2lS��~t��u��?-Ϡ.=���yu@�eB�L��� 'Y8�v4y������Z�s/L����9�T��B~.�p;�af�"B�xZɊ�VѶ��,ao>�����ěpj�m��>bA& �}��ϑs�@a�fތRyȥ"V�'CץNd'�S��N����b5�e����QO�^�yG���dv�"f�U]x5Z,��|�n�.���4��1pVZE��(j�܍I�8C᳄��j=*Y0��Mq�E؝l�����϶��@��s�)�l�Qzbh�a�A��q��0�l8�V����@���1��q�,�G&���-@����l�:�@[����8`h��9�D|�<�G�R������N�\,f��$�_�DB�0�D(��0�1���Rd�1�2��(�
�=�q�5�j앨`X�A��oQ+d�*WV&��s��Z���Q'��-Y�C}8���Pj#E���2���eq�u)K���G�ʴ����~�3Ls��:���;%�3tW�S	EU��D���ĥ�'��Zapg&L�5��8��i�i�����b-Ru�9�E�#�;����#v�	���ؘ^ـ���ďu�^Yt�[���90�����Oq$}��M͕���"�N��WD�k
��X�!k�°�-g�'���Z�PK`z�'��>\B��p��:�����!.pm���K1*0��~���m�L�z&�*>��4���6�y�(��t@��k6-��.�
�>~,�΄�!'��@@v��ǐ��^ݷ����+G��وu�'B��b9%�j{��|�s=8�,<m�ȉ�_�of���q@��lf �'�h�S����vxCw٫Y�[a�J�6��>��������#�s`5�f7 Eވ�V^�h6a�4f�}�ȝ�q������9m�����x�O���wH�m���J�5�E�4�R�l�8��:*~��-:�'[�o�ss$G����4;���j ���{�W>��ue��z	��L~|i��Y��K�o�+�=̾��EZ՟V|.h��&���9X�YR�F�K�:�FIl6udb63X9p1D}�Qa���E���X�;2=�i�<�"���W;��Tu�|�!�LL����^�K+r�<@~��:v�G�U-S���o{�n�8��B�Q� 'S�* ��ÝJ�@�k&����5����>�0螂�"��Xrˊ�w�Xel~�HE�U�������b�R�u*H��=qw�/,\�cT�"�)��\���Ԛ�|qǵ�Q/N�A@�J�MM�_�D������1'	�~� ���L�ŏ�Ŀ�5���>��-H���,��{��VoV���p�׸��'� �{�C 9~V�E���[�?����ѓG��/x87��p��>�5����z�)d&�(qJժ�[�eo���H^���r}��bBr�\,K�u�na�1	�*��II%!�"��d��Uu�o^�c5������T�c��"�w�Hl-͝|��~$.���M�k���#7�r����kƩ�����=���mf�(��븻>�����=C�8�V�'���pTEբwdڵ��Ɣ��$�w����r��Y,؄�=�k�M�嫲w�$���l��w� ��Bt� ]��E��!��2���M��-��I�D���[5B�%P��7�}������e�z��>���%YٹTT�C0O2�����H��V"�eٕm�7��ǰ>��1�{I�.�ĐS��>˳ �䁂b�{�����n%B��C�
�|]�~�c���Qo���N�4������-4j�mT�|�Z��҃E=���դ_��Ur��y�bW�6+O0f�>��ӻb���KX�� ���&�����C�b&������)v.BZ�+��7�]�B����)u�Eu47�1�\T%�Ｊ�xμ�9�mvM�L��y�XA���G�q��{��v,���ɣu�z�"�M�$�T�<*B&���K�F -�+x��,�pɯ`J)թ���Jz5���Ñ�RG�X&0;�bA�mk9~Z��M�8sW���P;�D_>)$�M�q���D[�I]�Z��MI��5�C��*y�Rm4�HA7���t�f�:��|5s�K�R��#)[]��kDԟ�w0�mS�ɭ��,T^�����F�I��)�� 
���+�ڎ���_Z��L�l4&�D�!���6^z���T����M�E��əKM^��pe�F�	��u�����<��������T�M�l���\��oV�N�1���Ё(�����ޢ�z����)W?pg��PҦ���I�!�/R��+�Iv��1���,:E�gW��'*fRB�S�����$($M2���s�@��7a��Ԋ���@T����g�/��t�v�g����T�u�hk}Wq[ݟ~��B�I�Y�ٝ�^K�9$>x7-M��'�,ȯ��[ʀF��u�,��2�� )c62��9S�����X�2�z�`OYu�W�;F��ˬ��=vȸl�~�e�'}WM�����9������;-zI&�,�l�d��1X�K"�v��/r��D�ⴌ�$!�o����a�k㇂�O�������one��������u\ ]�c�*��~Nu����]�hk�pt	-|�V	�w��$�@�:gӌ,����*z���=4\F2��g�V~4�3p�R���_r� ��	���C���s����M ~8,&rY�n��ˮ�|Db��s8�(���m;�@����'�o��J�H���XsI@����#@��G��/�9^�x+����r��'��E�O@e�:����'���o�<�����/�")�mL�n{�<�\�O콢t{�X?Xލ�6f�%U]M��\�j��>�^���~tr��3�U�gw���:�λ�`ܧA����U!0.�;l�-�Vsi@�����*�P�jTi\�G5B�Xt�e�
�������l®Q�AR�5Sk,꼾���g-�v�r�-
���g��]f� *���"����!�վ8���o��U��nz7p�2=��`Y�މ�ݽ�p&����.�M ����ej�Y���*9"$V���"�E�^I9��NMKYC�E�?���o�`���#	`q����ZNB��6�jg3����	M�V4�hgZhø�UEA��y[O��_��Ḣw���Y^�>sL���i�����ې�R�]�r�,D����]�d��� g�]��8<�Z�]���:��L�:�Ȍkȯ	5� ���8Z���_;�3np7�!��� ]p�nT܎p}�Ð�F]y�Fmn$� ���pjA���^<����K�.��*�ʼdя<�tC����iɒ]���o=2
�)g�c�b.��(ܰ_�K�a�qr����O���9����#�eJ��}Ro�����T&؛��+� �~@+�G�E���ة��5�&���Ex~����8L�O��el�%k����v�JTP��*v��'����Z#��.�f�o�%�'0jgU^s��T�dojQ[gw�p	��B$ju���5F.;��or�Kg�@�n_ٻsl�3���T����/���˘�B�d� ���F�xG���.�� #[�[����1l\�s�yԷ�U��ɩ<O������T�E�mNY"�[�MAFVUZ+�B�dvLj�#i����p��ĝ݋CE����^υS��nؤ?���\�)*�V�V��D�2Z�a&y����S��'����������YŹ��i��L�b��O�/7�$���|�����d��c=�ScW�s�b�����#al4{��z*Cy�wSV8�x����H�6�=�����%�<թ/3)ft���Xuz�{f��*ch�Չ'�9h$�[��'��M����B�ɠ�+�0>��w��HJ���)1���~��IB��5�XY:@5�@�F\���c�A��.�U:�O]�zR2T��ug�ri=����!`�g�-�d��,#��``˧�VB����AG
���V��	#�9̹o+\�bNo��x�����<���pp��?ȟ��y)�z�VS,é�dc|6�z�5���@%��H��9�����A[$�Xm��r�*�G��s�o)�1ftës�����I����)�\�vI��Ʀ8���U�BH2n��+lzi����&��Ҟ_��=�zꨬ�����J)r�ݴ�՘T>�lbǮA��`n���f9r�};�ogO��,\�.e0[�n����G]�ǋ�G �0gq��5���%�ErRQ+��v���I���$\F��͐å�g���J&��#D�vb�И�5M��\��5��<���ÓF���p�(�>��.m�͜:����*z��1!��4�x��xXi�����6�;���J�ʃG�hA��xكM�>�s���i����&t
���a�V��u��s`@��^��4�jk鼭؏`��b�-��BZJ�=�7��(�k=���+x�<t՟a<B�!��I�h�6�`���x7������j�Q�9��������']���bZJG�)��+�)�&�� )E��Q�*�B�%pit�h#��b2C�[�B�V�2A2���S?Ph-p"�h	�`�Ͽ��>d��t"d��8��a0���Ɛ���oݾ"��a[�	)A�ËPI�.����n��p6�A�y}�����׉�6�٭.���NW�`�:%������]V%�lk\�fŶe�}�����PH*T�Z]�m��Ó?�-�2��챷����#���<�,�6t�������%�:�hU\`�~��{���Z"��2��5���4�PCJ�R���L��d��)*���F�������C6����N�y��b����yrk���O��<b��o�j�J�?Ntb�cn=c�@�ǑU�jF!���y��I#���+8��h=��b��.>6��zx0 �b%XA�ES�m\�y�tB��&��(Q�ʆ��*)�P�R�����&+~�`�4��@5��ǈ)W�#�p[���F����R��i<��Qm���7����Z]�v�BU+.��S��ɉ����6�Ր�z��q��n�(g��)WX�y'��C�,"o�JD�M�~޼#`�:� ��<%�>y2SF8�?�� ��M����9n��5a�c�:(#���X�by��:)�L:N��o�݌
��}F���n�f�����[�Օ d����H��Y��y�r���(�U�8�y�6��/e�����t���~b��gyY��E�QL$��T���ON�o:�9TdP����Yn�)���cB'Ӥ�e�E���m�O��빍;��ˇ�(�n��JY�5��b!=ЬΊ �a�qr�:��< ���1m��^�#.��v�l�p�`�ԋ,��.����w�L[G���d��hP}���f�G��0�y�~����
�q�p��?vª�18���P�i%�{o_	����u�q�yd�.�4G�-����©�0� m�U�,��ǈ����YN�$,�XV�c�@�]>��s�y�ƎY�� B>��O��[`�[e��aS�:��G�r����>"~㖶9�x�X�Y���F�	�L�����z�pc�A�gȓNZI��ł�C��?����oL*U4$_z?L�#��Q��Xq9�� 0%����#[NH��c !�C���2�@e����\ٙg������+��P�d��m�YW�|x���\��L�9��f���ЛG$�h�I�9^Q+#�����f��f�f�EC4��_�����Y}�YN��cF39:H�?�`#�4�ܐ`)���J�t��*&��p���6� S�]eǽ�C�cV�r�*��wd55�ĈPVQS�v��9�!���彍�����u"���ށ��'��0�3�x��l@��O�8�P�&6��d;�kt�����>��L�܀ޕ����/X�-��w���_�՛��?��O
���c=&�o��%N8��ְ������bx�rj` �'l��裈�ʐ�Ĉ�!4�1r?ۙ�*���Nb�>�������5x�>��q1��MϯE�k���~L���s�5�v�{������ΈZ^H��(����[�:Q�R$�$Ӡ��̹�S� �Ob�c��b���c�<�H5p6�q���>���ɅS�x�_^���d��??6�|�v���;�L'K�Jv�])�(Ӡ�1��sB�Bg��=F��ZX~������\e'R m6�up�'�Sj<'a�K׫�TQ�7��E��T�`i����G��ʹ��
�٩E**0df��w���cٸ��۫���L���O��X_�{��-����=�U�@����墫n)�wm��ĸ"|b�$���Vf��^�⯛�$	GG{�W�f��@�d`�<��n��;�##l2N�
��*^8����j�hG���0�` ܲ?�/�皳��̥��N�}��B_�� ���`�N�񚯌����0�_��9K�@�y�3I/��c\r�� ԫ��g��o�M?��i��f�7�#��6JX��ؔոI�*Ų<�6W��m��|S�4`Ϧ;׌@�v���v�L�jᆭ���Z.�}�F�?�ع��F�<e�r���ҷ-voh��!1Z��.Y����eI�[��(��Ƹ�f�/W\�U�� ��QȮYwn�kyRko�L��cx��(m��}
#, �7H�d�b�u�70vA��86 Ҟ���O
$7��0qJ&V`G�v��Y0/ʸ��pU?������ū��������O��m�F&W@~L*1�|�aꦀ����3*ov��
O���L�V��n�׵��`��ƌ����8c�t¡~0�J�O�{8��=G0P��k���e�0���i��ٷ�)�)D����܉"F���F[Ф�C$��v�$�!�zW�͌���G�~���g�}���ԃ$"5���m�c�_힨0C rb4@z��~�K7Ĵ�_qI��&��������r�0���*��r��+�E���c��O�9�r�)T*tn���y��-m�,�1��Ww�~0+���G�V9DR�c�=5������'8h�h��z0^R��QLUV�+���{�.4W���
�J��-%���e�'͗a�s�A�#ٴ��"�{?�_p��su��#�+�%m�~�䨌�\�]��b�H�8�� ���E���S�ռ:�(7x��$� ����c��>�r�.N��֗�1����gu�z>�Vu>՚��גF�	R@{X>ۑ�v�?�?���;�ƈ�Bf҆j*(Q^�^~+�b������&�謁�{o��>��Ќ�I�.:{L�	���%!���MW�@
����Hk����KY������������H����\��R�ص֕ƕJ1&�>�l�֮�{����$|�6۬M�j��e���A�^�t�·�����Лu�h�3��YS��舱��7�A�|[Y;~J�2^�L�����9�^K�\��Q0��*m}9wU���9�����M�B�ڷ=�k�o(�C}���;RIx5&�F�'���t\DݶpJ��]l3��{e4�ƻ�cү�B�b=�!!�o��o\����C����V�D5!��%�j�p�=k2�:��E/��O{ y�Ie���VD��d��YJk�uv�7V�w��&����h)�ۭAr�|�=pC��C�T-d��2Å���z�*c�0q�;@*���X���"|7Uyqm��h��6�v~)y�l�v)��$||���%N��Oa��E|\aV{A���w���Z<��7��'��Zye�?�勦/���0]L͟��}� �֢i�!{#�أO�$ꓸ}4��2z���jn֥��ey��\�mHӽ�z|uEl�d䂪�4!rυ��G�w'��0Q/e>䓂�&8����}�-���TޯN'� � A�P f/n5�� `\�\I%�_��N)f\� �$CMa��Q0U�$ӂG5wYr��Փȑ�&w�x8dO��g��<�r��a�۞^�*zf���"	�L1 S�vͶ뚗�.�=�
�&Q�0�����uD�����1�|fbƂ�{���dk��E���y=K��`���[­�����ms�N;{�'�a&-��C��k��_qK�u��)��K�$�#GLW�a����JA�M=�Lf�8��`N�R�;ko��W���4�_v�=�8��]$ �]�/�=-��f�ŖZ�#=��'�k �x��=z��3:ǜf��S{�ȿ:�ЉxCMw���CV
h@�����|�kh;��"l�6�t{�!"+���� ��׽�c�g���[���!n��?��u�����y�n_w, y�(��p�����l\-�5��cu��g1B�,�v���.��N;�V��4�Α�̍eI�R��K��� _>��+aaj��kV�i(��n��K]xV�agY_NU�Rb��R�����qgd1��.G��5G<�wh/_V@<��^��;�oR(���/B�tx�FK(�je~��Ҩ��8-�����U�� Գ�7;�?������t_Y���%ܖ��,�:�f�8'P(_�.��2����ܡ��2���iz�.qc,c���. !A�oU���ޛK�IX[�v��%��>�d�\�1����7�Cf�S�*'�T�g�,J/��������c���^U��`w3�%G�!����8˩�I�CZ^��l�l�}���1��\��&��߿�g}�JG�%�{������m=Y��:�[� @������j_\.-�а,��01�/�Q�a�^��Z�AY�<�@�S�Y�*��L]���5g���- 2S�T����<9a��,��u�Pm�!����37�~>��2�}XY�q�ѓƎ����(M��� Y�4�SQ��G���G��K��˸}�%�`��N����ς��1w��ԃ�m,>��naP��Tqm�q�Z�E�}��� �u�<'*mA��h��u������s�jQۅ˟����	P�y��9A�`���SR�����r� dK0QZ��;����~���o�rS�ʝ�e����_-+$i��T�y-@yz�Y8aG���=G{3�P,�W����G�g�h������[�n�ԤT  �fyU����Wu�� ��C4��$zG�MRzU`���e�bo��"�C���M��]��m��fDǏ^YW�X�R,,V_����|�ּ0
�H�e��(f�Ǵ�_xDyޣ�{%˅Uw�Q��Y���Eɠ卪����G��jrc}���f۷I ���g
A��2����ëVß�3gX*>Mf��@$B��y�c����_3!����[�~��/2�Ul�E�1�1v���jc?��.fG���U̮0�⎡��@\�s���g	+�}�x�ڤ�=6��]Um+)��Y�κ35������k!?\ �8ˇU��qqOK2~�Sc�۞؃���2����T����#�g�_��TW׶���xx�u�4�%�rڼ��G%-;�JC��߈ڤ�*�Ф�;��k�����)��GGE�oee�o�P=�p�x�?��&�>�η��!��Z��2<['��T��zjDwF��U��
���Ꜷ���*�)[��l���#�)pV\���A#}:C;�I�$1��]2�=�
H�NZ��-8�BrIsw�q5���S��H+���\Ro|r�3z.ܟEwn�b/�	���Sr�g��DN%�l���$j�,��o�'�i���fa��5�o(�$n������'��9�r��3�t~�� �����ﾸ\V��6G߫x���f�0y��߄[=�?�����Q�<�~)y~���K�5�8G8�u���:��F#��U�=�����~a�d�źFD��=Nl��9-��4klJ����3��f� g��	�i��qH�g�ɱS6&3}o�1��.}��q2�Y~��������%�&p3`u�y��zh��j+Bw"�)��"SW*L��U��$��X���~p��`_�1{��V�W���x�m��<�b��i[��Pg�oOL�y�ؾN�q4:͎�.~�Ku���|�$�R���r�ʔ�W֓X��Y�B��ϱw���6�;8�S�k�)&�N|7}2�a�����F.�l�qt�4�a򽺛hl/X��v��3�BH`d1�v�t�p���Q	�q?�5�+��h,~��'�n�iv��0
!����e��f"���N��	a����-s!�bٞ2�m��k@���̳�Ϟ��0�ɆP�A�A����F<�E��lIv4Ǭ�6�ƌ�\����l�ǘR08�'�M��Wޭh�$���]�(�7t�4�]��e�x} �"���}��v�*��4��`-�\�
Y��w����օ�����`���*�4+�}�f.}c�p&����4���}���NK�q:��֓a��~n�5���>;��}�f{g�����$1�f��I��F�g��|��Φ�~X�EB��gI�i�U�wb�R;]S��@��5��s7}�4��a���_�K9�Lզ�}	��%�%��>��!�-Y`AQOv���{������[��5�.��� 1�O�&��0<���u4��N�n'�W����'ʳns5՟��Ɔ�n�s��-A� �df�E�I�-��Y�j�h���Z-5��j�(�`%��A���i�Ϥ;	��}���n�Y\HG�Hr�y��;���ק��2̉O_h�[pA���+�5%_�A�|���+GҀn�&�j^`J��Z!L(����P�t'�����ء�!͆q�4'}"�ʶE��>p�&��^��s�łP���D?�|�T6E�C�C����\Gph{�=W*�c��ǁ`n� +�}2
N�%������WKJҳ'���)Y���O��3'�<(�`�F��$\��qm¬C0E]���]� �d�Q�6�: �4�ָ��R#t_3�/cS�n���Q��$��zx@m��ه1�>f`-�P`ʅFsu="{J�L
���Z��0>��*]�Odg�?��S$8]%�G$��å�<�U����������;-'m%V��{%L�l)ϣh6�嗳)����w|'�A����_왮�(��j�����k%�&�fT�9��I#�eS8kb�����.��z=y��*�-��<��+|W��纲94na!�д����>p��&*�,uCj����9o�~�y�ǝ7@�Ѫ,zQ+����p�T�&Cا�Q�2�5�!\u�4�22&�
ִ/��:3^��ܡ�[{]p��9|��i���4�S�@��y�V"����Ўf�J��(��xp�T��H��I��ڢ�D&�x���4��iQ ���d�~�|����Us,ʴ}����F��O�ޓ��B���	�>M�Eo�x8g~���{:�8#���P�E>P��^�$5t���n�?�G�[�8O �U$�8���3�1_����֕�kmC�>�o�Q�P]�G�Óc�k7@]��8���;T�B���/��MgZ^���3Ş,H-q�
G9��-_����,JR-��Q<��w�r:BNI��2C�h �G�y���֊�F����W1�L�2�Q�I�7�%j�N��:���H�m��o'qm,�Wi��\��^��tk*'��=~�~zg��$���Դt�w�ޗ��P-��b3�.����D
z��?]�s$nТ��Z�f	2��ϙ0�����X�7���^/��9�	M#�2�y	!dQ�b��=��/��P�`������7����E�����Դ+�+3$@�$�wmr#�m`�����J���&�\����L�Dv��3y�Kؚk��Ē(0���#���Ubx
�d�@czSl���#/��FZfb�q��&p�?��q�̎ i@���p.(�sQ�P����
?�{71���|O�*�!���'#1�ea����C����ey����㥚L�ϥ�C��wHk��;�x~�)�`M���wFZ�����"{����4E������L��<it�#� Q���jj;f�N�-Y�]�{-$ڛ����s�ݫ��E�g�"��3At�M�<��ߨ7�?����U�"�|0��M���0	�7yo��j���j�qZ	�MF*�8c!���8	�k_odݟ�Sp��γwH�&������?F!���.V/�H_���ق�{���ؿ���f}i�5�
y��}li5�"0�M��"e��J�_���);�!�ly���!V�yK�d����U�]����/x�b��A9���}��'(ȩ!��V�.��?��N���3^jٔs���=���"O��+���mv��T�(�Q.�5���w�00���V�W��y��É�9
��|h "bz	�Sm鿽�`"�'�⥏,�[T�r�v5K.��HᦸT]�����S��� �¿�o{7u����'�O��R���TDt���i�W?��CcX�HЧX�n���]����+�gF��1S M�mM��/]�J>�Y��l�^�{M����i��'�dS�W��[�I�1�9 >�� ������"@Ac1}}�B�`6D�8g�e_���[|�Y�j��1{�������l��W�8���h
�����~��Mc��0��@ob��/�P�YtM��*[�����ʎE�P+c��|�U.��l(��|��0�!��6��e�8jD�Ս�5y�Nc܂'��r/axH��:�����zp�����P�v�St���7A�Y@�it^��nߪ9")�$�j��f��zz,�Jq,H	���)�>]e���3Lp�tI��X�1��¢]>�
�Lw2ӥA�����v���>=�A��I�ͧ�ҳ�b6ETTK���a���z��sA�,�m+�Lrd��W�1(�� B�S�h��8k8s�૸�G���zK�Qq��>� W8!C{���$G7D�?@
?��_5Ҿ |~���C�\���pO�\M)��1I�ҭ�b\�E�1�M˨�@��:��'��u����'g���Ufa-��A=v��n���/�q�����! ��Mv`l��@-�և�R��a0;�� 52���@�y�nmU\#�O�:�䝳dʱ	��5@��n1}[� �@���,M3��h�}&%��y�B��3u�����{+L��u���~��b���V��!\*����Z�Wn���wH�S�ٵ�,��&��0&NgK5��IEp%UK��@�>����I4����E0���f�ޮo9��(�
�}�?3g��oG�=�J�#O�iZm;v�o�L��Ә{���@7�dPt4׌Z��� j���L���\��:� W��4��}�[(�~pD@����qɹ*��%\�\8��/V�?���k�(hH����I�<&J3���|�6Y�;��zں�O	��)�D;��!�f)6���P&�mVvRf��NR�I?�[��/�R��W�_	��2��셢��b��S�̥��O����x���e�W�˵�C�S���PH�SL��[��h����DI0����e4u�l���TN�P}%�\#����U�8^#��� ���I���_��9�������|3`K��S֯��G%��7��?WP�['��:�ŋ��c�P~
���8���(!�E~1��	Z�N������$��h�H�A�g>V���G�&j��';j�`LBw:��\;��~�ɘ�h� ]�k�.�=�\Tq��l�L��:Ϟ�V>{�0���rʗͿ;�-[�j7�P�������A�g�K�e��50�Gߢu��_�+�@,�2��Es�1���=&J� _���Ls����`��9�L
���Y�7�����pS����]D�}`�![}�袏=b�v��҆��$�r��"�/{ �z�OI�g.����G���:w�W�$U�}9�C�r閨��3ش���Q��w�O��DM/c�("_ѷ��o���Ě��wc8����kٴྜྷ *5�z��"hN��ݨ��"�/�lV���(��J������⭮�[��#����^C��6�4;6>�V�jQ��1��4i��R��9���U�9���3=�~6���*��o�B0��h�{��;�����B#���j8aF,d�~��vQ)S�ĔL%�ג�d�2V�_q!�{��-bU��k�/XA/�g��q�9���n����D�M�~���Q�&����k�n�Z�C��V�-�� w$�FV�Ux�S�tZKRP�t%��s��h>>����:��6]9�id2coQ��fe�T~�8��im�����r�)�r^6���+��w���@��2-5]�y�G+z����<�s�B�3W��"_� L�~+{d��f��I�
*H����L�A�'}%��:�r��sʟ�v���Q�<����g�c��	�;�Hb��|�iӞ�}י�Ҙ�'���HE�z+����Z5��j�����e$��Ǔ_�`\��ǯ��(�lE��X�9�Hv~4�%�v(�5{��ǌ4zPB'{�5[��Ƈ�r)^��wN	�����߲MaI��DMr��X@��V�>h�O��P�iw}Z�z%��`���3�رdT|�%nd ����8,��J[�̆��A�9���D`Zg2jО>�C��SqC�W���� T��z 2�n�%�*���b�����X����t�%�������І{�U!�K2���QKw0pT��h�Ol�;�@�C���HEg/G��j���!���a�����^�w��L�!�$�#�Xؔ�xӎl��G�Uյ��=���Q4��+��c�kr{E���˻���?J���~T��h���v��%;3�<�WӉ_|F0��?����rࠋFv7S��g��X$cu�զ���IWy��ӎ��%�*���]%�@���U�.�*=����P������e��5�8���%-#����B:/�=:�E���h�w��/�_ؔ���+_E���t{M��pWVx���mp2�d�?��� �����K����B�`�?�\�T�uG=X�Anθ��	}�������V5⟳"*:�q��]?���鷡CjM7�,�@X#����Ŵ�#АGyTq�]��F�!ru�7҈z�Z�������W�Y;tnP�X�,nS,�(�I����Hٻ�/��=(�R�7,r��@%m��Mܾ��mj�2�}�N��=�& G	!0)�ʚ[o0	%x\��,�r��ph��%q��f�8Vؘ)��(&8~kzXU��q~qVT�}-w�Į�˘�T��އAo�B5D��`y^���b���7E]���K��؞oYSz��#�Tُ��u\����`��9�}D�b$�ܓ�Lf]2�����F�xܗ�!��2��Z*�D_T���5u� (T��Y���|�L}47�d
��EF��O��5(V�ht����ݮ=�`�ɖt������σ�y]f$�E�QsBr�Ĳ���RD&;�����_N�0N���H�����,��t�W�`O$.���v�ITK͝w��Rw-�/���e��FZ/�QTvAY���z���"66�#�x��E�k�"��"*�Z%���Р_U���E�]��m�c��Q����~uV�ΨUe��FZs3B_]�AELs�0�����|�7c��74�픆#��l�Y�v�Y�KJ�y�/��,����aM�(��((z���8�9H#Ns�,Ϯ̳�nߏFk�ĝ�#���{V1�XA�!����*�zit�����g�`�k�^�?Z�ݫX,���m4S)طs�Õ~\q���%��x%M���d������ ��� @����J�m&V��U�����P���!E� x[SE	,�e�|3����J�=I�K���r�|
Ӡ��M�����b��h�؇ݨ����HG?!d��Qqκ)&�����ߒ�E�_�����L�����9Rn����V�5}$p����L�}����@K�lM_Is����7C9�pE�?�)N�ڕ�T�� �>����]]���m�Ƶ����S�jB),�s�	M�B��җ���k#U#R+>�!��=��N���L��(�j�k�Q���z_ʞ�ׇR��n�{AK�.p�6p�ܟJF>%�td����<��)V-��E9�n�PN��&[���S�4GF��]R�UD�7�9���=�濅P�-��[G�fp���Ťt5�7���f�2J� ��T��]��(�4�.�%�G,�ms�ĩ��A�B�@ܷ�x�2����@q6��;Q}�?��Vg� N(N�s�Mȱ<1 �&�����,rPf}9�rX�#�F�jjv�}���������&�04�%�=+�������ǁ3�^QhF2��!8A�2N�(����(I>S�� 1�(.�mhr�����2��2��Gq�߸c�V�W��(���]13�1����W��̔K�(���������Q=^&���gMY�0�	�E:Ț��o���7c��W�Q�RE�#O�(�Y��;DI�+�D6�=E�\==�������m[���*Z����c��{<ՄR�w�A5�{�:p�m�'{�.�ȿ��8Ou� �^u���P�c����mH�kw��ྜྷ�	H{"ϻ~��P��]k�d" �}*��\�+SJ��v!? ���|��8���0�n�gu'A�9 @Y2���LoӃ�	Y|�W���3��%���h���S��P ݖ�`�r��R��``F4�Ɲ��a��Z�d���r�fDU�K�e4fcV���P)���D!��������R��>�L8d���Z<)��cmv0�4�@�N��/\_nM�m"��W-d��qI�I���-�,r�QD��M��s��_Q\O^�<_������\���<��I���*cÑ�ǈ�2��hiφ��Q���4
�.��#�����Q<7�o��K�·�]�i~��QyOyl j����i1U����>E���D�ݚ�13��I����T)R�x�W9�ƕ�>��H2VN{̫��=J�5c'}`�}��id��f�S2��xC���W�i̱|�7��:J� i}d�+���^�W6j�`i�z<I �{g��tB��f��Qav?,�/nA�	�aO��l�3չo�d�RyC0O'��/#Uf���+�xX`��{/J���x7��?>��Lm,�� �d��u��	#�vSx&S�CutDcH�i�/[#��$��T��J� �3�$��!�N��"��,͍x�s�&=���[����Y���o�����[I9k)�^�[�hL/�ӄ+2�<߱��^���'s�U��FMD����|��?8D���X��Ĳui��{��b#Ҙ�'�������s5_�{�YbQv����c=���n���]����`��mU��|�a�g?%�Z0����yC6��9������C����Z�Nx�W�'�)�ZS�����IN��0M�X�*�&�o�X�ȷ�5f�й�G�DqwX������j�G:!Q�b��G˙�"��30����
�T��9d��z��ߕ�t��.�+�A\]7��U�F��$�{Y꫓�3O�6qk�;���Y�Zv�m_N���M]���ՙ�.�b�^���(�BE�`��*��tp^�]=v y�>dHZ^W��*rȹ
�����lEgϒ%*�U�z�A��m��u�w?�ʠ�/^����6[�[�+Ccb���EQ&��Q{�M;0n3Oy]R�H��JCE�~qQÝ��dJ3������g^HS�m��`��B-�]�Vq�L��ֱ���Z/���t4>p7�k���#v܈(�h��6�r�}�/�)��Q����*Z�����w�fC��Sʡ)��$���#��1�Y���n?oy�\h�n<�(�>��r��{�{�A��~ӛ��r�q����o����fz� �1ߏ�哅�x ��hLev�kx���~�wGy�ڕ�S0�A�_�O���{j䙉@��.GS�UT��z>������:dTT�4���D�\v}WcN!�����Ru� -��7
�[1rQ����"{�ۄ�p���g9bk���{`��8�$U�&/^��B��	�^T<�����ãa��@#�������/v�h>�{���[1%[F�S��	ۿ�ͫg������9�A�<�6��ķ����@��`[| Uȁvy͑�B��S|�_ά!\4�wh�S6�]ft�ւẔG$ ��A�2!����N;!�Ȥ���r�=�_�w�'T<���h& @O�,�1/3W��ڑ)��nfz�� :}[�n�ܙ��f���M#R��o�P.3 \?����UT�vFzUD\2�~=�)�����&a�P�e12�4N��_���!�3��pHةq6ױ�l,�}^�[/ݪ*��Wy5bz�Z���9s�4��rh�"����'/�?=8kNC�,Π��U`��vث�\6�F��JDy�Wp�z9�+U#q���]��
o ���[��{���\��P)3�uHi�ZU˅�2D1��E��t�s�vk�LRnqp5���\O�b����'n@G�����#��g�}@�K��NWl�	v<�"⦺5�X4��~�����t��d_n/F��ڗ���Hmç�FC7i������݀����3�C��D�ݩ7ے*�l�]�	���K �1��3�q���2%��5��C�=�E�L�$�x�>��98��ywpѨ���߲����8׶�|C��KN1�T����@i��9#)m]���Ꝡ_XkuJ'����	_Ɣm�`����A]Z�1Jd���ޖ MA��{�of�}��U�F'.!B�#x(�<f{5D`��v����؋�ڡ��?E�Bp	)��$���3oAm���P�$w���<������H&-8��f)6f�!��&��bC/w�D����6��3�$!��	=�U��$9~���b"�_'�� $��J�͎����ȳ�Kq�،R�A¸�Qdw�5WFYS���-��A�����F�2/V@�f]+�f�X��X�g�U������Q���{j�2�ob�!�2ЭAbtFL�#��s���ZF"��c��?����D���U��ː���I�DL&hR[�x�	;a���N�e�HӖq�&㖛s!I(��
g�נ������{�;C�G���jZC^P�%>���S�[0�؎���+���8O���C�I�k=���qB��!�d�@Ď��v�:�0��5�D٦:l.��B�D|=Ŋ;[�֢������,  �h,6W��2N�	�-���.��&��tw]�2M�UJ�]	��EI)OV��R�M�I\\&�j5�P�a�G,�l~�X��vG!���&A�rvf+��L����V`"C$h󰔣��}^�}c8�� kb����ǯ|�Xqv��TjK����XgT�F��mc��"��2��ʒV;�X�����0d��B,�Մ}��׳U㗒;]R��t����%�n0^�qԜ�	3�sx�.CLg�D�_�FX���T��٘�.ٓ�̔��n��-��&�D{Â׾M��F�E}V�����f~	��4���E_��On�zo(]��ۧ�}w�����L�;cs
>&���� |�Z�&�![���dO�:�/�\%r(�Kƿ<�@8r� ���'��)a�T��(V��&�H�\P���y����aA_B���ްfE���������r�a��C`*�,+��;gz���i�)4��,�OX����?ŷ7mƼR��o������'�Z��$��������M��[;[W�s=4����][ĵ�/� �V�ia��C+�:~'q�V���DKG_�1-T�KBMw�d%iF���n�т��e P�}�:� ���P\M�R}�$/sK�e�`\���K;Ŋ	:���Ey9G	햘$@�?c%��fw�b$_��{E�τOW
a<]a��,pqw7�ZZ��h
��c���{Җ�@��H.�hY�׊d�7X�8j�����hV+�/3�|�:~�Q� ,*��)�+~@P2f\N��uJV��8����kx�a &��b�i�yy�U���;�4E^�`1o��É���{U6�q�G�W��5N�����e��b3�͸��c��!��йf5�������[nS��iyGyH�M&���ko$e'��[*�F�$Q2�Y��&l�BMk�~0¹��@�b����$?�6%�g�4��o��	��*�ε�F!e��&^)��F� � ׯaԀ�_�oHAq���l�O�wV�3��5�σCϻH(��6�{�J�o�OL��A8�I�%��Z#�7�H0���LO_`� �ֆ8q&��qX���r�H�zs�$��&�]�*	�Ԋ��*zY;�;5��F�q��n؏¾j�����o����iO��(�$��?�����rymο�,O'��r�T�F�\�gm�.�q�OYg��g"_�����Q���SD{�*{e M�7�*�a&;��{}�MRĽ,�"1ˌh��mG�t�Wweq��'�9��~�,?s��o��+�P+'�F��>�}-�P1d=��1-��QHQ5Y:C� �?N�����TZ�.��:�a��F�d�u�[��l!'�f?��ed���$��~�v�\��֥����32��-˩p������@�F
_GT��c%�iOKs��^�i�|�$��E��\���oMa&oo��
_52^f�)N�O�7�uHG��m�"�sOt4�&�ag���D��a
��h�3X��fƞ�r�"t�Mm�J�#-40=�_t*��W��Ѓ��R�#q3������|��Vz��M���2*�ž�n�K�B`��)�E3�+�������M,�j����u�q3�
�Ү�D���7m��Y����z��Q\���AҒ���(�M!e�,��,/��S��R~��3����"La���s��LΈ��ɣ��U6I�U;�������W��U?���hX��5<�>b��g����U�G��xIm�C�6� P/��S^�,q�B`?�����ݲ�^��F�<#ڻ�b;
�1�{�R��zʍ���[�����(�{h�:(?'���*p�=�/���� �HX�mS2��ⶐ�����Ǳ���tZ]��d+o|�#�Ǘ-w���ڤ�"�������m������F[��o���:P�h}�_x����gT�U�Ql�و�=i\6c������[2wu툇�E|i?���o۶��.>�^��5�2˘Hu����T:p7��j���=�~�D�ѺE
���wd�.o�p`�=��өK�įۦ+	-QY��g
�S�k�ԂdFp[�)V�7�19s�y=& ����L��Wa�T��B/3��!׽�m�98�L��DL�A�[�{_j������e�wߌ%��\��P��xx2xt5hB-Om�z������ྃ�pUY�jH���&4�ە~����ZJ�=2f�O���֘$��i!��P����/�=�
0��:f�gM�����+�˧*Ө�~*R(�Z�ێ��٪)�������Ҏ
����T��M7�~K#�]���:�z��O<`�DĚ�yǼ�������q�e�Δ�}\�ɼ��2��@�����ۚ�٨���)�t�^�Z��6�����ANnM��`���a���"���t��e���~A%e���]���V��@��4Y= �{m_��3v<�w�f�f,�䀐n�-��%e$�~���JL����e� �����>��ԳL�Y�tm�6�0��PEUP4qYf�H����ɯr�b{p�gJ6���6q�����D;�s��Jj�n��ٰE�W����~�����������+�@�p+�R'��o5�R�/�ʦ�"\�O�mԇnr�!i�������:hp��Fl��m��el�\PO3���)=������~
?���:����YZ�l��Z���q;MZH��q��f2�mx�l��a�4�7l=Ld�}��<+�zHY�ȩ������ 'i��9=S,TNm�=ۯ���t~�X��J/}���	���"V5�}�z�gqط�8�"��&E�����޽�㐖[�?���?i_&W�9j(�y���(��I ��Qu��;U^���:/��@���H+�F��ǏF��Z��+[���{�S^�7�s�D���%�O��,=�"�����GŴ<��v�>�6�v3��&ܢ���W�z�U�����ƺ���n�M#V��).���q��-c�{���kLP[�_�i���NI�>�E�x鎋nςP�5i�R�q"/�����`����K7糩����Cױ�f����+ׂX��T�8�
�0�_ [Q�=`6�#w��O-�]��Sոf!�h���5�G�>Q�G���2|Ȼ���WU��!a�m������n��N����:�`-`4�u� ��Tq��si��m@aVи8��t���{h��N��D��KU�< ����i_=�ϧ�w��*�w
�ږj[r�'s��BU��Yw?@ߗ}�����2x"h�~:�Wk^�0�w0�)�z���s�2�U�n*=�o/���:pw��������u�\�u�M�X�5Vx�5@�WN?b�Iي�T�-$]jd�(���Il�o���/ {��g}�є���s[/���ΟޓÇ�5�R_7�z�?�3��7AӬ{:lk���D�Qr,�1mfq�Ƥ�t��u,��%�h�g�s,]�t�͊\�#����Z��u�I
\������×-�=G�Iu��p0g�=�Gpj�p?d��R�+~����o����z$\Os6�`3�<MQ ��Tg��ZL[��޶�	,�ow:m|y������SmR|C(��1�M�� �!~	g-��vKC�6А+�h7qO�zV�ۗ�d�{��'����H���e�`��
����;�Xuq�Z��4v�ǚ�P�s��Z�;�l;ǋ����Ęn�ze�QxɟP�n
���|�p�q�U|���!q�R��A�1�	UО/��)F|�C�|��60��I�r�ꥥnHQ�7QF��;ewm�.��N�y`��'�o!+��y>#�BI�N���m�!�!Р�61�Z+�F-�2%@�ċ����n|��X{y�M���`�!�}Ӌ�	���.2)X�ٵ��;G��7�?�c��'9;�d�!X��@�um��OZ?��Xb�^՘�m�������K���*f�1��S�D��k�	"�\�d�a�*����\ �5*�S�P4�DSb�����E��c�� 4UU�%�X�IM�!+ҧ��Ohv���%��܆Dzc���	��٣��7�C�bCB��n��܌xv���M��[��q�R���f6�Q퐏�o�aE�����S�0:�@w�e��Ey�GS;nf�� �mϘ/�2e�J�~Y��_a%`��2�KAc�*ozi$8��6�?�X �u@*�Y�n��o��uVTK����Ĺ��)�4�JzO�LT���l�kJ�GN��y�h$�	��x���� 0:Ѓ�q��3�$��t7W>�R�A�����4:��rD����]@�r���NPhU�)��%(�}V�APHM�y�ԝi]R��4�Y}��h�i�#o�o�Q}�J���M��?��:��&�c���T��p���GD$E�L(q�Q���,�xbBvl��|~��ʪg/����6��G\���F��?�����e>��F�����\� �'o���L�br�!E��В,��?�-��U��5?����l��kɮ5��VOF����K�+� &D������Vq��ǔ=-���N��zD�RVk���D���U��!vk�G���X]N���&<e����U��P��8�N&	� �.���ܖHO�NX�Z�n�W�+�p��������G>{D&F�9���C��<Nؤi��/��T&yy'M�X]XB������ڮ�n��!&ʉ��X'���y��
�X��iO1��Ӗn���he��4.��#��$ m��S�2���ps1\���B-L����]xjX�$Ӈ�끩5�/�E�2'g�J���?��nrfQJMO��ˉ�@F�e�gIx�Ь�<�4 ���e�"����F��64[n�vZ�!�
��Ne �1�2q�B~��A4~��dxF�8�����|[B����
�K���UTJr��𚥙?�?�N�2�4��)zZ#wݷ4]f�����H�}�ok��s�TD��M���Џ��AV�l�&��k%M\���P[|���Ԙl��2U�׌	ko4��/�M�}j�K�i��Vu����i�!-;�_�6{��c=ܠd����W��zm��|�8�la��W�<���E�<+�����ϱ�*���ߐ�r�S	���ݱ	s���l��փ�>��C���CG
6T�Q�T�.[���/����~mU�]��c����Se)��ĚsI	�(,�^V=%NW�ܺ�3��#��'5���E(k9r�)TTF���(�?ʢB��ʯ�^-��̦�`�cK��4j+eg�mB:�J�5S���t����'��wIi�����'�e�@���Ƭ�D��#i>��u~N��}�R��_�,�o�Y�t�{��Zn�YC�,zϮ�k@�֝��e6q���l%���J���f�[�e��`�gh!DXMW�3U0.<�{��CټKoՃBu|'�8�4M���i��,@�g]_FqF�]����D��I�ɏ]�[��)k��X�|̸3���
^Z�7�I`2����L������$�e�G_z��O)9t�C��&�j�8�����-8h��̱KY�dX]�Y�+4��m%����@q)�o�#V? ;R��V3����
^h;�4D��v6\E�7	�ȏ۬Q���\��"~{�,3Z�����ν��6F����3���>�E�g�����Ϝ<%߹|�`��[��/��ڠ.K����ό'TF^�b
r3�4�z���%��o[*	�[��>)���x`k,D19]u"�ܧ�ф{�就;4G�;���B�	��<�$qs�
�UBrcOqM�V���o����	6�!A�
9THa.=��I��B�"�t%���@��ꕸ!'6/��&�)�������E��++̚���!��߆��g�t�2�NS���� ����;k{C�Q;�VXƶ�H|Ԅš.$���/���;%����G�����S�s��S��۞U'2��Q���
� @u��(���$8z)b�o���ٳ�$Z:�*u�Xi.���|��o?}!�M�*�+?���޾��j�-��4�~�`7Jz��!��l{�C���읞A�H��;?P���GV4�i�RX%by���Hfv��,%��K�ע�^c����.�%S���S�ʽG&E�v����(�dF'{��A��9w�����Ƭ��8MS�pa�R��^T�ߩ+ޕQ��N��N`���బ8f|}�sx$)�AϿ˕S�βDQ>�K*噅�2 ��uHg�A'Z�LAw/�F���)�Y�����q4���O�L|��+��c�~�/��X8��{�V �ɭ���)
�n�K.�F�[�ϟG<�Te
�0���WIh�Kt�Ǔ����`�[����Ջˀ��0�*E��N��ސ�xq��^E�P�\�}�EdL�E0:;�kɏ��ي��I�9������x����4k�G�#V�2Lׂ�ٵ]�hn���S�7p+y	5��Kک�8�xV@���t�7�Dڳ=���T�}��b���E^W1����c;�\���D�M�TЫ��GFn�T9�;3r���6�;"	>@�x�s��2�"O�.+	n�uu��Wl�l�Dlg��K�F���пõq�NT��@��8&�}���vQ��¨�X��(��W<��@mP9�c&[9�P���z��\�׾�����g�19�9ܟ�1�gιV�����@�5��ѻ00ƦnP��4rВ\Z�MǻO:`6|O)�@u�=���T*�r�� � ����R1̶6(٠��u�J(Ѣ?�00��S�;�
R0즇k� ���ļ2���<���`^� \G K\�t�G&d.w�
����vY��;�l$�贽fG���P�W�7���~$͘�Q6�J`�N�D���L�xZ/�+ː֜vf��:�.eI��w��
IJFV��A�K#M ��IB�")��o�@_r+�1�Gy���|Fc�/;��Z�ĢX8& Z'���P~w�0��G ���T�ˈ�d�*ä���s��*axD�7�|_����v�,i����T��B�ޣ(@�����#����>u���(xڟ ��k��>)˼�U$xy�#Z�i�c���׷�]X��<�^�N�ȸ`�}7��iz�G �oĝk�=h���k+�=�am�����M�_�f��r8���ْGv*]
w�`a�}��y	=�5Β/OЄ� �T�����#�w9-�C�P��s���`�j�ZΧ�{�C�Y5����A v�!^0�'�T�)��j8�aqre�5wVN��*t��x�Xp�Q���CӉ#�r���,�[����I1O'UJGD٨|q��&E�$^�f��\L9�b1�\	�W0�+����ٞH�k���U�y���`�f4�r�΁Zg%9��8�W�s���|V!o�J,�]/�%3�3��Qpn�0�1}���4�ړ�]]���������զ��7bL��p%�n����F0R�k^����ˇ�Z�8d��T��"�� x�� 7t�3;�S�͛��4�\jNq�x�o�(]-\��K����'�����Y����5��n���C|�uH�W�J�H���	ɀ�n��'��{�kB�TǦ���Ӫ^eh-�7�n�{w���[��IJ���`9c��t��$vn�48��Xr�+ѵ+���U�gJ������ �5����h�%߽�-:m	��Y]�ld��RMP�|[5��~?߮t�Ll[�\�7��7�;���Ct
o��]*����OW���HLV8��R�b�T��¢_l3��Qh�IOCmA��E#)뜔�c��Eig�S"��q��@��X_��Z�g�ު�"a�܃����ɿ�l���d�cI�� �S<ol����s�<Y��J���x�1��2v��W���y8,\w���l�.Yb�`z������C*���u�* ���~�|p��-��M���+k9��r�iUJ��,E�MC���G�b�!�_�g�x�:�����\�r�b�_�T�c���n�EX$�A|&Y;m�	��� �8q.?�ղOt�:���p#�w�����8��"*��V����@�����t�v�WQ�o�\�/��ݲ��B_����]{����H�\T�$�GR����R�,إ����ǋ�&�+c��<վI*�+7��۽d% {T)q:�{@��;����3���O���`)j
���������{�[�[�Y;áf5��(v�W�I�A���y}rr��ͬl�h{-��o8>�⺘���JQ{T���'
������@=�Fnk%a �.!��o�|��p��m�/|�xn��͵0P����r͌Ԑn�g\V�@7_�`WO�`[i���+H޺R���G;����N�ᚿ������D�z�| P�8���x���$���y'�Z�>�!|X���_��f�gQtx<U(w��P��?8{���^�D��#�*1�z��D�0�N�n݆��K���O�LI��7��`v����f��.��
w�O��V�S4ԭ�"u`�@K=�L�d�8L�c�(�T�wRq�}��@�lW	& �ݡ���$O��$G�2����H!U�Ჳp�p��	(8N����+<yĉ�{p��8�e
OX:�W����N�ve ����fߣ1��`<ӛ�"J'!�6
muhz����^ѻ��e��t�v n�g(�,f:F���4W`�}��ϹQL�3S˦#�VӔ�Rs�V��w�^/LY��=;U*�ܱ��u�@6*�44�(ݩ#��6֏��ZWMMQ�>aO�<������	���#���8��6f�t
-2��:��a����n�y�S��Փz�-^�~�h2���N�>5�y��"�o'��j����U������+P�Y�d˅��Ț����3��	���4��ƽݱ�[�Z2'k
���D��M��/0�첿$qr��W�j>��"2�[�}�$�>S��4^���F��ݟN��Y���q�A"�{͕}�%(�0 ��D�8gƢF�k�{�6��8#oZfL9ˍ�|Q!�4��Z!�$�o5ǟ��3yd!J^�րC�ܮ������Nxeh�Ӗ(՛�8Y[���}q�[��0$��D�_����A=n�{9O� `��F����+��Z���s�4#9���y�Vk��,G�F�C�[��l�_4��~�,��E7�qb]�^���˸;���=*}��Vq�tmy���"��g+C��b��Oz��8��D�Z������$�e��J^���j^��a�[N �o�l�C�����c��΃KK�߉z�F(�_��\*2M��E��	���o����;(E�m�ʎ/L'�ז��^@�Eט9f�x�H�X�*�+fYCW�f���E@DT�g��nTc/?!�Z���n����ˣ��I��6DPy�rk�XA+��la��-��d^m��b)s�%Cwʧ�fw�\��I�C6����������A  �}I�/��E������a�ľ���i����C`��\A���Sw�;��.������.�y�����GU�2�g�3��o���E�A��`��y�yd����"����hc ����L�:�ȥ��	ݠHt�o�B|���	�	�_��_�l��$�N��@-L d�\�/�8�o��3R�E��t3-x��55~�ڹ䝖������>����+w�~���
0'���T�ρ��F�?޸.��֪r4b���PTx�����7���w�r1�Vl#����@��Ue��1c�Z�mM�0	�/�߀�h<�(}ۓ[̬F\�S�����oO��D�:8�&�K�f���8�x���8��≾� 7�NOHc�����R�p?sW�r�\ػ��i��n��o����ڍNݮ>�Q��Y4��1dV��N���ڝI�k���5J����`���*��C�p
�Os�������1q�Z��gh��ӟ?�)�<	
�)q���Ҥs�P=�*^a`	����{�zʈ.��@���u�e��a�|`��/�����K�|CP�����j�&$w��5Pu΍0��=��"��w�bSr!����7�^��.ύOQ��lo%1N��t������{2��g�n�_2����HQ�S~�\(� ����0��^k��>�l5ރC�ʏ2�� �[m����O���!��ڽ����G��̫HBN�Ҩ	>�	ȸ�A��zK���H�EY�l��:��z��'�.�;W\�Ò{A��p��.j����(�Leұ�Z��޿Ӝ|aί��z;����ܘ-d�$���<��ə_q3�\�f�u�O�������4��7����#cqR
�zi�y�	�k�Uӏbڒ��|Ո��՜t��%��T9p��V`�����#?J)��D���-��g����N|ڛ7�ֺ�Po�}L�z��ne��]������= (>��O����C�PWXwT��D�|eFe��k�6�p�y�W/*#���t�mrK ��j�D�wB�bWO�~`�.���V�f�X]���S�^����'��l�L�j�f���~���f{:������^�^�B*9_�"��]
_��of���j�_��������8ݹ�%���M�'��u����}��5�|�d�n�]�pʺ�����5�3��0���h���"HǼ���?�K��G������a� �'X��&�ey�s�;�=����N=v�H4���(����gS^'c��f�2��S�q��Vy���}Y[�8�=��t+X�Y�X�em����M�7������s��z6ɱ�}w.������ne��4g�Jit�i*��n�w	��v��xy�蘅�iU���(�p��Iۉg�&w��~l���.���y$��\�']��#g��TYK��le8'\� �
't��87�G��e�z��TTN߹ <�Ѱ����L;j	���\߿(�SC�K�..�Ȱ��ou%���(����S/��w���k� Д��E�3*�-���D*D;>��}�j������'MEwKO�z��|��,�����f��t%���gĆ��Ml��K��a@ʺ/������6��Q��b���J����������h���s���M��1��u��Q~"�!eH��"`G��,Ґf���-~�t1�S�I��wQDy����5�E�,�kw�l��wJ_ta��"���Z��pƠ�@_��Z�V�S�V^�n���ؼf��o;�iz5��Zpy=����zRS�%�0�0i�ak @���%�n��BxxF 7��{����\�r�q�XDR�R�i�8,86���Q�쓉+M���+�1#����l��kP��	��p�����>���gƼ[n��Ц?I�����j�,�W ��#��\�2$�Qݛ�4Et+t����p����e�L���+��J��٘Dew :�X�/�p3�)����B�����TBM�g���k��>j��*��|�+5�u��i�Xg�Y��e� �����Ҙn�"�EŴ������ٺ,a��\٬�;UO�È�ZOȬ2�gU{��t��/2�*�tz���U$p��~�L�9�w����}X�k�a� O:��A����n�N�WϷY/w�S�M)N�sE�'�u�|l�B���/��d�`Zn<qrIE�3��1�iu
9��E����� #G7�0�mJ|���_�
�=�X�,^���T�i����]B���ba��$�[�Q��͟G���I�@h�T��@g�Nk;Z�R��`N���ֲs=I�f���r��A3�S��/l�����ꔐ�.����N,܀�@��UY{�H7�g0�lZJZp��������tԅ��m��p�����u"�c8?e}�$�8*0��W�0�Z)�8o��.L�t��KL;�X7wKv�ռ�ւ�ӹ��C��BႪ@����>�����~Wv�B�R?��uL</���� L����Q��2bU�����m�<NNeE���@,�E^��=����*��C��4Bl�	E,87���zDWtB��o
f��Ѧad�:5+H<���Ε� GG�v,�X0�c�{<cO�O��sq�gR�D��
&��ih�&(IC����\E�
�U���!��=#�q���к�B�q��Wy����E�`�~���7K<h�QAw��>�*�C�@�(���L*&<�3d��K�2�1E����!	qKaJ��Զ�93(jtգ8�ZuF��,����UmRBc6#�7�
�6�3�^�%���?��8!�>��9���E�Y��b껁�56b��BAQ� �����E�u�'`R�A�C�TK�`/���p�u�@�-��'ΐ����*_��"+���DcG߿�M��@��忠5�$���c9C�}k��f5�y.I��Z��a�;o���g��������3��8x�/�`8�}����+q���I$߯�ƞ�������(����o:���p�ى8�PkW{��;��\haE"�,j������.��hD��:���:/&�7�ǟᯚ������jc �/�������w��>�"�t3��Ttڳ\8�3��K0a����h�bJ�=�xlx|_O�k�����?I�;ȉ����@�����GW�}g��&�pFɔU���dz�i*��=@>�2�oLi1	Ь���س�;��O�)^���0�%6�Q'n��;AW�/��fQ7�|h�{!�&@�/n�2;�_�8���q@�����eR؉�8����z����k{'Y|�Tk]��L3�$��+S�J�l!�|p�7̯�'��'Ϟ�wdq����A�`F�[\~��~ �hY:T����j�Ȓ5$�������Ȼ�epn���e�ػ1���u N%�����&Auݤ_�m�����U ����D�G�d����ݓ<,9� ��u�kGI��f�Y>t�iM��h_z_x��D����	�j	���'t�t�[�����AOkT�#bd��T�=��K2��]F�jaep���;��94��4nѠ(|N���:��4�/��fFIKq<�c���+�� �YR�	X�y�:7~1x��-�RQ��悩vfڜ�����2"�q?�ޝ�A#�@�P�e��+�F�r�Ȫ���^X�
;|f�?�J�V�}W,�ݲ�G؁^WJ>�8&�ŀ�Bw�!�+�jkS�Yc��PA�����ZT[�d� ���-,Џ&�,� ��|��¶0H��g际�#x�Mv:k\������;K��*��C���;�mm�P�27���T����:�A`v;{���Rz~����ǟ.��.s~��hQGQ��t]p���x%�U�%�*@���*>Öo�Uѿ�ѡv<�+�g�Y��������E�Tt�d�[s��~�f��u�?$$�g	V5���0Wɠa���A����5س���B�i�?(�e��ϯM*!!�/x�mH*�'� (1���`�Lw�C[b��Z@�'�����"�ٮ0���Mj!f�mυ��q�~��?Ea2����ae����du$*���f�U�h,nk�Oh��bWқ�x���*�Ts$�32,��Qͻ��'C��W�b6 �����-��-_���|s�Y�9]5��o���>�/8'{rc��lSzn�o�U�6���և�鍜 T�G�0zkT*9,p��=��(��-�)�	;����sj����vц��=�9ȤP(3��[�$���А8��x0�QW���*SD!�s��b�*�~T���kUb4�_!�U�P TqH��8���~�	��̳��ܪf�7Yuk�"Nwi)��P�����x������7�IE&p�h�-W����\D�ɼ�!�#�}�5�L.�`��T��&
 ��=�3^��d,��?U�f�[�n�=	p���o���[j���c�"i����|�S��[o�����E3�C��)�ՄQ4����夨�P�C4:1Ꮄ��?�5Շ]Į�cvCg�bN��|�,(U+~���g�b�]D���G\��(���#E�x�o�UE��e��n�����6j�A���Y� �!��)v"���C~RSa`����H�]�0|��g�HU$����/N��Я�P�����/a��@��ݿ�k'�Y)�W���NnK��!q�j�nb������ݘ���4mH�G��=0(�2��=.������3�SL��������ې��;M�ř�_�'�J.y5"���K�
-1�78��u�|��|��_Ў�-��T�p[ɜ#�~3�,�5�h�S��2��&����+[�4ϑ��])v<�>lY�	��Q��菭��8���=K263�<����Ѱa�=��,��O��#�Ӎ{���͏F3�WH��Q�H��V����a'L���gi��=�9����bG99+s*:�)6���}7ZAN��-�"���ph�ӝ��>�8�3���p+�a:�.h�k��^q��K�L^�.o2�ހ�7{ߘ��ԆC5'z鮂�"L\�噰�"r&^� �A;wq�,o|���:mnJ�3�^ �Jk��&-]��ћC��-�
���*~����2+ VG�n��u �T��J�� 1q?F4U����^����8w���p��On�Z ��NT�β��x�i3���S ��&��@���ä�K�Kl�#�;��J�}V���%Rc5Ahdl.�[y|_���ѿ��1�5�m�'B�	 Q&k�Bu*�ag��Nݶ�ϡ=�{K+cOC��O���D��?��=#��dK���f�������+_Zd��&�Μ��3_�Y��kp�X����6D����.�S��1�`��fv-[c��U:\_1xZ�?Y]�n� �h�ċ�)PT����r�y�ĉ����"vlB2`X޺��FM�c7����]�ǂ���#s(�,v��BL�`��7L=~��Qv� vu�@�"�Wh��V�$��3������ܼ�|
�)�Cɏ�GB&K�u���z��鲖���s��\�Lj#N\�@f^���^!�K��[�;\N�<~�`�d��6yGH��-�1x*���䮅�Vzk::̇Ӟ����=݅~�o'L&�W4����/��E�j��=m��T�N�v��!Lz����~��E����-���1Ϗ x+ ���LJ[�L`����<8���DM!^2d� * ��u�X�<�x��?�<�%�=D`��d4/�P�O[4�O�-i��	$��Oիy�΍�R8O>L���ɳ���Qim@?����Ɂs��c�؟��`��f#�Ǟi�V^'N[pEM��Y��t�Qկ˚�
1))=��@<�u��O$[�h�bF�,�|��^m@����h����0�|�'��p���N�ۯ�(z��MB���JV�V7z~�����6�'L�Cu�hB2f���Xa}}�Ƌ�#�}���J�;K��N���������2�'��i�bL�OS��`�"��sR���Z�R:�8���Q!�6�4��C{�k���U=�b�#+����.�Hz���(�)���q:��{����흡�%$*O��n����e#r5%n_�T�/�N��'�|5\-�R-4�;"V�i���l��2O���#����(��T���<���,���D��uh�3J$,i��ґX7�	Pd2��	���?�ܮBDP-������f��8�����Ƕ���WA��(`�K�~=�� �oN�C˺��O��&������'<��*��P�#�2�,1��^F7ǵ�Z�W����:��Z�T��O� ���c]ћ9�\f�~�x�w��G�`e�q����}���4���<[B?���UF��{�t�Ӎ�3$��D�Z�:��"���tn�nE�c�n�5s[jl�٭�W��%U[��t.�'Ɲ�"���*}/rf#�j=E_���3�1�4Ҕ�����ɼ_Ĕ#��r.�?��N�`�ӂ����C�:zf��X>V�u����O�� ��<���A;#8rQw��r���ޗ������H]�����!� �l0�~����2���һ{A&H����"�}z�W����09*[k���|��(�ϧ
�@���GZ|�"i��]�]0���ss���t;�_�e ��Gk�����K�� �Ag���
O����sm3�A�CMH��9G�}ضI�s̬$K��OA.���N���6��Xd�����*R���XXǮ[,�C�al��.(i��;]M�՚�/�V��ȶ��:f��/�����0|۹ӌ�8��ޥ�؏��)`�9�`�����3&�m�S~0���iP�{�н�����rex����@B�?ğQ#�j�hrO"+�A�t�6JB.�e��{��I�����u��f��k����V�t�4q}A�iC��}�@�*�>2K,, 3sR���\Q�[�"�«�!F _s�K'��bv�c%9���kBGE��Ñ:��<�υ<�ép3�en�Sث�P�[�3��$�;adD��a�/��fGI�:�e6:L_oVmd%Ix%�>jLx��s莐�\�(�@���AW�ļC�Y������d=g����Ͽ"-��D/h�	WO`���.xr^i1��)����<O�ũK�u���^m�j����ٿ4h�׹jm~�����5˞5�A�����A�p����`C����	XW�h�vZ�]Υ�2��D��s`�1K�M4�7'�u�T��.�:�>�,�f5�;r06t��9��c��� �a����ߒ�lv��YVV�� A�gw+��P2�7F�ҽ"(�e�Bw���9��A�d�2`�Rb�?�f�g�W���e3sA\��2 ��,:Ñ.��q;��C"\Wv&�M@x���v)�5�!\O�  �[��Y����H;� %�L����C,M��7�+��Qi�>�tZ��	~�!�k�y��+����%�$?Љeu��j�����w�N��F�%�6kG�l0�/�39!�X]k؂J���d�dy�Wjw����,��j1�c���Y�u�S(��iT<晽nXad"�&������|nv�cN� b���f,���(b񀇤>*�R�2�dNR%�� �-]��0�H�9�;z%�!�R0Xl�%�ҷ� D�ӆ�l�QX M5��M�+�R���8,�w�Y�_L�'�鎈Q�7�Ĥ+���>N��پ�S0�gb�~m�������T�Ո:E&��n�9�� Ի��
%��=����g	w�:�URT��Q�o(��.E��8�=�?l����� �R곎=�3�4����8���nF?��̟B��)���]C��f��_pTFܻ��D���E���`���^���&�������UH��,z��_��oHji��PJ+t�L�DIW]�I�6�H�0)�'��}�+CxN�K�?b�@x��F!�Mc�(	b ���=���^��6�?�nP��YeN��oJ(d��`J��U�����o�<Μ���Ӛ�)�0E<?x�&vbY��2�4�߁�U��{S�Wǻ�*�}�qB(2Q��d��Wz��C/5�.��w$�:�(PH���-�_I|�mL�{e�-Z
�GT��`Q�0z��5�q����t������G��vt��J$��'-`K[�6t����W߮m�-AId�4ސ1g$��M�Z⺠d��k���mÂg!����q�֞r1�|T�|�Qi�gS���%HM8��}ѓ��ͼ�e��[�����K��0Wٶ�g��v����ʗ���jh�Ӭ2 ��m0k=�r���&e�FQ��|l���+���jw�A��� "�a`)Yl�ލ�Q e �ln�P�Z't:
�-�_{�s�$���'�tд"�f�c��dmn0����i1�m�j"hT��-�X�c��B<z�:��2���փ�Ǹ[,Ą(q
���D�qB����↘v�]�F�란����t��G��T�/ZR�hQP��6$&,*(��{�l��O~/l�Bܫ{��\���3m�� sӔ���JdH%�~���g��� dn8ݔ�eo�DE��%�6n�˦W�z+̷��zB��2���� փ�q��f�x>V��n�����%�g	&���X�R�U�y|@\�i�z��&P�	���C�\��r���:�<�L�-m�'�~� �ap|iH>i��U�@b����ɛsn�&컕\=`��E��֜�7B~v��H,'��G�b�h��gZ�ۼ���R؁�G�R��sF����0���)��p凧�؝����;�wo5�	h�O��F�㭌.��1x�MȈ���^q2Ư��6��%nϦ�$m�WP����W�Y5�y�ct@Ŕ�����W�C9�t"t�J3�G���/Km�����k`�$��=���,õ'\k���.S}�y~J���tydq������f2�P6Yܰo����Q�Г�@�D�~n>��G��s�14�H�9������A��N�ĖW����1okM��I��qOt�1�(�n-ǀ�Cxnd��O弔1�5Cp�h���0Ń����r&_�2�	�G���X�im�4g�>�����q��B5@w�>GG;�h��\�ϩ�*�j���b��=�L��̊���֯Tv�Ox[N��=o.��$��!Aq*͋��*X�1-��Uf�F�@0b�xm�2U�t84h�Ȇz��u�?����N|:.��	��M}��1�(�*�6\�?"B��
.]�	,�8(�##v�xT`q��l1B�wAj�c�AW�^�O����δq�\����J)��/�t:p�������ZE��]�J��B���K�7��VȦ�f�t�Z��}}����u�+��a��g�]�-�����-]選���B[��|�:������TNɮ��c��Ii�(����!�)e�hBQ�:"��}Z�����}�/�j5�m%@���s�T85�g2��T��tޭ�K�w�\�"���*پ����VSde}�@�,zQp=�}Y!�#^��:c��$�be�:�*Qa��o�\��ú*g��&�D����@�͊�7н��.b��_��/���DAM�q��}:�Pf��`xY���:�7W��8�Œ�h=��v����C:�_rFT@�=���%$��s���1˧���%uFl�.
0�]J�va� �����V��T�ۃx��4��N�| �m���`+��=8fͮp�v��։t��J>�;-2�Iz�_Ã�孛�*l6`�9�]Q/�q$8��~����U���*@�bj�4�}&_K6�棋���br���$�[�����`��kO4����Rq}�lN�V��������p䌱�Q��J�<����yf�>g;xiKD�e����2�Wv0E�aʿp�K��l��T��@4���x��t�̎�(�.�vc���
H�9�)�͗�8������MJ���<Nt�b�%����P����2o�Q�chևv���5����9��Wߧ�` %FË�ڀ�U��>1�A"c�.`�+�E|P�M]x�$�<����
`��������� ��Ox%GNË\���B1KBt� �>m~��p�C�9�|�O�,'A�b(c�H��H-F���n>�B,�e�u��Y�ْ5�q���v�����X�k#��Ћ��[3:�˝Z�`� o�:Xxd�����q�$w�SǊIL��c�������jM,�CDǰlc(k�$�*`���^޲�L�f����ڪ��r̋�\�1U��fn�ȰǺ5�ۻ\b@�|e�Ʀ�X]1K^��%��]D�7��,��F���s��bWɯ��y�Fve�<�����t���4����m��HX�"���������96�'e�ϫ���tW��)���8���X�w��bª�V��� �#Rv���<4�G�{u:�t���j�	*����M$�I���w5�gW+�q MW��Z�#��*@��bF_\5���2i�(�!g ���=������R	�����(p<��r_d��H���MO�i(��.}�M����q�o�~��x��I��٧�>�bv��=Ug��y�[Ƕ�%��#*i��WR��(�GC�//ӷ#L�@v������_�|{��|��Ĭ!]6.[b���6�����x� q�?uCÍ%t��ma7M'���'���c�n�ӷ"���%]��}�B"�}/]B�T+Z�kƽ���r����T�EuC#q5�.k��:J��PY��
��X+ Sjl��*���;� ����ͪ:�*��kI����N��ܨ�7H�@�+܆��	�P���nm����{�HgD����/c]ʣ���SZ"/�פޞ��$_��I�T�U�"�B�}�~2$e�l�tl+��N�<��%O����<�vr%���/6�����@˯�����:*S��#�+��`��ac��ȜӉ�%�vh �����*�����w�8��{��/z������J��vA�uKp��o��ahI����$�W/�b�k�]@X����"�S��29!��9��'�:�V�e���\�"�	���(��QK��9�J�~/���-$szk��1����B����R�P��v鲻S^��w�߫�­r�\�d�9Ӓ�Q�����7�G6m2�aM ��.���CsK]󱤭ɽ��w�*9�~��A�"d� GJ=����+'�z�w�H��RURR�
m�7�<;P<��B����p䝤Q���B=�B��2��Yi�H�oվ��s	���F�r5�N�? �˰aD|솼��YK���5����;؃��Ҷl�=��(	0�Hk�bܖ��-t���n��J[���'q�`���|���O�:ؘ�������\R5�
��0�C��_���TuW�����A\�$��7z
����=h�=���k�����G'���y��yI�1��"Z��1-jݸ�w$��@S�1��rz	�D�CE�
Ә��[-��bS�W|����.&�i)��|�3�i+��þ�,�I��;��R6����m�����/�|qݠ%#%��3ph�(A�o�(�F�jN|c����m�]r{�g�DC��'K zH[3c�YΚĹ�^&N�y��@���%j�%!��^��>M��� 9�S��zL�_sl쫘p+���%��.;��tN���u �'���;��68������̠!�N�XǦ�����~dbЃ-�X�"�iv�|.����(�h���D� kw[�p�p�Q�Cc�)�M�><�Ԃ�_o���3��C�&[�.Vh��w�j��Gԟ��b��d�b�Lj��x��a.[����jk;��x��i�`b��WNb�=�4���	�Z5�@����D��0�@�#�wm�	�����5u%���s�ϻ?�j[�(k��GF�q�����Y	]iK�Q�|�yԶK�N���!�؋'���f�x�1�i�s}s�r��
E�"��&H~ۦ�:�����h�ux��2�S7�JR��M9I��6�!F���G/Q�|Q�W;�NR�z�Et*�>�u�-/]���o��y�|Z5�y�i<b1&�$>u��GǮAv� ��@�MF?D�8��z1�e(@��+��G�C!���mD���Ȩ]�#@^����iZ��=��}=z~�/�`��/ō�%����n�e�����_;��L�W�HM��\
I^;���`��*�q--ː�H{��X�:�*���cfl���TQh��G���<�W��(�]��̷��7A+g�|�I�#c����W1�_t��V�e]�bM��n�Eq&K�,�N�퍟�ߍ:�.�F�hr������N�T6#�em��7��y,4i�:S�ō�XF��g\����I	���qC}ᠪZL,.�߃�;~�v7�҉���|lM�KZ+<����` ����c�^��� ���kĕ��"��"Z���;)�Fv�`�!Zt&���=����ES\� ��U���Ѹ�v�@�uͬ�Y}n�����c��*\�I����q��^����^k��0���h�E���+�Np��
��:��k���y˂+��U{nF����ؒ�m`M��0q�%�0��p�UϞ��}�^�әy(��ܦb6��ױa�b�U��wp��_�c�l�<2�;W�ۖ��N���m�"'!�q�D���n�Tޓ��2�����<��&����9��1OO���g���<78��w��u�U:��~�����7p+�~���Z	�8����7e�ֺD+Z�씗ͣF �$����2v�LE��✫��+K�g��3�̝:4��Tê/㙲y�k�'�d� ���cP��k��::���͖?d�@��}c�MkH���P�Z���6�kf��5�m������X�A
���:�։.<�������V������~����W����������B�&$T�~]�jusS;r�gM��>��C����nh���M_��RC���R�(1���'$���~q�%�d6��3�T�B=��P9�NqՈ�I!�����2��=��ubН�հ���]��{Ѹ<�1W��
D%}��d���Ү��}�A<�,i�Gh1\�k7�zG�����3�j����:W�y�P�:�G���-��;���1���/j2~�ĥY/V/�9�,��0��J�-ugO��@#x�J����i?u?�������p�������rD��kgH��S��Q -���O�j-�R��AV��᳛�^p���D&T?u��+��V���v��:�����Q�� ��	Xdb�N��}6���x<j$�0�F�³�F�Şo]�@PE��M�b��M7�*���<s��ԥ�rJ,��>x�ckOGU]�h���4��la�$0ޱ�7���N1)�Y�Nu��I K�xK���/n�=�kȜ^�dQ^�xd�v���_���/��ӡb��BMD#�LO pK��E�%Fd�;ǵ�Nc�Lx[Xݺ�Y�yڑ�'��/����Պ�ݬ7��|k]�����WB��-����ڒ��A�(����bN������@+�g.;l�aU�8�a���;����ؖ�R|�ɽ�_��PSN���폈�Gz�ݛw����@o`�c?�����u����na�xB�����2��& �8�����;��k�TAl�6[�<�8�;G�%�U�>�[�j���[ډ�vGi��IO�T�����c�|��-�����A�B2�Tn�J뜄<�`��Ό��*׻�ч9�5�a)S���U��{ D�������q��{���ܘiq26�Jv�q>�¨�O N?H�[�o��m���Ƅ3�I>���w#�N%��D=A:xk�|q�#��S(�o(� /�������f��r��X��]`�5�j�� 1�R�8DE�K�s�{jL�\R�I��~2q����f� ��Ԃs����܍�L�\�1���l C�����^�Q/[�q	⤥��L9�՛p��䙹�h����*3���5��Pk�A�}�
�f�(2A-�K�u��HA�����G���ޟ]�{q�Ѯ+�_k`�U�ې�dM���ጸ
��ܣ��ɨo�a����	Y�BS�+�.p��$a��^Pa��b�KG����n�,���D*E��!��t�(�.�P*��l*�i���1@4;;�"�R���`n���at+�UH��q����䘳U7�1i^x�\U�d����k��J'u#�k-ܰ�°��@���I�¦	O4֎WO�o{��\�u�Y��@�N'�{�fW�KXv0��!gA�������K�r]8#���J{⢷H c+��ʹM�u��)�]�q�"���jB�rl�r�ϋ�'��^�u���A����F�1]�ٳcY��[�x�1J55����b]��j�1)�Ƕ��g6�ٲr<��jB�q�}�L����	��b��!�z���I
,���G���t`W��_e����T"�����̌P��6�e����Yz>v:Lid{��ц����(������S%�k���OL������ �Ӷ���� �kۼ$�0��}VT�k�������,�9u�!�i�4�s���,�g�9�J��,#�L}v危�_���z'�k�t\ר�u�m��(C��?N#&�w�{���mUWO���Jd��Bk9�q�۩d�΃��(IqI��wM�yJ��*����H �b�H���tb�T���a�Pױ]w�	3�8!Uk���1�5:��	}ñ��3q\F�:Js��oQ��3ҪRe-���R��x. ��c��W"O9�X��뙡'$�-���8�z5H|#nW*)�r3z��ƆA)��0]���������_`_�₨�:��4�j�h������0vV�,E�d)�����!�ܾX�:�e#Z�Nʎ$G���ܘ���V���K2�s̐/����x�c�B�r�Z���N�#����\?����:�#�*Ѩ]1�d�X���r�D�_v��=u(���&�
0�a4 K��2��:�*kSllokk���%x�C`y���9�O]a��imq_�5	:w#�c֏o��^�Uy=+b�]vĒR�16�fZ,>��O���+�ƈ;�)x�F�d�ظ��?__/pk7!�j^"�a#[�m��Fo"b�\�j��a3�q��i��?�tK+�Z��Ox��� ~D`� ����z��q��Tr�ZR�N+�n��7mb�2ȶP���*��B9�@�.&�j��S7)�gЂ1ڍ��ì�����E��p��T�\Anv�����D��7ny/��'�(3�"[���z~�Ϥ�k�3��*�lξ{��?z���Y7xp8.scLS� 玕�E>'����]
�����7R���hJM�T���ƿ�`��ח�Q�
����u�/�]7�K�=-(��PW�Y�^S���!���蕭�J���b���K�������UNY�V��-�����/����AS��k���& �+��aߌ�'�|��,�e��u�Re�K�[�=DIJmS:MMU�a�b�*��i܇+��O��E>m���Dj¶:&֙n3�`3�:���f�Z�O�]y��P�{���=پ�s�8�Xve�׺(Kn�>l���,�d�%�=?�Fƫ~X�l��s!c�Ɩ߭;#.VL������}�}Zt�I��N��CƱ�&�ڈ��\��]����JgU~�5+����SՂ~����H�J{�DF�e�h��ˈZ��t<�"[W^���{��P�K!FU2�5����s�_� ��o�(��0��K33��e������7��X"`@E�X�䧋"�T��̉JI��aX��K�V�k����4�5d�R���<l�n��3�!)��4X.(΍�0R%JY2J^B����ZD%�q�M��!*��*����;�����Q��K�ۄ���z��&�9�S�?�$\�`�Ȏd��'5������;|���;r����_LЎ:|_$ۧх��+*k�+f.R���q�- *)r	Y�#i��b�\�:��b���5� }�z �тL�aQG�C�>�Y������?D�!�zG����Yj�G~��u�,q��u# ��2c#m �H�4&u?�	�˲MWG�=yX�zR�-VV-����C���7Z�/Cw1��XF��?��eL�	�\,��9R���Y+���� �\��7_�%��[-4��9$i%�������(���I����"�|ΔY���Jo�,���R��&���f.��5
��VS��v1�L�rs;���^���ϧԤ���.�Z] e�٦��Y��F��s�����F���ʄO�~Fzo�=Ɇ��/97h��U�ã���$��%T�@�V፡�m���V��a����w���+�8��¸����Cm���Si�JhG����b���*_e\sk\ޮ�Á�6 ����h� �,h�Bs���9���+��-�o�%|��Do%�oO]tf$�[p��E�D�V�1�6��ݩ���=�/�t�����!��}�v��
G��\��b˕+��%�}��)*�}�?�%�lm�闠t��K�=��"�TtX�ǚ�̟�N���2��z,�u�D����n�F�˪H\	�!�]�0�K�fWWh�i�x����P%�����eU�kg�-O���B�Ӯ���?/m�}�z�'R⋞E�9:-[�/Ҍav -�
�ý�˚h�\g�2cY��K�|�0���6�V&�����ZT��'��ų!�	�������P
��7�'
�%�Z��+O0��^INF�=��Tt�e`�b}��L%�cq�>kT�O'�X%�a?I���8���S��B	9HC����a�7�`@L��?�Z4T�̘2M�a��r;�f���r���}�ogz���A��V��T��㏨��z�h��pǁ ���ַ�.�Vk\��4�4�;�īh=� ӹ����#��x0_M����#�m;�ǋ�_������'�V�����[��$��^�����E�ڊ�]�S��%.;���pҮ��N�x?!*@B��.��ı����,�/nb�*Pd8 "��*#T�T`���~<���z@�5:�H`.��h_���ͬ����ե���iBoc�<i��3�/�-�\�{H�c'�Q��¿��_�H�u2,ho���Չ?��D���\�	<��vޔ~�`(�KY+����X�lx�p�����o �v�yD��kJ��B3�x��!xu,k�*s�D/�&1�TvC_C��Ȭ���Sx�(�5X�1�G2���4%���w��!�!^�"��s*_��J�P�p��M� �&���m��HB*޵+���d���m#aN�yI)K��t2��!���9l$e���ᙄDYb�*��]��U��"ѳ���O��)fLˆ(c>
PZ�X>����q�̝g
.�؞��8��TYQk!�/"{�`ye����] ���]g��	�Mu��� /�w}~�O��q�~���m&,"�I=@����@��߷��4h�O!t�	�Ȃ�͕�-h��HQ\�Fa"t%;Z�$v&���Gp�"���e�hy��$j�L�An�&����XZ� <.0,�wP�%���p�P��R �a1�Ba֗e��8f�L~.�`$��h��a/Q�_��o���		��d��^�������ك���i~�t������u(c��O���}"ah�#��[S�o��0�g��mqj�<�Xcy���@2.�T��Z�2��0��|0���)+�G��}� �\xg��X��|�~����v�U³&�w���^O�L�?����,�`璈��R&I�X&�y'x�޽��T�5��� ��ݳg�U����ݵ�~U#{X0 �o��۞G����M
=X�
�:e�����i ��8<䞷�/$\��Mt�A�K,��M�@�Ƈ�Q:��|�)���)�pL#e����'��cH�"�r��Z��m�A�,N(�	�;aS�t�>�8��}>Ǒ���g�bv;#�9����׃�#f��~_%P:�F�'OĲ����'Ck[Yi
��Zs�j#�Q=��u>��j^E��!E����F$�b�����I���EHZ�ծ���q��ؔo�oe�f�m�1��k	d�.,�~T}Y��i��(6�v��4!�a9~*A)5�}�qFqc�����
Sh�9�F;A��δc�K{<�� MΦz�eddq��F�e������������]�y��a�*�ߦn��QJ��R���ľD�q��@�V��.��(P��d�-cҞV��|U���W/����e�7�O��qָ(�6�y��!&�/��>�/ߠ#��t�|��vy�YBn7ؐ�5V�Z�T�鹪�f�-����>*��Ƕ��iR�+q�ǉ/#]Ҙ���0ۊ��"��`
����}�#�RǣbcD���R��|ݗZ&�-��=B�Z�<��M�t��9����#� ͐ǰ��{��=��V�z��N�u�4J��ҹ�C�e���ݏ*�h��6��L��W o��w�ѠkuV=�:�i�w]�
��X�+�E�>��<�#��篡%v�$���tp����)��+!5Y]Mf+�^D�.��FN�C���@���Tk@��
"��{��_�?�8V��Bp���R��^f\��.�>�"�
��c�@���+��)�ar`d/���g3-�f�y���1�ph�-K�!�����f)��"�^:io���FY�q@����o;�0V��]���䛊�n�2�0��\Sw��Q���)�|=�{���Er�v�0�j����xn1�����J�|�_�� �����xY���#��S,������B��v�s+W�/.9kGiE�9�꠳kЅ���!ߘ��8P�:Xi��\=W�&��"��]�q�(�=�������=4Ȥ�$���>턯�V��R�����̻n��%��D�]�AaBm���=��,3�:��M=� ��*�D�Q�|���\�ކ�\[˾w.����b�+�{m���_3�L���l�G�� ��^�d���9� ˓}�2+X�X^�CG��"H;ǫ������5�b�2��I��B��C���rqe�Ƶ�e�G�՚.�kTͩ^y+���_X�]��
_<���e�G�&k>x�� �:�!�{��������o�B�h]���2��ȿ�%�Ft�8��p�Y��	��k!`VqQ�P~U&�[P�%��0���#n�Z�|3(��ET�yƨ`!��B�U]7�$���_\B����K2�HoS����'+Ŕ�,�i�}g�P�І��h�7��0�l�{-+;��w�e�ʠ��+�K����L�`o��ml���7:�$u���LFnl�"��B�m_�v�Ç9��vA�0����k�mRO�����ʽ�7��7ҫ�Ր�]����G����8�����W��Tp�u�0Vo>�u,sUY��h�o���`/���NV1������
ʰ;�wucu����&�}+����v��ߋk�lo�K��j�v���7}(��ɚf������</�}�$��	�'쁍H`�3�׶�H��ܱ{s���+�f�����[����y�X��Zj?��+�LSf��ҾIO��]�	'���<W�j�iPSIޱȂiYꙩ�����WRp7BU��i�$����D��C[�b���53�3ˉ��;Ox���j?z:�@sp�V5|��Ɠ)���𛥸k��w���aK*���4�lyvt��V�vTW���\�*�t{��6��ĉ�8�����q�a9�� ct���t���nl�,�E-��̇����%�a��W[�i�(���)�9/��1:Wƃ�;�����bG��(����F���[�ۼ�f�	դ'[^�d�����Hr�c��F"���=�.VB{�zk.򂌞���O�����|���+[���OX�;6k��͔����[��ߵP�]�w;�'�8E�N���ky�NC�SH�l��e�L�z�q��\X����XxG/T��
"����r9����eز_T�	[Ɍv���S!R�s��Pu�uyZ9�&p��B��4}��l6E�����{f"�A��tU�(�"���w<3]�>,3*��䦞S�ҥ�bԤ���n�r�f���
�-s4��cI\,-��.�d�P�z ���L����M�Wq���%��|C�ë*JR��G�X��z�Z��U>;h��'%q���O��z
-����.R�����Vtqr=�J}�0�[s�!��K���_�Py�ą���瑒�~R@d�Ql���E>N���]��5�r�T��[�m!9���)4{��(yC�qs�����Ϸ�L�� �kz`ݡ�7f{����#`�V�g4�%W-�	�4/��!y�k?{6�a��3�����O�}Nm0b8t��F��X��o�b@�hD���\)�b�!�>�Y�%gL�`��y
��m��39�y�y�[#�������)�j=�4���_�en�V7�-���%�PU����y�6���OJK�]�@y�l#\I+��HB1lM��[� �YH��V�T2A�m���R�ܠ/���r���?�a�4��0,��EN�j����ݴ�]���;�&/"q�X%;�I��_��U�_����[�G+ъ�od���<�X�g2-J-���*P�@Y��_Iv�uV��c�{���6��><l��q�.�Hf�Z�luM���?��\%EK����f��l]��o��]�Ją�H����W��r�j� ��D�0�����㗉��x 9h0��[�k�O֊k'���R#`�9�=5 ��Q2`����LOfѵJuה�Xj		PE�{ѝj�ʎQ���x��Vo��öN-�������$��Y����-�o3�"|Կ��S:��{���n��M����h��`8�$��0 ��'D��ou���� ��l�]�7)�Ƭ����HN�Q�����t�PJ6 7�-��d7]����E�+Lھ=��N�+��!5�G�����^�~~�۹L���'ؐ���[�������B���k����
�h��M l�X[�ff'
���|�kX�~���^�q%�_K�4����k��f�T�%E'Čn`�<��7�.+��tf�XW�^M.�1�=R'=7#�d�^bӆ�h��� S�r��[D���S}C�j'�����R��a��!�+;m*lZ���\��tc��ل�3�8�T�q\�>���L
)0>L���6�`�G�k��.���;F#��u�g�Y�v�]�y���M7���["(ٲ
c<��Iu����y��hu�p5 4W�H�uj~�\�}�?X����\!�6�ky��H"�!��A��#�z���ݬ��8���T��j��Av_ִïξ�ev"��x#��y����lH^aO<�vX����L�AM��߁XK��w�{��=ld�l��.t;N�,��ET�}��ЪD �[�Qy��j����P3������B�!/���J*�j������.�a�-y�u7�߭M=,X0^�:�^���wݮ�(���U�)F��b�AL�P.�8Lջ�"�IqX�9��YW%��q�婹�_�*�^��S��ŐV=��'����@���{�8O$`3r���g)yS�M�I[5ҧ0:��k���K/����K�؇���
���b�Z�a�P��r��y~��x�)�Ύ��2]@���B/߬�Y���Z&`���V��}�l���tޥ�#	�c�<(����ﲪ!��|G� ��1>�a�i���-{_r{�*���C��n�8K��=�Q�cS&*B�:�!㱢�{�?)�1��kM>��1Օ��Ua�C�$�6� !��)XO7�?}!�Q��#���"�����j V�a��_;��J���{�u�R)����M��w�ծ�����L�OM&:	7\+�_��0��U5���s�a>�u�����x��fp):t�;�| �fPy_{d!.n�9��:�]J��>����Q�9}4b)
�|�M��/�/���cRoU���P��;4La�KE��M�3���P��Җ���*���>�t�z4cRp��, J�K�6N�zӻI�\�6@�̌P�������~����^�Y�1�lή��O[e!��x˰�w�rgB
���׭H���8����<?�Z`�I2nz���x����@=2���~gi�,�,���+���c@�=T�#��|cz�:����2��
"���H��μ2C7�/zf<?h��qi�᲎r���#A�yq[���.</��4��e�W"��)�o>�~��n���U�#3|�uF��߷ �I��HE��*�?l�Z�ۊ��F���$�ct����=~��HA���}���:M��TD+�E�}tm�u�H7B�7DIM�ZwC��f�2�
�{8��	���Nτo%7��Ƥ�w֖*��'�������4�>"��F��0�NnA�ƦtRgi�6/���L��~7y��W$�yf !OJhY�p40T`v�pݕ�-��ސdr�WC<-�/��h�2�!V�1�kO���Kص|>��83��$��:��}�(`^�q�?��(}�#؂�b?=���*�+ę"n��OD��P�d���B���]��1K���M�砹l�� ��,_�WA���#�Xy�r�����P��0r�G��/�,��$���u�O�SO����w�m.�t���d��(�{���٢�E�1��cH�ě���c���{^��ؐN���i�|S��t�\[��B���> ��u��t�9%�K�}��&��k[vm��YJ���ט��T�[�G��Kb��S��*�V�N
�v��s�t�2A��!bm�DM���WrN��������Z���_Zh��^�"Jۂ��r}{��Ua�^�������g;ղ���Hl*���/(��aN�v,SM�"�.)Te��݃o;��d�)�9��[l2F���[�%����f���/UЮ��3��:�ר" �>մ�3ƍ�c[T����
g��
s���d|�0�kA��+y��m|̆1��4�d��4��{��5	Z�����*����|�*5?��K�dbT�]�}� 7�U���� �)�V�m�mf>��,�c�mUvxUq�t��q�K|#K�ʔ�����������ϯ�P��'H��rEQL7��2W
` x{(�bx�����#��^����ÄY�$H%W����q�@�z��,Dm.���l LD�D;�E��M}(��^���z$%(��Qʫn��%m@��8����Y���j�I���ԯW�X������F'�4[Z�e,����h<n�W��p�R!э���oM�K���R��%�t�8E��5��j֭?߽'c˵���"���-1�U���1f�_�$�5�ָ�Q�a��޸����+����4�`J0�0���
�8?���Z��i��78�Y�4�-t� ����\v��2L~�'zKaz�mp}�_K�C�P�㉿ƍ06�Y��`�(�(�N����4W���n�4�ؗ��[�t�;�x��f�5�M�
�p�!���bXqz���h�"��^��*gJ]��_�D���o�i�:!��f}�Xd�{���C�gT���u.=-�uvR�㩁�ę�d�xT�V��N^]>�R�'G�<,sxi�I�6��N��4�b�7�g�oA�8�h��H#�6�J�J�7@����j�##��� X�<���3L��W�t(��+q:d�>�J_\$�-�Fl��L+�#���0�|ɀi������u}�<u�ڬε#�j�U�<g9k�/Q��LH��b��`��/�������=���eգ~=m�`Y�p�����"|t8Z��7�dV�++���Ѱ^����`N�!=�K>����a:��)u�Z���T�笗*%kH���<�~2E���ޣf�l����މ��|���{��Jf9��`pD$�b�ǹ���`l�DZVԹ6�cݾZ
\�4�7R$"�4j��s�e,p Q��4��pe�/�\��;i��>f��,g'z_�]P�ڡјe��(V�pKZl�uRhT�m�o$e�����܇�k&�H�J}��ǕZ��,������5J��9�Qߘ��(�>R§��$�-�\	Y?v�@ps7�]@"�7�Um�s�m@{�dexKV�=CKUAϻ�i$� �5k ��Be|��#al�x�(�u���"g�>���e����e�������/O
����RD�3�<�ᐞ7�����G�L�D�r���R�/����;`&wnr_�e0PlF>8���c��ٝv+��jC�yB+!;�ڴ�gM���?U�g-�kr��`$>~=,�tx%Ҧ��G?)=5�2.�5n-4$�MTlFθ�V�PPֽf(�Ϣ?慁Ե蒑P]4�E�E����y�Z�`���\W������;v�!�=$�L�C,\�W}s��P�K5��r��7�	�_���2�vL����V���ƍ�t7�R��"
~Eu��p��I^|�}_9�w���/�QY�\�g?KL�-�Ҩ�Fʶ��]�m������.5�qD(��Å�ca���%+���	�k�?��À���U�^���D��ek�l��W�Ρ���l*�/���	�����0�ve/ꏃ� ��k�nSq��
N�>���Э�ȥ��
��gOI(J1��=�_�bR�TƟ.ਂ� �ȁ��W���H����)����3_hv��ܖN��Z����B��uhA�S�w��#�/-�?�]�=�iM�rW�Z2I������f.;=�\3����W�uͮA��c�ͥ�t��2��xp��h'S��܋�_�֩�oaYL^���(��4:��lv+ɇ�$�9%�OgN�my�B��~m�/T�5��>�y�V8�u}�ݲ
���k��(�`h���*^��s��
��+�B�l�E 5I�P~�l�Ij̍"����a�M2��lY�:��r7C/�n��W�'b�ܛ��3��3��V���C�s��}�P��ҿ�;��-e��L��� n_gFH��TI���Dn�M $������j�S7b��*�#��`�^ |%x��X�0�M�&.��'�����z~�S{Q�.�l=?�
��o�l_\�mCNޣ����4���(_v�9��Q7'�ْ���Xj!Jx�Lk3�v=� ��ܽP�����|�A�R��X�}i?u`��_d[ �!�V�7��L_���8��[���Nj�V*I@#���t�!@�X#�O�`��Jf �v�2hl�I�;U1�ΐ��X�jB�[����"�;"dLSBi�>aƔ�Ү6Scb*��b`[����?]c�u�X@�	�w�A��B�S$�ӎ�����:�U�0&�F��x���y�R��7�w�[�����]�7�x��x3��j��]�������F>��BE�����7`�}�-B#�k"��Z�LF�_�Mb�09*�����mk��i�<��Ӥ����@8�<!��8��ɻ�AQ�__(oح/?Py���Xi׌�O��}~a�����84i��tsR��B1�I�k�P��07M���Q��VO�&��x���5��z"���ʸ���1A'�����ץe�D��v0�����q�;�1y�5o�a�F�)B� p`Reuz�y��+G�,s}�x�1��=}r��Z$�Ø&�T����>�,h�0�q�A�Z\���ef��ڨ�ʧ�C/�%㾟 PʸX�?X6Ej�\�f٠y�q�<d=���MQ�7'/���B����B��Uo-d�e8����zaPjC'�D���<`1ҳ�h�(������	���b,g_y��qE@��Y_�c�^�N��̠��O�"�IR�;�OA䍿�x�w����s<�N���>�P�Fq�~�b0AJ�[ʴ���kp��Qi]�7�زcau�x�9�ڈqn�h�MLB�gJ�#z!;���S���X=7�SLj0���wɵ�OӖ&���A�}��<�g0���`�S�0s��D�V1��ʕ޾��UK]E�Ň�ΔKbBp� 鈡!��M<ny�bzy �z��)p�.��iWʍ��R���.PgLN�x=��Z�l�ɭ��
����;��n6�85����������~��>�/<̼I��;��y�e1�� i��^)wQ5�%�N7�h��f`7�C��	���S5�_gh��RՎ��홗1����b�bY���NI��8N���ό`��iIG�eHE-֣�e�h؊��X�:*���+D�>����,�ڞӊ�=��W�QC��.`k}�j�P2�������	=�SM����l��`1��QW��ٷ��-�w�.s�[�|�iP�hU��C��(%���E�o��DV�e�$_E���H�,�q��6lՐ�*C�=��\���6/:�����۠;�����V8�q3眬����1zkf>���~*Yx���-"��#2�=@?`HyZ�k�T�}9��l����g��F�R�pV�	�w�k��[ ����dwؖ�*:[��%kz���ph6(�w�_��]1��8�O��h��X�Ι�D7׫9��)`��e#���{!�x���$���#@v�ؗ�_�q�X�N��z1E��Nr�}���K�z�d�Lz�S�(��)�+����o#��/��C�G��2Х���#�M��}�w��-r�5�o�%rw8�O?)���K�_�g�&��6��rw�.��}ݔ���Q��?�5%�.��Q
�͠�b|B�����F����O�h�u	��ZC��F@��h���w��I��V>):q��Q)�`^�3�,\o8�V*��+�I�!�ci����AKI�e�E�C�ҋ�`�ݖ��}�|���ў6�^�,O��}]�Nm��?w�C��멽R�r�����ʵh_\�i~P�_�^,q9����EV������%	�����ڦ�h|���ގ���9�!Ջ��.���GN���:�pf�U����Ot����*!��V^�3�	�x����H٘�:�3Ǟ�=������E"f$�����x�U-� �ιQz� 0Bf��P'��
L N��_๤W��"/9�_�1�^�Fe���-��Yt}O����փ䜴1 ‧&�
��%� �M����x�}�U��t]c���6K�?J��\K��~��JGּ.�+���8�c�x��At?=sM�����*1����Ұ/
����F�O�7'����DE{��7m��jȘ�/E�H�)�t�U�8�ɬDZymd�S��f3�=��b�]�]�at�wr��3;�z�Bǋf��Wp@J����C1-��*T)l��=��2^e�} �F03e���@d��C�EC@$#��/A`]��ΘU��3���Dl6����+��}ݷ��W�y�hp�L��t����9S>>v"���Q5A@�2�u�J�1����̹%��o�[%Is�?*�%!o��Mf�1�Z�/)�j�hkMD����[w2� A�Q&��3i�,'��l�������S���+�O-g#N��jм�?S�}R����1�yT}�xi#ڕ��u�ai��������n4�ܠJ�)���Uk�;~/�||��yK��m�=<d�FO�q���I^�'�����YaJ=N$��{��M:9fE9�V�}�T�A��T�2��]�zV<�l�}���1��i���!<SVcj�bD
�� ?
���M|�UB�zɕ����|�$x�f5��4AuB_߶�ݧ���&ի��,�Et�<������ևq��w�>0��N������'��o�{�!mȘ���h�ʰ��Ên�9��}`��U���$����������џ{�AG��ZM��(6��Ӗ� �r��.��56�ɶ����Y�$a���1qϞ�c��,_RP�7#�SL�C\	t+$�B�,�)�ʈ^(���H��KF)SI�4�Z> /�|
$N��_���V���i�u�}���J�,�;��H�m�ٲ�0P�������GZ��ĵ؇9��j�� �l+�a�	Y���l0]�sٸ�8?2綦��*��d��P�i1�N�P~�(K��%�~������ߜZ!q(���'���0���{G�ү��U�u��\4�E�z2������;x\'��e��ἠ�_�@5�A�J��.��wЫ��*5vQ|!�h 2� L"h��g�+���<�z~�L�|��h��J��,�]�te�@d��Қ�D�>��UC��D!\�1�
~��xݳ�<n�~_��%C�R��C��M��e�r"�u^=��u���.���xz�h7�W ��*�N��j9|HX+�֒򟼥t�M&˗�2q������lPcl�B����w��e7.�9�.�*]�RN#s��!�BL�����ϒ��?��*M=��&44�ޣ+L�MQ�ܟ�T1P>�xʢ�u�'��#�c���^J���E��ˍF���![��I�7J��:��*T�� �������o<�%~�(��gZ�4� r|  {4���7~ �� �Z6^������"�=�X [���]���p��f��5��BB@���/�x{!�Ե�):�ʿ	�1���XOf
�cOp��r�ț1>���x����ˮ��@�s����\'nm"b��@M�v����1�|�?:����"��\��1�RygH �/�QX�u�~���0�ze D��u�^�
t�(K��x��|�P��#���ߪCjc�w[�I�r��1x=�?�<E ,�g{�U�=�}M ue|���5B!�-�@3���)ñPw��H1י{�.,d>�K�6�2�����E���oq��]l[F2$�a� �� 8B8��Y�K�����%@�S�+�}���zV" -T4T�GX���0��B��>i��P���svx�4����/��(
�����ğ��1�D�6U#�peCMoL���)�mn�G;�oHW0 �.��5�^�v���sfr�~q*ɵ��Z�4F}�',�OQx'�Q)�Lا$�B^�>S��"��1�mI7��&WƸI���������"=w��&�4� Eh�l�Ah��v]*�v6e����x��q��?%Ձ�m�&o�'wcKקț�m[��,[aj?��\{��&gv�yyTJ���|�{����U��uUk��46g�m�wh��� [w�y!"0E��rK�]���٪�� �&o�}9j��2Vi����x�e���R�TC�� ��N�f�V����o�׿�$�uzB���4!A7��쇸)�H��r���6������K(VV�� @~��H��)�.S�9������ٳE�Z�+A��7ʩj��+5kL�3$4(��;g�.o�'�d6	+�Br����8��2Yj���ǯ���^�_Tc#�,J�X&��{�qR
��i����	
��G4�	�[;~i��u��hǗ���{�����w���A��XA�T��t!B��������	7����a-�T�F1��߼��w�!!p�9�wH��P��gF��dMeq�+�Y��o~���mM�3Ų6."�9�/�"셮����	��Χ�~5��ؔ<\^MP"{�]����D�
��_�������XD�P��cL�y:(ڪ��p�+�\OA΍b�&V�VU�n(u�$O��R�F��=�4#]iK���\M�⹌8a0�Ü������h��::R0LL?��י�W�ik0��&G����M��~��P���-8h�� ��l���]oZC ��C8{��UK�����
)"(d��I<~����ϫ����/�op��l���0�"Ċ��U�1����1�#[S��\�lDΉ�9�P������(<��D3b��b�mj��~�1����p!�o/y�䧳#����N-˗�}Re�t!�N$�l���~0@_L�{���X��J��55�ŏ8)O���~Y����[��0��T(��F��I�|x�I�im��Gy���<�%�$I�ސ���f�I=����Q�z���R܅���~'��?􀳫_m������ g�=HǷ)Tͽ��$�E�{�8z�m��bΈ��Z����ⷎɽT>�XA�1���C��#l��yd�'K\�|�?-f5�h�&6��:?�1�ӕ4gD�����U>{4c��*Le�c�<����g���/1��o�^duǽ�|r��>�9���������/}|�p��+�r�v��N���r�r&�i�k�%h^�H!�D���`��0��X
ú��n���g�	�'�)��x:2�:eέ)s/J�>�"�����P�Ɵ}$u	�y6����M%h�.�v�z����R|��xT��c�vJ�`�h���7�k�ˬx��#"���Xt��a'�-~HżZCJqp�,�g쯔gi<d�w0�%5�:����' Wd�����!-5HIH�4rM�s����w%l��H<q~2F�h.;YF�5ˑQ��U�ԯ��?c��ܩ2�i���2$�E!�à���Θ�G�TB�Ǻo>*�]]<v8Q�v���`�4�9�\���kE�r��Z�#ɕ��F��x#���ݮ�`�=��`[d�sw+����+&F������L�:��a������%!n���������M��aD�{)�`��(d�d��۵�W�Hh��}��S:�]�Y�3魻�c0
�u-��2'��u� ���rV�X�H r�i�v�!hRw&Y��ϳ�;�diK ��>��FЎ��]�����g����>��s&���裂l���1r�_��.~V���(�2�H�|�d�Q�H,�I����N��������+��"��4}�_��<�m��23�ze0aj)��[,x��a��t9�-
��e��I�+�9@<4ȴX�O}�K(�H�`��x�����d�y�cP��T�H�4G�L�\�A���f�eQ>88Ӊvz����󝷞M�m蘡�C��Dr�^ߚS|!wM��l��o&�{�E��s>������M���:����'��d�i*&�,�"
ĭ~v�{�`oO��?��[Ip�I�ƹ�Y�r(�pQ��J��k��!�^M6���ش�R��D9k�����{~T�Ω��/��!i��ڠ���:�O0B�6����m�0)��q&�~{�e� �zvKH�������������d�b�k��]�æz~�)(�ׯV$���I� v�D���f�r6Ci.��k�WQ�6�n���d~eC�	���Oe��z�/����T���arf���uPVI�͏
��d�]$��ۭ|�[��1$�����[>�T��9U��ɺ?K�M_r�X'��1�"o7u8���L�yZ��}c�UV�]+��ibJM��^�Q]rH_
%_�����"M�a����ꡟ�ks����14)@(�O�IM���7���L�P�;!ń=��Pu� 5����'VJ�Gi}�I����?��t��;�=5��>�w���D���P���P��$_DrŃڕ���)�3a�����fhЃ6�%��)U!�'�@ӟ���T�%X��G�ȓ��`�9�f^���O��t���/��.�|Ĕ1�"����I����B�2�b�f$�ey� ?OU�5��9�RA�t��0%^�D�H��"z̃j�!k�g�Y(�gU@�0��7)�B�U���$��*ݹ?�+C�L_^�*�i4#�Z��#ʄ�Im��s��������>~x��my�BPT�ś=����TNV:LE�)�,�E�k�n?)���O?�����	Rs-n�EK� ,�)���6����<(�G��r�eȲy-~��5~�cP������aG�H�:�IXN��/���EsӇ+�%�ɰ��0�����|�p}{Y?��۾�_]E�^C�	n���	nt�#5�ߺ�.���I.����C�_�@�+��"�4T<_7a���a�V����T�)լn ?��d58�
s�۪3X�\��9�np�1�� dfd���r�4^�*�<{3��x !�3����Ы���h��B��q�5�n�����^�\P��B؏�v��#�b�z��
,�'(�i�T|.�>�>_p��������\��YkU��c��]�nw��*t���Q����rXR�o�����&��q~;=��Z�"ؗv�R"�TCv���t1���mY=��`1F2�Sp��ġ���9���
���E8��go��8.1��޽rU��<|mb����-���|��2yhW��G�)�3|�.��5��(�d%��R�Y��NQ�&�H�}�r,(�;���|�U�e�Щkf+R`���?(3|�Q���~�^��r6<T"R
�x��9������L�`GG��ܙ���Ad��$�y�}ֲ+.�eͬ��Jp�4��_�Y��;�\3����A2 x=|�<DQb4�qT���#t0#ra${=Z�+��$a�l��C��G?�ߜ�m�������{��@?3p5cs܆�)u�fr��J,�}�J%��1$��[p|��Ѓ�^d��cGy�Z+�}s��$1��pK��^�p�$��rv|т��B4�g�cLS'���d u�Ӟ�w?��F�Am�@���` ��`!(�x�>m(�i��EV����5���/~7�*	\pQWF�R���ey����Α#jZ�����V��#�P�P,N�y�Z?uq�a7]B�֦T`&�����̿��0���/٪�Q
�k���[�h �B`Gw4^�Z�ꔄ*h�&ϓAйF���^�`�C�O@^�� �#�$���'�v�.V�7�����o|�qNkO��WR��#��f�=?i�D�'M�yM�?MH�U@B����"�p�o�k� ^ǌ�$�咠s<�E|�j���Z�b�O��b�ׯ}o��:���B\�u�2Ә�1���L� �T�r��s�:�xf��$Eѹ��8(�4r Rm�������1K'�Խ�x����l�f�뉜՘UGŷ%�9S N�-
�Z"���%�t��J�&�~0u��'x��⎵ݛ�S�w�i,e!؞@h]^��=�@I_.&t��#�&&9�.�8���MO�m���Gz"v�6����.�;�`õ����7��/��]�&���ˀNZc.�	��<���>�me~��$3K��ĪW�:�{S����_�X��$f�kr�pn�����N�}*��t�d�j���[�t@EB�5��^��{΄0*�DVy���@ZS�՞&+��ӑ�7�V���ރY�r�B3���[!h�i���Kk��=�Y�'������`Ƹ�8nQ{/;=����5�{�2�Vx��j�ﯜY?o��v�v$��g�!���7f���Ud��$^K�Qz^G�^9M�NO�դ�r+W0V�x�vR�^;z*p�Y�@8^�MӀN	꾙Yp���2~�1��GhR���$��`�㐓]0�2��|�7�}��*7�����CCD{f�}���m8@����{�37Y�y.��:Ee2�& �����F����Ǘ��d�t%��
�XGJ$����H+�<�'�2R!�c���}��adV����I2����q�	N�tj�E}�pXLb%�4�ɱ��x�ߥ�aa��gk����j����(��bf='�dH��~��O���؉��!��N��3Y��,�J����n��V��2�c����J��V� M��%�H���7����쇫�6[S�������G���ן r�~�8��\
�Ի$�KUQ��g�0���n�'<���'��i-M�e�<����J}�",�HI��,�k���Ȩ^I�B��i00�o7줌������T���#�|�%S(5�Q���h̡+�	�r@��_�wJQ`�n]?���Laxd����zt��n��c���N� �ԕp�Wu�~_18�>+��!&��؝�e��>y���\�L�
#t�70h��p�Z�a2��Fg/)�M�:�U�!�ӏ����.��6�-���-�+�m\!�vm�ׇ���ûZ�~���*��
_��Vq����X�wp+�zl�jyR~�YE���d����B��)�@��͆ZO���N	���/���*�Ǯ�l�:���r@�WuV$.�����8i1�������j�!��k���Ȯ��/SΤ�0U0[�?ػS�	�N��0�ovQ����)�&~-usLd�����k&����A�5ֹ�䅱&�����i k�`y�?%KF��K������FcU#|cW
��^U��e��D?0p�<�B2�0(�< ꊼ�G఍�ʹ�ɕ�� J?�2�;���SlzM�pT(��	49��X˧�t�*��ˎ�NM^4����%�+���v=Zٯ��?�[Gs�"={(7[BK��Z�j�Hd�x��YJ���N-�j�$8�_DGt�U X����̍��^���ɱj���3�-�>h���4@��'��*�p���4�>NiO�e޷�J�FS!5q/��/�Z,�;����W�K2�uO�SP$�E9N 
�?��-��>Ž~5H��1���4�u��H�?vy6~𞂝K+�pe>�%�:G-�](*�=!���F����@˹�9�.�Y��Hh�	�o�s�	��r>�/Z����/Mh'�R�"���޺.�ѪB9��f9���A�#@@��m��ք}�UKK�1�����fhQ���oh՞�l~5:I'�D��]y����>?'�Z�3ۋ�T��(C�cw��7h��.6��3޴�ɏ1��M���Ôn���(���Q�zc���C7d�h̭ ��c2�X�Y���^�'��źO+v�iy����;x�?�U^�_m�?;M�R��x��1���O��B#*�,��Ky^�����	�����mB�z!�	0m�� ~E85�d��"��n,_���i��cn��������vn�N��"�3r����"��k�ʥ�ŵ�]�׮�HM,ވ�6P�����?<;g��@,nf@�4^�,i��8$�TK���<2)���;����2NF��f�V]̚��C�u�;ڑ@gص�ͼ�Ul=�^<�d�`�&��v��9�&��S���� �N���,�&2�Ë�=�䁾 fV�j!`�ȃ���<e�TU��
kэ� n����R������g�3hDA�Dg����u��fw{(��iv�qZ5�����z�\ܧ�  fv?�ku�}ْ����e	64�||Ԓ��=��4�`�ʡWD�'ITa$`v�t������G��F�#��V���z��z�J
wn��1��m��@����>��L�	S�5ksD�Bw8��/�g����cz��c��JZ��us�����JmlP�D��\Ot�8������mE̫Mz7|P���S��9Z���&A��+��Y�(�GR�T�~������O���TY�|�;s)8�Mw��>�e���*��ë�.��M��K��P��Hז�ԡyD�M�f��:�!�Y��H���KrU�f���j�r��@��?��p���~?���m��س�%.�8��I��U��i�]U��K�b�3��X	�H �ɹ�~���ۼ�=���s�s�N}�.�1I�Ce�z��YڡhC�Dt�]�5�X��_���r��緾�Z�X	Jf����o�9��|f�������P@�@՚#�>�� P8Z�tb��{�Au�e R�h��+*�@��3�nч�t�Akڑ�N�����-у���9c䬘GZ"bpS#vi����q+��s4�gU�5{is}wzD8!��ߜݢv� ؐ,�)p��=�(Lo�ޭES�m����a���ШQ
:��ų�tzR��eSo3`{����"�����]l��KH-�[>��Q�u)�t~M��g@�`Ɂ�B;#���q-����|t�wc�@@{8�S��zʦ,u���=)Frp��D���#�HrR����փ��)�d����I��t�A��G�z;�fƘ���l#�x!��]��Y���u�νof'*6A��}�=�|l������I���\l�-�0n�i��F���	� Ԅ����￐�d����i��9���J:��	�U�EY��Tz�}F��o{�g���7OY��"NR`�X�|��s�G�.` ���,�����7������6�j�*��,0�dj���c��J���A$��A'N�	B��&
 �z�x����]>�/u��o�/�Q�N����<��N&{�2���,�����q-���ir��0F���CC��O�g�
|-	N,����Gw���ʱU�5�4���f>�X��[��?G��87L���A��r^~�'����aL��[����$�!�-�s7�d����_̽� ?���l�=�lY����4�T�pȆ��In`�簅��T*�����Ƞǒ�*�L#U�-���1�l���6mP��o�'�)rNw�<עLB�q�ٿ�m��fW�G�I����Y���T�P���X|���]���'u
`�t@� �11����k���Rwmǹ�׍SdJ��^��������֗o<A�d�/8�^�M�B��$H�̳��[qB?�杳%�ry�cd54��)����e�9���$���eU��^ay���N<�kk[��0�Q�'/��r�u>4ϻ�MM� J��c�;[{*�}��g���f���nHI�}v��M���J��K��>�#֗<V�~9�R�K��8�q�~,=e��AU���{7sk�ޗ��@f33"[�k9Q'<�F�Eg�h&�޲V��fI���7,�a��=ڑ-6P��:HCv������v�W`if���BH���R��I�(֛�۬�i-�d��Z���@\�!�-�)>��HS(M���)��^K�[����!Ԕa�+����#h1v�;�%G�1��(G��J�W��P"���Ug�0�I�C�������3_��W���X��U���KN�6���g���ðZ�}��'}:o������P}��{�<�1��)~���⠴�h�1�I�.���f�5��L`�a���c��E���6�����N ȍ�ם#�?5�	Ѩ�d���z#��[.�!����L�*�;�f	>�����)͸Y1%�c�F@���8��I_'���|b@������@�b�پ��8� )ĉ��I�W��%L`�`:�;��,�M�@AdH���~�8f. Z���$�v��r�o�4&>���`{݃p�|�����#��s;7ᡏ_��!��X������&��W #
�P��BBq��Ҽ>&ʁfݛmI���L_�K����DLd0�!Iv�Wm@������L�V廔6����!�Fl C�<ӍYZh�� w�ww(�5�#�^��:�p��4>q�|����/�|�]ǟ��o(<6����1�4����MD�v�a�Yԧ��=��:����5��V���
���L��V�����B>#C%:S�o&��7�XYJ���o
І0e�x"n�z����V><r��6�ɛ����+�9�w��g�)�F��.�Ǭ@����.��
�?��g(�?�����¬�X��3m�����;p�p��Vޙi������u>�����u6�z{Yov�u��3�̖�!R��k�R��^[r�J%o������R���p���%��+m߶���z�C�DuS?�G:b���Hs}y���G2���!�K�yl ӗF�2����h��S5�| ٟ���t���(��oBf�a��q����E�fޓ
m��P{\��z�/�9G�C�ߖ��1"�2j��Ѧ��ِ��J��5��y�4��K���:�ac޷��A�["?�D��~I���
i{�z�Y�/�'\L�^0M���̵z�4T�ʾ�r�?�齻���S�����ݑ6�՝�9`��&"�@�_���Ҽ)�/����Bɟ���g�Gg�mH�25(G�v��H�m��.%�d���	=�D+��s�"^~�����y�Qo�*�8@���L,��$�J�1��s��~���P�	Հ5�>�o>�Q�q�c���Na{,�륰�^�,P��ʑ�q Z��G��O�7QPT�!$�؇�'f�җ�:V%�V��	�"P�ܼ�vu֧2G2���f�[(�ؑ��XȀE���@PL3yGҖ�Ҋ.��+��2���8�=�(��'�� ��������O�o��T¼��7QV����{�U�`N�[�H��Y+�5؉q�j ZK�zf�z��vG�J7��2p�Q���30$��j@L�DOW��tG���۱E��B��S���O����I �"��V�@��pa%�A�AQ0�b͎�����$��{����
�x��b�QX��R�w�v/���f$���G��}�Z3��+Bx�%��6��0�n�Sl�@��{�J�;��=���(J⊴9�V0ݾ��&��o%�L������!��A�t�vOåqѿ޻xD��	�ܘ���;�r�w����@�p��?�P�P/ε���뮰{����.q�"�n@vgEw�pU���������#1�D]���<_'o�����3��)MOZW*]���L�V���I�<�b�u���E'�I�Q��c���w�	x�aG��W+\�<��%���/4U���hn��(CF�+��3���� ���+�&üS�yF�����C:�E�w���٧�q���a�YcJf�Ez1o74���YM�LYP�U{������O��X);m���6�<Re�|x2��לYs:�d�ڧ}�+Ƚ_���=V����L"��?��.²+�t�5�]�
ՑZ�G���է��"��%X֍��~�YT�����ίӶ[�[��}�j���`i���U�E�S�:~}�Z�Dυ&��e�4����9��:Z_��ܣ�kA������G����^�:�)����3@'a���|a=����|�]2x=Ng���k��
9���:`�1� ��p94}��Vz�pUܞ�P�d� �����_��_R-�\���9+�B�\�j{_Ӕ�=
�/^��������uK\�]��.+���z;v�~��$#���6s��*�HI�O��7.%[S��J*�5�]��~��� �����	(^���V�H��Ӻ��s���Vm`u<���,PrDLÅe���4���\�l���?F�����Y����vCZ��G^�#%� L!�!A:Pͱl�x��� �g&� �5����X�Pp^H{e����^:3�2��	C��@����� �V�v��,k��
����~�{����y
1~���=pF�V���y��S���^Kp�~4SO�#�Ġ��h���%g�q��(I�E'%̒�/�t'���A$=�v�c(H��P(3��L�qתD\�=g` � L��J���w�Ū]`�;�\�1�t	���9Y>qщ���&}�D��a�+�P�r{����^#]�����^.����>�ɵh������u�yNm�h���\���u�/��u��aۋ5���1��c�����v�(�.sġؙ[�_��/Q;�n[%�����GSL���9���P��`�[�q��Hf�։`XN�sD��]�lcmn����+�-�V���k�)jH����,D�[�+���dRf��� !����y�y��pݐv�<O�����'#M���I0�T�6�'Ї1̞���#� �=K��������*S�P���8Dj7�3��	8�Ew:N#�����Q��v��E8ad96��^`;Ò�<���M�e �Z��!�2�%�?ˇg�Dd ��7�T&�1^n(#�0�����s�d�NN�q�΅4��%���ޯO��p�2F�R�~�����yb���O�6���oT�����d���t1��_�U18�����*`����V�["��D�֎�5��R�Xy����{�Y�K$;��1�g{�u����q���P�Z�XG��6q�aa@�f��n�\��fQ��k�^p���ӊ���y\F3��+���k�_#�)�*_j%/���2�;�q�������ܚ�c����A�Lu߲q��j��u"�^!C�e�MZ3wρ2�=�O� )�a8�-�#&� G�%����↙��]J���FG5o��<rɲm�G�G����t��Eױ׿r� �(IB�Nj���P����r�N�1*�PN�#��<���AF:���z�oM�V�ɥ�pJ!�B��=�4 8�'�pRE�L,V���֐9������̲B$5ou����c����Vҧ�?�jD[ɇ=�i�J�����F�ج�N�ڎ<	5e�46�|	���ĕ���Q��6d�A'��HO��ӄ/��l��®
5nO�ᰧuj�#l��żO��gܿ�y�AK�MCH�tn�4��km[���>�'龛�c�=eY��ܶ�Z�A�*I*��3�Õ,OFr�6�O�v�Uiq��xN=��l����o�j��L�L�|�¼c����JM�m �i�=��vd1� e�����D�"�3����Ao����*N��|�:��	� 9��ՐQ��S���_���~�c͖�GΞ�A�D�X���E�,N���$9�v��0��0��tF9���X���,(��A����_�lY1�5!��8���P�oC+�X�jN�c���NÓ�X]yC@��_�����HU#r蛖�^[k���1M�bM�p�r�܀�"����� YBg�rb$Q{���O���X+�ؘ�2&��WL���~�G��&-M]�/��~@���LV����t�:PX#���Y��e���,=ʚ�cz�V����1|�]�������"����vj=S7��v[ :�D�t�q�W����Q	�.K��{Fr�I[�<vg������v[J�,))l���E_���?������6�%��޶���V֢��|`����$QKw�7�?�Z72hD0��M�?�(^��E��DĤc�k-�L�C|��:�yh�wfY�=[@�uF�"���7�2P��q�;S���ԙN�Y��?^�ys8�nc~X��o���1����}���ӱ~��{���5"��/���쉏�ݣջ������X��6.s���Z#r+9D�"Н��5��@	_��v�M�;����ΰ+�H�ψF���H��;��ӎrx�N<t��X);�$�����(iB�,��\��,��ol�
nxaͱ���y���R�I�ߘHT�k�*_A��&ym"�~F���e!1G�1��j�Qc�u o�L[9:Q�A
?�g����D�~��N>XV�2��{%�h\�/ɛR�݈h�=WyA�?�X$��ۣ )~>__v@~a�� ~�bx�8o��,!�C̍��*eh4�g��j���/�J���j�<XL�]�}��E3�-r�AqH�
�A|{|{����eM֪����嵛A;��c0�\�<֐-��A���s-�S�C��T�ŷ�bh����S�G�^f��œh2(Y�������Yv�,�5����|BVR֣Cۡq_*���+���Θ����0�E�sH�ZCb���H��V�ˢ�z�|�|�JU*J���0��]:��Nͥt�Ĕ���ݕc�
uMe+Q?8V�����G�E�'�~�&��Z�W�3�����+���M����uA�g��hP���TO���U��oۚSp%Q����P
V|��U/z���Q�'��u�m��7�5�`@���k�+�	�Pa�y§��ѷ�O�M��-.�+��c4�@{���4��՚a)*����=�E �v���c�%abڝ��,fۚ�����u�n���?�sۜF�b�5�>]��AC�x�3)������9F`����~Q�-���o��V�)Զ��.���"[��b��������r��2 ��+�>u�ѱ��쳦͞<�h�#o�+8Ƒj�z���rY�ɭ�!T2cDr��H�����b[W������7��7�zZD�u��q�A���ɧ��=�b�0]�oI�!�����x���pMX�[�6�[7� �9o'�a�j�a�d���t̤Yg�S26)�Ǣ���Z��B3e 7�^r��3�&���%�d25�	%AO��[�b����ަ"�SI��́�Ld������Y.�认|�=�!}��9�R�H~�:�rJ/�_/�-TΞ�T�rxt{şw�a��z!gK������l�㹘e����`�X�˿x��ݢ�d�~��@�A�l���}�޾�"@�eW����.�dR��ȕ�>��I�z	!ő�~��48g���̱�P�]�$s����bo�+��e�8L��Gć!�Aƃ���ͥ҈k8_����( �`�AJb�2J{���KJ3E���{0��V5��q�|��z�QW���NUSau!e�ە~�죢`�ȸ��~�D;)�-�6bgM�����T��#���������	�q�F4t ��{�\NsUk��byݛ��?"�{�kIӗ?�d��@����M����Agl'�)6_9��j�b�ra�S��Wfi�ނ�Q4�g̸w�%����Xm�!n~�3K�o쿚X�Ҳ��r�y}T<~\�ݪ�?߬���[y���d�Bv�]�z�aW��<��.)Z#Ĺ~ꯐ��!���0{�o��j��9��Ni ���g]W-k~@Թgqb72��mb��!	�\L�6���?h���{� �p�X	��K<C�3F���Ɵ��n�95BO@{�=]U�����_-�����5����m{��\;\O�������`΍�ϩ)�}����P��}b��x���i���2!��B�?�����~�����ɳ�]�����P��&��o,zP���7p@U'q�7�B~x�,�@:�F`��f%��_,",ڪϰ�T�@��Cz��(���b{(	CO-Y�e,��I:��1~�u㜆Ct����#�<�����H�8���c ����Qm0P������7b�9+`(�c�W����eF�����WyОc���Q��o�7"Y�53�u���mh8�?m�2�dez���{� ��%1_�Mb��J�D���ۜ�睓h���	�h��c�dB��;�R�����S�5t'͍��r���N��SA��q����J!�/}`�G��\Z���Lq��3�)�����u\gM�6���F�u"�O��ȸ��M=V��߫���m��%e��y���-C��|�M%�۽V+SԶ��͋��qz���>I���X���g��8�YCX�-t��u�2Q��u)E�E���Ξ�T]K�u,ov�&�la�Y�~X�H��_K �k��d#�:B���W��j&b�u�$$҄J\�g�E��YsΘZ8ٗB���)bQv�;�7�xn&=��yaV��	d@�fX�~#;U�酡>��v@�vl�����O"�B	�r�/�����o����N�:W�2v*�� �����\����*�J�� ?�Ĩ��]�;+uǲ�I�~����\�brZ�~~�o��s���}q���M� ��/����B�e��լ�c�{ lN �-�~͙��v@;�-&�ŧ0C���޹�&.�C����r�k7�;]	��)oجT�<e���������6t�
D����l�:}eS&�7Tã��u���|q�Y��,l�Vtє/��>��'�F�����g3��ME8��e*����\��+�s�w`и��M�2{g˾Q����#nIjD�euvҾ�?%B���/:�]>Q�(F�D��u5?��i���1]13��W��g=��a�Sb��$�S���PZ��u}�F���pdOi3+�5_c3�{����ӊU���u;�(�i��b��CT�r Ű�����j�N��?	W]�dw}0��*����a~ӭ��u		uC��)���0æv�)�߇�e�����-�W����]��Q
1Q�^@I^u-�R[R_�`�+ [������&]�f�>��}<��f��++�v�ʕ�1��F�E�>Q-�8�]&�3U��M�gD��%��	�l�Ȟ%�����A��@kM
y3!�g�Ļ��J�> {m�2?ZU<*xe�l�
�f��sC	�jF?v�aꗕe2X��~��;.&G[e���]�!�Q��sw��[��-��:�ɲ��l((K�܌�<J�0��aV�܂�th��@�+{�����o�:\�i�~ۇ]�៮8��[l=�Oݝ*{X�u�l�ԁ-#�|���''׳ma kA���<ZZ!E��KRr9�1��P�+�Ss���;���������i~^r����e:-�
r���z�X|\N�A������1&K��~��
H̾'`��Y�ɵx��,A;!x��Z�1��Aj�׽�S�A�HO%�N�6\���@��v�^>@8�/^w�Ȭ�T�9	�_��w��E5t�x��yǢ�`��]=6D�׷a�&�	<��}O��c	Q�^�faoJL�$x�÷fY���q�׸TN�>��i����j��&�y�Nv��ϡ�aM;��L���<���O��5j}�Q����눜���`B$[�?����'-�7�<͞�J�Wt����m�*m��0N5a���U�9-k��� hpz���|��z���\c%��`����6ɓ�ȠU�{�Ը�/�Lj�H{�Dn4�y�ٖ8�m��-�'�����A���H�H�g����#M�ͳh�C��@�g����+��ɨC1�SuU`�3E�W�~�h��|��{�vX�t��
�-p�*�+��j���U6��EC^2za�(��� �ʌ�5EhkM��.���pN+�2����^[� 78�C�/�s����p	]p����A:y����P~����c���,�/��&����P��#�\���߿�呴z޹�3ج�kO���%�g9|��y��M�P섹W��Yl9��6���!�Z#B�s�A��nK2�f�,�NV�xLw e�ګG��	��J�DՑ��Ș$mߔK�8�Z`8��K���><< ~�RT�g{�4�$:dv\��kޫ�/N������Xa$�;�k&�&˂�iz~6HrVh��,�DEU�0$�����wn>fd�Ys�A: *Tr7&��_Y�7KH9	���l[�\�r4��s[��S��X�Hq܂8k�[�m�������_w�wl8��K�?9��/@�Z�>��Ay֢;]Q*�ua�6d���ܼٗTy�&���p�WRx-�|�<R+�F//�*ywr@W��x�M�A�K$.�r�lY�|l�Zk�Y����m�5.�e��B%Ӭ���*��c������P�8,�{o��FQY���ec���m���1���p�v�39ن"�����^;�����Tů������h���W��U��6�n�kNo��z�gP��&�tK�T��1���lO��6~#���������4 L9���Du���f7]ԏ vFHy�TI%,�Y)u ��M����x�F׽�MAy?�L�P������ER�8�E%]�/Z�))����>A�Jw�����D����El���=C���	�� ѽ�U�T�i�P0|��!~�5�4�=�;�4�[D�7��6}�S�=3e�N��'���G�6���KHck/觫;�A����HW�"�Pv����=CPqE�R��;sjxI=}��8���[��>C���!��'��bV���j�BlM���BaM�IS�����2�ȓV��L0�iR.����6��q�T }�ο1�\D
��|�xo�0ח�Bo�y�Թ�)ze�?�%&ܕ��0r��gN�c�i�IWd�[���T�����1�"ӝ�Ŧ.y�cE������	�ߎU,�v���vaG��뇾�LeW���H�{Kp=�'5�Z��5����t�RWX1+5�\O�k����ePØ�t�%� �Su�����oDJZʤT�����N� as�Ej��J����}đ|�b/���sWƓ�>�w��;T X��̈́�]�t�`�O�j�U�,}~n���t��>�^R�F~�_�-��4Q�b9�v�F�EЗ��T$��?��v����he~^7�>!����S�#�'LM f�q+)��x3
�Q���R>�u��,!b�V\�?}�^��|�92Ѡ&��̷s��T���u��>,#_���^��������O\H�f�����))�l7�)x7e�@���*�u1��� ��BG�-����+y��e`A�3浞y�5�}2����1d��{+����!2g�K~A勚�E�sG�+'���5d���T����q[.dߧ���+x��ў��y�{ª|h\�l��+� ݆Ekk���DakW��Ba�D�����=Hya��u��Wl֠ԏ��p���Ӟ�[¡�MI��qI?��M��o�w]�Z�f��CD��4/P�d�s�.����k@\C���®o�Mɸ��'�#7�UCjJeP{-O��Uв��0͙""PF�����Ȁ�3��!�m��⛾G8i��8�{*�Wa�ʱ��v�����s�Z�ˢ�++���S_B��m���J��d�bZ�<�A���2�/ܶ��;���ͻ�f����ٕ���k��j=n��a����6?6{���b�X)ܲ�z�R�B�/v����yX��XG[+��oK|�E<�9|p���{.��Jr|}�O��D��)�ە!5�5����u�J�	v��Y_�Y\(�= Γ��jrP�YF��~<��-��i]�M�-KN�;/��U#� X�Mϕه8c���8�%���
{-8�uy�`�u�NN�B����m�u��o;�5K�y����ZF��;�� �[�}��)qY���LX�W�� �^ * ��,D��#�����c߽��UDk�ZY$3>C�7C��a�|n2�zu���U��%Y~spj�'v\Ґ�G��b��N����*.'0Yu��!(��H�����܇O�ߤ-u�!��2 ��A����BHf��3'0���);
CdR�M�#'����KfK���Ի���i�E���uN�i9���]q�=�!^4���K��2-�����#��^�]b�A|Y����͒���)�D�{R�|N߆�� vj⻡id���� h�3ts����[fTA=ؠ��K5�+��N_� r�o�',�<ޖ$�����;�~h�޺W�D��H�Kߴz�7ȨM��T2� Ӳ�ٴ�����7���q�YW!bĬ�9IIڈx�x>ir���P��W��$7)�!u�l�k�M���7ڬ�-%��]�'R���I��:�JR�5��M�,;�2�NU���I�Ε�G�cSxӝM�u������8Н��i(��](�OG��!���kco��늁q�$UM:��;�d�䉜���͸EO�gU�9���F��Xr�ҠG,aB�M��+�Ɣ~�s��Jk�"V�Z��~g����:���Ir� ��쥮�"�U{.�:���N��o�j�<򥷌+�|��p��kŜ��#��Ö�P�rߡVA~=P�|�7ܟ���(/(C�W�C��)����s��CQF�؆|�@��I�RE�c�]�k��^B呝n���JhJ���A|ʞ��&b	r�S��+_0Uɭ[�Y�9%]��#P}���[��uPe?V��u*B�?9�y�jt}�Hl�ӡ,��eu��U�?a�n(r5S���j5��B��Y���!��M>���AB��XC,3��M�g���\�AF֣D�f��7��A(q�@�k��C�3�?̔�������ءQ��ZY�Y�g0��ݵ��-�H�k
����(n�m��N���Ԉ�0-~2z�#���j��$��Q�����_DNtO�"K\[�vbPg�Y<��%��a��ɚ���wq91P>�w��k���ۧ�;,�g�Z�x�m�ͼǋ�j��۱&Ex��>6P0�Aαu�]��*4��=*�07�
���ߗ!�g�a�n�8�=�{��2�=y�A�fa�^�%l��;"���n7�1�7xL�(�WuJ�@a����x�H�8$����_[�hq�GeZN��$�y��E�~������mT������1D�d����gU��6�������\fAڌ���	p��at���0S�	�گ�[�=������ ԫ��=еN��#�l��t�c����J�)u�ᮠĩ�$%����I�$&����ѯ�n�ǻ�S���&T�⍚�ш{$��С������i�v,�(��Ct}�Qҍ����3���l	� h�S�C�nM��X�2�n1�9к������%� �gv��+���y���5��W�!�v##�4<U��L���Ϯ=�U��^��T�'����p�hlc����v������� �5U���Y����)1?�����R��E߁��P�4�b�&�K^ V�뙭���+�،߳�↨�N��� �B�ޙ��b�pV&�xA1�Y�n"0��I#%��e��û��3�&�m���oc��d�}��������`�4�KA~��_u���q�m������0��:�����HNOfp�E���܁e����w\�C��Cq
zsᯪ����\%"C���Xp���q��F:p�*��D\���96�R��������
�I�p7���k�Q�h�!������wʨ_��%���B�@��4�bg0��J�k�nO�����p��1Tюpo�5��M���:U�@���v~��T�����R�/�7:xy�A��Z�� ~@�>�~�wY6�a�J��4�0���	��U&��4��Vb^����5}!��Ao-��]"��"���|>p���8�ĭX`)���deds��\h�,c��qΡ�Y��FF�Ɯ��	q4��pP�M�9�Y�k��F�E�x�p�:L*b�9���ɲ���� 9L$���E%�^����L�4u�(G��� �/O
���0�����4����O;
�����c�Vl�>�r�k��Z����v��/C�:�(�����e(�J�˜�@��!�$>�e�vi�9Kv��X�N1 �+�2P)yJ�B��i)���/G�H�b�V5r~�[�h�)�k��+��yL"t
�	-�WzpM+i�sϕ���D:�5V��B��b?��3��%ky�g����j��l�pq��j!H�5��zl%�.���J��O(�0������N��"�ׅ�k�6J�EF��Ȟ�|���}6�J�"`ҫ
ݚ�VFs78)��4�������p�%�aܴ��E�#��<��5K8�elC)a�V��O�=�yO���q�x8`�ʇ_2fA��rH��OVy��O(B��V��m����5�2��������+`�KoR|��a*�`�����G�rD�
eĝRlV�U�V��c�(*G<%$��艕��o����m|���h�;&K�fc�#&���7?��S��k��h4��[��%��+,�m࿟��]i��V�L���T/����y�t�uG��[�����>���8�r���@mx��JQz�P���6F���G��yuYf��`uݡ��+�cvT����ȱ?B�%���!�(��C�x��M���
����������������q'�Z ���PJŢ�}Z�Ah������+��<M��N���J q?�$�����:�K��+XZw�~�%.�9�E���9	,D�ፁjy�Yy&/��cP����0\�4�9��p:�iv���Ƈ�j�!����2��v�g�����ճSK��5/Ӈ���յ�J�a@Wbx��}L� �	|U�����-h���a`y:��?￷�zZ�� ��p��'�$ܵnlԏ��2H>��=���f��#T�O����8��)���w $���E�3j
���S�}�m�O�sH�~� lڪ��#�Y"�[	ķ��<�v��L�T��cz����#�BP�p|,�R���Wq	`��5O���W!����Oi�*p�6�q�[sם��ͰՁ����6	M�"W�-� �����p�f*�c}����)��u�^&Z|�D-w�B��,&�XK=��ze�ᆋ}����d���Qc��t�	��:_��2ݸ��݅&�x�9����l?Pk�R�*5�eP:�x�DAH���3���{Xw�[��y��1���X6������զ�yZ������f��!����9OJ*��x����5���nb��i���% ܦ_���S�_1L�O%�����iR�i �.�D��[纯[�[�X��l�I���]���6.��������l����A_��q���n�Ka�;~7� z̦gH�w���9$�Q�_�E$��ۯ���m�����q֖秥��n�8U7(�y�I|~�EӋ̷�k9���'v9Ό��XM�/���
����{C��0��YG��|<N>��?�� �6̙ma~���B�x��y�4�)��Zv�,�/�}�~/�� �g��e`@�������:�^�А�7��Z���o��	q�p�ym}��NF�/�@�}��0�u���F��)����;cB>E|�lE���
��IhX ]{s��\�D�_aT��3�v�%w���HI��	1+n��ѓ�ޥ��iq�T�3J���T]v���
�1�@�`�כ̑�_�w����J��0m�ͩ��
�e�+b�[E��n�|ڜ���e�,���b�v��4��N�l�B��c-a���)qbr<��/u�]��S�#�;�ׄ��^C��.�A��n�վp?	Vvl���"�`ct��N�.��K�@@�s���cq������؁e�cW_�2U�9���bz4�e"�S�էX<����Qp��+%�lv�yBK�9�l�^����P�?-�3�2Pˢ�2)��>Jx�-�+��%s8޸c@!ժ�)�����;�)t4z�e�
A~^�0�||�L���MurW�1� ��K������\��z��!�
+#��xL�{t%�b���JР�����/���a��V~��A� g�rV�ESsR���e͏��lk`i�p:mc�����O��
�\�`����� ���D{�� d/��oچ�����m���F��q%�L6q�DQ���(��TPǹr�6�1��"�;J�0)��4�y�.�=���ChS��z��]2���[&��KPȳF��3��1�}ս"�]E�Omr��&��E��E75pE����+�6H���`X�c�S[���b��t�xq�2{���I�b�<���SM['����[�d��b��!�v�`c}`��Y����ɀ����<�Kc���j��}R����[���_�5��ɢظљ韫�&������!ρǱj���[�a�A3^W��l�"�/�da���P�� ���_7^u��F/�6�s��w.S�Ȥ���	�#�b�MX�գ�n��	eW(:nD���T��J���
˞F
�>b���#���Jꮾ�+�X/��D-ݒ:�
İy8�/��vWf��#b���:����q;R���GT�U�$ȅ�hB��(�U��LUE31J�2�m,L�BN\��!_��\�I��
�s���ˏ5�FPx54Zp;���ŏ��{�.��p�'���g���u�8�{���h&(j�>�[�� ⧇����=6Bo6����Bk`;��xr�|i�(4RK�p`h��`M�S���̽�q�j�mdy���|�S��'�)�xE�ӡU�0L[����p�a�蒇��A���)�8�w�٬��C�U*���y  :��ե������dB��3n"~(�t��)Cu����;�A@R�[M�i[p`
��bG��U8�ty�k>lJ�{3��h�Hm4}���D�җ����Hm[~�*������@�z�d����x���b�r�^HH2��8�0�'V{�Gm�����P*x�,����Jeߡޯ3B�S�m0��Uz}�q֕���)�j��̓B+��AU��-9>�%�c�xv��z/s�$��		o�r4��q���m?0�W�ԧ*!��ٷ�^qQL���#x7:�(y%�{����ַ�p ���o���G�A�<�|�KQi�Q��;pdi6�<���%���o�S��ő�?�r�kکJ}��%/��Q���	.!vo$w=���ѾL�ڏ���:wI@�.��Z��(H���ڃ�8�U{���#�?�I���i�J�>��d���GEv�R�qw�:t���L�5�&�4�h�r��#bh��ʢ�c�CG}������e��ڙ�KJňaS-�6�.Xy�Hf@�k���5T/I����/_��Aw��˰;0�mθ��]L��G\�������N	�t���d�3��wPow|~� e�� �	i��ځ�LU��)�&��G�yze5zÀ\�@���Ua3� ���]Bq}x�^纜��Z�)ƠZ�'s�yoAgrK:�̔ol��r�Ja&6��nd��F������)����Ēh"�r���!m	�DR����r���y�FB
E���m>$�QT���v�iF�T��e�`L�}t���c�Ĳl�M��|�QJΌn/\�~*-Đ�a�	>Ti5�:CE>'trØ���R���T�_�dٗ����?"<A_T`6�e�|;�T)V�t��#�pe,��%a� &C7���)i�?�c_0��m=]�Ix��n�Hy��!Z�%��|��Er:w[��е���� �ģ���
�y'#G��|��7�9ϡ�v�ɗ����4�����P���C�w�i�s�ݥ�i(l��$T�`�I,O
��A�2���E���'�n���v�
�gbrp$J��g��x�w۸���c���J­e梁��y� ��o{�����qx��/ᰲ�����-��I��̴f���7B����rsu�߁��D�A�ԡm��k�z����wٮ�|k_ �^	�H`����nt�4k�4kTMs��
K>I�QV�Loky:�S'LU
��ץ��c�쥋���m��M�.�^^X�_���z�	C�D����&IL�3�VcP��P>ە���Lw����M�g�<�����fu��4m�5h2��v���^ۦ�����n�/�_�c���W���,�E���-�m��@f^����&��pQ̱=]ާ�@��
L����V�4�b�,��7���Xe�(Iv5���ZXU����*ƴP�@ܞ��Wd�$ZX��`���o���n%��IX�?�l�۞S�����~��mSD���h��$�� 'X<z$?��
�U[y$𱪭���/�j���D�ౚ���nZ>�1Կw�@EwO��`-qL{�%��a�[�)��*��N:Y����r=䕳qʤ8=�Ȣ0�C�
*��h����i&>���%P���=\�ͼ��Q����*թ;���vc���l�{K�m�%�����RdT�w�ǒ��܎5F�=�+w=%ҽ;w�R�����Uq� ��K��T)��,����5��׿͝]VƇ,��<�:+�D����-P�>͋#<�D�Lw�����ز%�Rx_f	�)to�%C��\|6'C�`�m/�F����5�X��x�P���B�k��Ʌ��,���]�ű�+`x�QheG�큸OQ&�+J�ťǍХDoYo8���f�D��fxq�����M��7D�3��Ȇk����K�g���C����!��j+�V{_��ۯ��۟C���y��(�I���Gv ���2m�?H���'��|�>34�������/�%=�S�uw!�j�	�F*N˧��#��j_�ȽTI�>6�� 5��^����Øv\[�$�>	����������lL���g��G��Xs�glJ��$���ʧa���*ť(a��JiJ���ȭz:M���h��tY��=M�h~X]��q�A�J�v��s��զb��oG��1���$a%�pr��帼�k������#c��M��Ƽ�.ƅ�U��\�r�c��k:R>��+��z-�z�؜^�����Fg���f�B�	�����i����\C'��E%�P���>��qB90����!�����Ĝ�|c�k72�]h������ͻG�vu����`C�-�') �;����.آ"$�ț�3���zQb������/�Y��G�H�.K�w=bj�Ӧ��CupS�����.���A��c���5��Ldd�Eo���hi�)��#nTM���G�6岐�	�RHY�Q��U��kzD=2��G���?:|!�G��m	w���.�q̦
��Kc�A2��	Q���F�/�lJ?��87��N��^j�P	���L��q��b9^����/��tCp�q㿬.c�-1�gɤ����q�;��3���uY�-N�w�">B~)�M�L4��As����fncwE �2���B�a�
���Pbv_-��k6��<i[�"��c4�/Y���ΎO<�5\�	]�h"�yѐA�*����h��e�ʢz�����:��*�)�7���,���Y�@ ���&xoo�#>W��O� bu��F�3���Wn�p6ے)[8Z�9�8"�*��˳��2�Z+d���`��<4�/|^Q�Kq��7�1��	�������'�x�7д��$u�r0Ed�cp��}���%Q�go�kcW	'q�!���/9����Q�F7X.N��7��t�}��b>����!-@�j@TZH����t_7��!I�h��fWV����-dA|�b�5ߐ���q�`�
*�����W;ļ�z*�%���/��]��ʾ艪6�����U�9Qi�3��Z?}��!Tz�Jhע9z��K
���t/Eh؅�L�C��P�ZB|�	O��ɶ�7҄ˢ�N��Kg_�E�O�/=ܲ|�kS�tT=Hm�"*{_�9�{]��gKc�k��U�v��6L [��D}(���,�܇V�����qfGu	T��9z��\�ccK��1��V�xP�9�����ڻ®&zEFw�)�MF�n��R�1�� �f�V��ɀ�z��+���Yso���{�eπkFK�d�O�{���ɺ�Xܪt{�V�6>#tcx>q�������~��<ŧe�p�$�o�ͽg~�x+i��͎�'6�:'�f����څ���!M2˨4w9���譟-JA��At@�ˣ�!1n�O����DǠ��êK0��Ar��u���mkx�$�A���p��wѐ�+�#���H R�h��,�'�(e���C��~*�f�|}�y�8 �ڟ ��0�IX��w�Vaoo�G�r�(V�03VAS�������*�j�B{��||0yr=),Y�G0��#�[f�m0�~ �41g�F��8�75��7�Ji��R SՁ37��l����i�X��$X1居盆��>l���.����Rݷ"[Ǜ0�`����������ԳV�@K�>b�V���.���E?x���~����u/��8Ց���ОI�1b��
 0zF���]�UW�!�;~�y���:?>֍�Q"M�E�B��sg!�/ުů�t��M"w�q�\�bB�ݿ�dO/4N%�im>FMӼ`�v4���cw�����Ä�~��_0���3�Hzje�U8�Ho3�����mq,�-��M'ˍa��R�X
�@��� �T��9i�Zg_��U�vӴ�D ��SD\L�&oO�������$�E냊l��=�>��Mt��]�v̉$�O����Ď�≋Z�\j���� 
���Ǽ%sq5�Ц����/I�sNd��J�v'������Ӏ|vg�r������=�,z���0l�U}�j�pW��꾇�Y�/1Yx?�>��О
�#��X���k�@Xm,��2�-�EŎ�R��w���1~+�/�1��'|E�A��3�FJ�f2h��I��j���Q��d I��J�)�G
8m�f�����뛄��x'��|	{{͓l�[�l�.>�=�έn-�߰z]�V/d�]3����žh
:���7Zqڻm" ������Am�b�~O�0�g2�^���^����<|*�ļ����މ���,�A<���]s/X>��4Ȫʸ���080*D�3V��(�;0�J~y�-��b��F§��W`��671��q3�'����,���:�@%�P��~����ѡ�}����������X�l7�����X�7@��V{j�Ǯ�s�EVu�F���Z�5�Wk�<�ד��O.A˃F��4u�{���:��W���^֗J+�Hk����#�ȝ����nR�4���?�Ťaà�6�_��um�\�Li�C(a�9J�������58��Ir�;�~\2��K�<U$��~Q�ڱ�omS��lO�x%�u�TX��v�V�����;�B�rb��YDg�ċ03b�u{փ�mV1��E:��7�9��;6B��=TU��ؒJ�e���#���EK���{껋g�n[p�R���!����6<=4I$9��6{]��6��k5�"Pڻ�������m�23�u�ۤg$F������R��<:�u�^q���g[���������R*Bfe�R�T��
+H"��wa�٘��ս��d��I7�ǽO!4�]$#xx��v�^��L��X3-;hø�|�W��s�(��>���&�)�d2�B�}�<�s�oCV�Z��{�R������̂_E���0ذw���~9�%+�6�{ZN8����-c|��U])(���8B�(n{��� �M���0/�=�����'n�6�>���|�1��U1���u���E�@7<�S�)G��2�6C���,s�˘�M�8֙��)fK�a�=_��	�I�`^(��1��y(�+E���S7�U,E\1kC��h{F-F$)&����L�1h��by��T�#7�#¯?zk]~���`�������Ww�{I�Gf']�!;.[��~k�dk�[��+�x�6��u���:)�$������Lx�,�6�	�q�c:0!uz�}�fs�#R%2�>Y5c�K�sS���M��䨿�����#�b�r��;�b����AA�[��r�Dӽ���Y0�/JL7'~i��a-�W�6B��цU�g_�靵x��?\VR�؇2s��j���D{D&�a����H��RhҀ/Pbjѽ��΄	��[Ժ���3ż�n҂8�F���c6��Q�8��ˈ����fu��qWI���ߏ�X�&�� �aSH�0�sz�F�2��hZ��UٗvO<|5�|
�Ð�R:���1�{EK����$��3�ϳZ��+T&FT����6'�i"rS�OHU�sX�c�A��6�$CұK�v��Q�;4��@��A5����Q������*�,-a����`V��o�HR��ѭ�<J�,e<ŧu����xm&�5~X��@��� ������=������B��l��~?���?g9J\�l0���!���-u%����0����D���PRԭ����= �J��h���E�����쭣E&/Ư7 ����Q�W6jy�Ͳ��`�����=�[T��+��9�U��)3.��XDJ�c����B��e�c��i3�9�U���b#�~D�;�ľ`�-:��ȅ�"| ���S�F.���	��pP60 �}��FHr��2����^�/�����Eq���=�<Y�[�0��#�.��gi�E���޹�-�?�t%��p�@�~My;���Yp�-�R8R? �6޼!}!�" �)�Tq�:�s��3杖�#����Qr��~�h�;\@��K�.��ANT�fE���h�?�g/}��p$����zxh��r{�5������B�=T#%^6�h���~�O`��ҵv-JpVR2֒gGK8�1`4[HJ�G驭�x��E]X����3�}rA����3S��|��nwJ�@�6Q_�� �Н�~�c�(�uYަˠ`?�^��F���5]�8}z���[�6����i���� .M̗I�kWKB�/�TAǆ��U�U�eŰ1�-��S�PY�;�%�f�����h��b�6B.
:D�!,�t~�3�]�����f���)e�)�1�� �u�ř,����Σp��~�<�ـ�U8u]��w �J���ⲥ���c9:V$����J��Tj?@�19��[��n���P	�ѡ�ę0P��M-��3�^TU��X�F�F��[�A+�=uс����z)F�`ҥSgkڱ�EwY�Z﹧ע� "o�jt�i�Q˚��o�k�w��]�vBg�����#�����Q����-Q��H]8�S���h����l��Y�W��#얉s�����@�fs��|4�ٱ�fp��)/�.��G+��gvwĻ�`K��x_�\ą��X_f{8���O��i�ss���`�C)��+]�&ހ}ק�=�	[ ]$M��QP)N.)���fq��jP���m���<�a�G.w�ʓ���fThI-x������� ��?35q��l
1���W�]7��.b����ͮvm#z�>���4��I5L����gVE��-eB�X>m���D�89��>�젋D�M	 �zDs:_����-멋w/��*�#<�Y�?>s�,��FDZ<~�P���P��6�z����i�R�}�%��(��iX�=a��'���ꗙ$;���}�3 b�҆Q/>�=/K|e��\nqS2�$�f<º1�N�|07��l��  |��z��uڊ�6���F�e�Cot�7	ˑ�¶-7[��%�)$`���Z�N�
�]��E�/\�t�b�N-�%�\�`��>�.�ᣂ���ZO6��}V �`o5�Y:�z��jп���Mm�]���y�M����o�yY���ű���h~1Gf^��/�v�w*Ko/� �5��D���x�6Z:���\��;�#��Ju*�f��N����6�:*7WP���}fc;����0�Ï���6'}u��~y��%�M}/��)gL�`�D�.q�ԄUq(��ǚDo5�Y�k���8:��MJ���~+����}d��Dם�1l9�ȫ�[�*T��z�ǇYiK�-���|vӖ�`���U��Loh8O� 8�1"����/��%oTC=p6N`��`K3g����\E.@���i��k9��N(�JY�K͋Ԑ�� �JЖ����"š�������r���;� ��c�J��t(�����Ɠ�?���o�G��Zf$l�eē��~ۧz�����I��G�0a�����[�E�Ki�>�nv&z\����E����"*���1��7Oz`2ֺ�b��=C"�a�I� nPJ�Wu�^�>T��j��xG�-�n2��L�{˳FU�ā�/l����s�pf��>u�M{�4�����r�jC��ݬI̾�=)���u�6/
q���M{T*#���|��l�Ы�pc@��7ӣL5�u0�>�(��^���{���U��Mhp����xs�*��
��wi�
��_2[����Qr���=L$.EA[Jꨭ�4pP�U�F��蕢2v)&��8�H��! �ly{�7D1S�@�T?�k��oԯ)f���ዙ)�6���B>�S]:p`5�J�M�Y��Ow��� ��}v�/B�	��{���nث�|�;=|�� X3��Ґ��kAl.���f!�y.�t�k�+D�6��_sI�hC�ft>�@����ȼe��/�O@T?{gQ'
��Pn�0q<e�.�����#W���Y͓��#
V��;!Z+���X��K��?��8p���j��O�F�{ʹ{F�J3�D�b+pPZ$�|�g<�7ɠ�S�L�{c�<���:��9�c�5<PV0�D:��nd�y�	߄�L�	��6�-���|4z`l7V���>���2�U����?7����.qJ��hs��+�m�Q��3��(q�q3I�Kv��L�F���x�(���Ͼ,��z�-_%���a��?zڬL���$=q=�dU�Z��D�]J��e������n���>5d�}+����"z����e������D�n��/ua�7�70�]��Z���{�'̓!3n�[�i�>��cj�c�g�S�N�GS*�22).�n.NJ��"�j�mR�|.A0B�8�]�4��k�}���&���7& ��a
V�Pl-�GWH��$���Ci������V�^3��	w�ກ\�c��j$)��,���	���`5��.L3o~��S:�;9�iccq�o��=��sX�W��N+*cg���]�c�#K����^6{���xq���6�p��X�Qk�����`�=J��V	��lP_b:*���(�
B}�=:��-�}�gf|�,�=�x����ҋotS�܍?��Є�y��>����K,3��AA0��s#�`��Y1��h���$�ͨZ�' �W����>��azx�r%J�N{4���bx����,u�T�;Ϻ��E��ak`��ȢXa�'�p�ݾ�E���B��+=�\` fV������nu�*O,kŬ�	�ْ�?v�MR���K�� �5�ޕ�D�;[aX�jKx�Z�;�[�1��%+)ld#�Wc-Y��I���VL�T�k���4�7�fB��E�l+X�����I��22~��x��7�F��	TJ��C���h$��g�&@�f���G,��i����-�u���oVx�1d�|�٨�Q����@��k�F�ݧgr�W��>ck�t=�ro�^�B�$��$ظ�|]�B���SY6�r.�����*9tʅ�ץt�NA��?��Q��[�Y�2��� v�"5)d~��)�ɻN��7��{�Huһ�.8Ə�u��PF2�/g��F4?DOB��(iˇ�4�j��b���DP�`�ʀ	d6pT���j���8&X��<��.� 7 a���v�h[�oO^=A5����ʥ#�xQ�iKs������m�%�b��P���EոKj6��i��T��q��F�3#*մ�'�ʠ���ƑM���D\��V�q	���_p������#�zA�s�T����6N�>��p�@r������c�]C=���"�u��A$	�"�~�P���[" m��L�$94 :@9�e��fj@"�6�][���T�&v3QW�˼ʧ疯�{�h��"EQ�����*�4�D�ؤW�^�s��w�	��x���4?�yҮ��W��p�����ǹTRNc �F;@��yͩ�[Dy�5��D3۟& �f|t�x��LhKi�qN��9N'��q�sRd��1�e`e�@K2���@����Gd�F3t��N�Ŵx֘?�ٕ�oY}H����oYC��J��:8Uf��ai]�P�t��U~Ҧ�s�!3B��g�0"ЉZ�����+j�[8S��~�z�m��⬪>I��o1�7댫�y����&�?SX'�8}�;_n/,�=E7�,�q�;+e����B.�/HU�J��{[?����fx�@Vh�����+�
U��*H���!��LMCos����z�<z$O�h��<E�@�X��,	=9��=���8|>��v m+Y˥<��}�W��rr ȗD��e��^��\i�-^ײ�Is]�E{�o�>jZ?��w �_�˦J�}�� )��X��l�!����;��{����-�W]�Z�A*z�̒��?��t������>����ƎOY&2vTEQ&�S�G�m!�؉������!�-�`x�E�_��~�`ͤ���J���}J���Ū�����V3�ԙ��kFu=�p� �P�gA>�{W�Òa���,��)�k��� ;�dh)V� 턚�� ��32,����H��@��W#�����c>Q,����x�-�K�#�FNXi޳ɐ�UT0ɟu�6�^�+�'��M`����l�����F��N�X�lq�?Eַ2��^@l�ʳ�%B� !X�-��,S$�w�������s�|>Ur�|�L~�һI�>�"�ȼ��z�������$�6]�ʨI�*!V�@��t��z3�
� ���/Q�K ~�N�0g�Yu}�BL�h��)M��&��-2�J�+��Kz(��n����g��CV���Y�*��`S0M����QvG掶G��x zK���؎�iPXa���E�����#�8����Y_-�X���SP��JL�T*�!�W]������C(1ك��4��o2�d̯ߊ3^�ʝ���3�w"����j�E��1'WT�#t��D���>��§Û���}$(��#9x�����f:̮�����.� iT\yڋS?Y�9)h�E�by;묬��t�=�|��������@�N^�� ?��9�{��R�m�&��,��4Ӳ�a���"O[��-��)]��[�W�d��J��Am��{I��{׹	ܶZ��M�ҳ���	�@���^��(�jg�i~���=�U�Q�'V�`T?q�Z8�W��Չ��G�ԥ��G�P��*X��~�����	[�
�ҁ߿(;\L"�h��}:�� �>Ǟ����<��"��L=�]a�R���<IA��LeA�>��ð�}�
�[���Y���B֛�|w���X7\�F]Z�{}��e"\��e��"�ff�B��EB�5�s�*
�
٘�uo� �Z�Я/�8ѳ;z�G#����*B0A��X�6�k*�)�/�ג�q#���4�Dd��P���>�oi���(E�"�14����lw��o�;�����矙_p�F���i��2M�'��f'�QQ��"���p��0�{��E�I��U���l)��	�է���os��g��wUu��x_��mS	�����C�2K�r���X�����~C~�!���!��9�&�$!������^f��&�����I)�E΂<"�]�#N,y"[_a�`�@Ȁ�(u�b8c�L��@솊���9<��7�M�b(��Җn��0��G0�l�~J/�Q&��}U}d���^ss#���8�{麗_S?ԾkӔ[_	�Ġ{ܶ8�"���^���<��]�c��*v�_L���a���'���
-|]��W��l�)�W=�wyz$�7��,�d����,�~{HK#n��ǰi��ir&^� H�49a�Nd4��M}�9�huB���Ąy�`Բ��9��g�g3fa=0ۣ��e�?����`/�o9�W�U5I��W'�ĝ:K��{uQ�d����-�@�4T֨��zYQ�\? ���09��'�z�pMJ���o�u�P������㇕�e-��eZ�w���qI��Q���?���I���$�).�#,�&)�o��%:�fpxY��gD\E��7C#/N�|�ԑ\Ǘ=V�#�V��s�2�� G^��!�,k'�f�dJ����(0d}�x1����Q����
��K�$���s��^Y90sa�����5�Vn�j2A�ǀ���<�_��&���x#^�f$:S:<%��� ��!ߢ�Y`�G"�VV�Z�7vI.T򿩟�g�N{L���|����<~�)��'�%�~��VO�/����X\���o(Qڳߜ4}{����q'�F
���}�JN�q�4�\g�m⭁�͐"P��3���cY8��(*/��w�z�m.˗���)x]��h�a��Y��M�c*?R�&Ξ�(Q�I�̝k���wz:&@"i��`���K9~�vU�/�,H�j�3�UD����՟[�K�J�Xw#������-+����1x�U�F���?s��ڟ?��_���:�.�]#$k�^��^By!�zpf�j�L,�W�p�Ry#N�[�"�h2���Y}r�a[���ѫ�c7ٙM�
]@~x��,���H��ꂀ�>��v�����,nZr�]���1�THnx�Ӏ��\"�M ��2�!����BX�=a��Ѭ�q��gX�̓#�q㯿ڽ�OD,��J�����(��]٘��8����|�#iL(@D
Ql����~�QN>-�����zoj���I�́�s�~��s�}@��}Ft��ۑu1�e�2y*��80�Ǿ�5���[��|�U�c��Y��oaq`���s����X_�����ʊa��M:q���9�7�+u,�>��s��{	�2�����ߠ݇Tq��uk���.J��aKXx_9�������v�8�O92ec!�I��ӒA_Vwu��lj"�D��&-���!2l��B����GM|S2t�D�&&�!���<��LΧ"��d@N�ZY�
8�	�}��]�
�m�䠲z������A9�ԖH̴Ee�UiH����\l���U߼�&ӋD#)[/�?h���NחqxG�����'��]7G.�Zpeeu�O3L���F����gA˂&��h�
�;U��Bܛ(P��@�$�:*#R����R��Ԋ{�}Z L<,�!2P��S�07.Q(�L'��=U"CY���d�s/����&�B����A���R�A�����)J��l�,��;Ľ��`d�U6�I��t���ehۍ��n� HO�	������D�u)$��x�d���6�G�����_h����![p�����#9_�[eb����z|(|�g��6�WI$x6�6�����-	hmt�� �{)G֭6��G\F��@A����������y��8�}�n�� �w`��>����|ص�Q.��Vu��C	���?�3̙b�%�|,P�/���/��TD�,����ۄ�����D��ݖ�.I�  ���u��`ʜ�J�E[/X3�s�����.���~N	�S�����;����o�nk[��i�'q`x=���?�����Y� �yy#��?,OM) ���QO^L/�C��� ����H��_���ЌP��	�B���5c3y���Ѯ�hEU7���{6Xg�:	Nc�E��|�~"��m��_��J眗�-Ð�)2�	6Qؑ�NCt�I�V引4�,�˯�����q�s]{������7�hF�qW�qqڗ��ؗ�a�QK��r�/��4y�i�}@<���N|��MD��Pv�����:�^\E�k�[?ߜ�9�E+���#Y&�x#ГR�n�F�OE���j�~�r�vZ��ܾ��f�%7�Zp�`�o[nO��*Ѿ1�䏖"�4�����-�]s�Duh*,ji���e��p�qJ=AEe���=���n�o��۷�XY�P�ԩ:a�Q����'�x��U�OD��8[{{��9L�m���N�X�b�JC��t5#L�v�ؓ�k>��G�z�a8͒�:n�D�2��D�����7����Dl����KT�|�����"Ɠq��3�=0����g2���N�ܛ�԰���q �X��i "*�xC�
+�	w��._m�!^�l�8�0)l��-�0XNdۙ�B� ذ�<�Z~b.6���0A�~���.����ny��uhf_ ��ێe�Z��ذ�6IO��]�أ�q��#��,i0����/��m8A�Kb4C�$����|՜tt�S!=.���@7�O͆u<�3��wK�h�;�eI���ڬ��l�X�������|�v�b:$�+�'���c���KF�I�܈���}�d����W�mm� =QK��L����s���v��0+���rG�"�r]ó�g
@/)�+.�e�4lm^���*��vh�M|�:Ձ�VP�R��:���X@��0ΉU�V#B-
&�[C:BfE�5.��F|2__>麻`�Z��/ۑ�f��]�)�����&�]�pg%�F���N$���Yk�bP]�ꊛH��lӏ���w�	�銴�?�`��|��MaB%ڠo�Zˍ�kl�iP�E���8�Ҷ�췖�_̾�����g��Rm�Hk�bT�F�x��@��Yj�W���+ν4"BF[#�1ډˑ����[�T]���H��!u�uࠡas���I�֘�����q%����04}R��b�ՌSZ9̫��P�!�+�,WՐ�^g��2.���k���/�/޸ns��y�D���Wq����?�G���G��������׬`��]-�JF�����J�����b %��nhbE�H�IH 4W;���S�2��?�;[́�0ۭD�����$n�LɿS���g���<��ԅI�/���DM����{k��y0U�'�DX�0:Ю�}�Bx������Lm�[;�,�CM�i�[�P�Tk�%$�w@�6�\�����ʤip����iN�K�	���Ci�3��M��}p��.��d(
��}"���?h��b��pl-�׍�La�FMG~`5tw�=���u��_i�Br׹����A��ɾ��V��Jt*O�l�I���bn�aZMӟ���[���|�=Mk���W�!� Ve�˚#@S���x�:^U*��1��d�U�N!�@;I\ ��v�z+�Z[Z�����rx�n��=�E�&Ԅ���Y�u7G��$k�>B5e �ӖQ Y#���W���9��1y7ٽ�B��"yB��)x�TN�S�&�myT�ߙVX�Th�>�~S0���<��� �@�b������4�[�x��m�N.y���D@�	�շ�� A��c#O㛈�=�g K�2c W���a���c�����p�č�a�L)�k@z%ɯ��=�x�I�d�o>	�ްT]��ѿ�Z� ��30+�j�b��p�-�Y���T	��{3��`r��.�*��R]1*�D�_'�q*L,O�[71�����'��~�(�Y7�s���+�*�V&��hO�_��u�w뉕��K��C� s(u?L}����3���>�X��.��^��w:u�gXK��yo��������22e�@0u@��Wt�2�tJc0\����3��KV��d ��c#V�Xb03#��S/~�i��s"�&�rZ���ZOO!� tcN������߷��b+�Q�2�6�\RY9:,ٖPA���V�a]�G����i߮�P\�Ѝ��]���Z�S�.ݟ=_�]g,��y��<)���J���,wm���/�g��:�v	�[u��_�5pgD�P�mLV��K�f�����3���M���{gL Ќ��S<5!�k���9�0Oaܞ�up�2�=@�CW�p�.ō�����啨@�r�BXB�:�:�࿦64�1y`���Bm�]sʖ~�6s^$@� ��Hqp=����2���ޜ�?�Ȩ���5�ߺd�i
�Ξ��dT]�4�&�\��</b ��m)�N��5X���
H�f��j\-F-X2�G����Z�KW��G����1&�e�)BU��b�5jWf��̎�X���n����Jw'�t����6��N��=dֳ`�A�otS�|��6��e$7�1"�hwO��ް�������x_��l�+a�[5�]]���(M`v^�ؗ�2ܓ��A�`�nI�6��)��PGK<}���a,�@7�<�J��Z��>6��)
��*Q!r+qs��W!����� <N�T�~Wa��Dn��*]��4�U�ᕨ5�8 � AMk�CA���o�`�O���tK���%hu
�<���g�T6o��IF@��/�1��@���;_�JO6���ޞoe¿���dmu�D�Q�l��]H#��X�����S7jep�����4�P]G����|�O�f3��^����p��lP^��@�:�W;���N�i�7k;6V����_ӧ�r����  }��x&PyX���X	/�?�`��j�����z2��AJ�b\2������\4f�j$iS�e��8$��-ِ�Z�P�Ԡ���{��Q������!:M�ŧ�6z=�w?Zk��qY�V˙�9r=[.�Gf����yb/���~��fo�}��2��>i��=��T��7g���|{=�X�]�A�'^�e�6�s� s�{��w�����/��̊�V��!h/���ޯ�n��%���u3�{���^/�G0<\h���g0�f�%�6F���ޏl��H���Ө���v௙�~�, t�:�u��1��O���_�|I}���N��-�E}��b I���I�-|t��x�7U{f@�peML�/G�2�N�\�N�E�B��rqL�%h~h�!�8�=�-e`�����<0�N�IF�L�9��@�5�ۙJ`���IQ�1��0�¼3�ڛ�2l�R��F���س2�2�E�!��5��>O��{Y����ђ��ü}� �-���<�Ng;�S���w<:�|���!�l��U\��%Ν��޲G�j���aL~���V�{���_T.��A'g C�£��"�6Z���p���D'�0⬊r��˔�;�v=�u���(O�g+�$8t7Vgقͻ+��2�5H����)�M�tD�G�1u�I���p�hM��S��1DF�4������F��B�����̌�3�~hnCWfd+�~+�����'Z�>���^��y���#���1.\60Y��BC�eF����o6�d�KW�����@�9i�K��E�0�q�N�׍�Q՟�:�,R�^&~�i��>��w]M��[�����6:D+{e���'y����K0�򋅌rg�$��r�(�6��a��X/�ݿ`ս� ylo���q©󙄋�Ys� q��W�,9t�b�5;�8���4z����k�Zn�h]�;��x�z㎪wn��λ�[�*��:��٫8u|��q��	��� (�_.�Y�^�Y:�A�KBaXį���^�������=1�6ӃT@\�0Z��-�Ԕg`��cb��B!iEO^�q0s���Ի}��ű��9�dvxzpcXڐ3t��pNgvv(��B��4 U򀛺^9���IKP�"��?�46(بko�Mk�p���KTnU���Ƨ��.+c�j1��'�O���4����M0�d�R��\B�Z�����^���!��&"��H�#���r�P3�A<h_��H��MS6hM�=��Q������8*���_�2�V������I$F�};��Sq +��Il�ȡPk����Q�u�T��<um�e��B�n��}�����Fn��eX��7h�vj�Z�?'�͘��s|�L�P�d0�7��U�<"�}�r�<�L����� ����R���	�c�����uB�e�1�|tb �S��E�]�[�0Y
K;
*�[ƈY� ���3��Xw�6Q�2B�m��*ǣ��j�d��{k�$4���͸q2E�Q�>���G�(�8D�/Bi��F���jpm�Rb��/N�n]��Bn�ւ������+Ec�*�q���֊����i�fF,Kĩ,x������9�fmџ���?�5������2l��]}7�"���V��I��%�����/�4Y�Ţ�AL�C�
�ۆ]�I�9M�!��	�ne�0�����? �%ՖF��V��1����\y���v �>��7�o1�g.�<�5{GX9��.�R���]E�L�%37�w��F%��W�#��~k�����8���p�l�1T�uf�VV�����(	l+�L3Rl$mk������������f�p^���R4WaX�	�;�Y�Y�ʾ.L�0̽�V��2|t�.D�q٬ŕ�ց^Zc^���|J�����F����A��A������@�0=a������^�aտ8�()	��s� ?RqW�8�+�f(��3k8��Dj�T��nR6Ujm�����to�3��)ʞ =5^��!?sx35?���P��h�7Jc�Y%����Dd��h���ܚX*J���[tMqj`+�����Vx��k��?�6rj֫�:?V2\ԴV���I�Zw��(�4��B ����5��:�LېY�b(��\.N$�;���y�����*y�+&qd!#�g���쫗�T��
j�~!kx��{��	*�������lI�)�ϺI����?�!DSHM_���i"�sad�h����U�=�{^S��D�bw���܀��+,B���;'�9�E߮<��ז���PR�㺒o��2L`6o3|~�(3rX1P.��eΣw�񽃙؈=Ƹ�i�s���wI�Cq��
�4�����.���o�:H	9��9�c:W�[=a��"���C�=���*��{~�zZ₰1顛�,E�강��)]X(��|M��s��=��-n���-_N]MS��o�� #@�G�f��XS�fhʚ̖()GP�e�p4�%͉�%�n�)�R�{ɛ��w鱇�_����0d#�T��n�~��)�sN�;�0V���b��d�%�l�`斋VTm�������wYm�<f	KQ&瑘r��VF�\��[:?�_p�^%�������WF���y!:ț�{ʝ� ����u�*5)�h���|���ߴZ+G����z��'� �^ A�ʡFP;�HtT���r��M��JtO��&�d�4�T�D=�F{u,�O�㋏����f��l���WC|�H:���UG�_���P��SV~�~��.da�s;2���I�w�
;E.Ǫ`���3�K�P~dm卢Lp��*���nM.�}.߯Og���t��Q�'w��������YV��]��x!uE%�
ڍ���Pfn�!���5t�ݽR�`:�Y�4+�;������2/�P<!Ǜ+M�a�j
�Ώ��O�L�:��X�!D���J?�L�?��N��ŉݼ6��G�9fg~��9�Z�//4�t>=����SfY��jH���I���̨�<����sW5�g-w�/��Jk���Tt+W�2�Ԍy���7[��D�xb�W�Tތʯɽ�63ZU4�E%�=�O��Xl���<N�|s=�e�a5��"��e���������v��d-iι�xJ��B�aTYՎYW/���ۈފ�> �?� /W��yQ�FE]jX��䞟� ���X(*r����Y�	bJ6N�8`�&�wT�-Sv��.^S�$��A�:΂v	�6i��43����	>��� !�	�m޼=�t.��_)=�LZŏt�ٹg6j�&U�6�*
�G�	�p�E!a=���р�/ � "����*%��-�M��'�)#JOt��Y8�H����;i�h�N/d��Q`=1"�q&�k��Pn�cơ���lHװ�μ"B5p�`��Ac}�zA(V&P��i���
��gNj���u矏;&9��u��$��L�T�^���R(�ϑ�{�a� E!ߌ��:���� �߿)s:�!�F��/��<���:��j�����M���:odW�Ů�ˏXߗ�'�U�8��WE���vxr��ڲ||��%�[�Ԫ!�Ew�+����jG�1���9W4	�����i����SfB�$�c�k��`�)R��J��P��R�<��:����8�p_��_��ÒS��D}=�^���	�?�� i���Q��I�G���n	�e��>7���RV�'��� /5���,�&d�v���ˀ�E��cv.�p�����ڣ���
ʘ�7����좗4-߹(nk	A_��;~p��#"�]i��O�5A%�>���\�������j��Z�Hǽ��߄@$*)/�cԪs(�N���t���Zu��J�x�DGkR� ���|�'ˠ���C�q��Ϗ8V]s����CP�WC�����4��ʳ�𣣰�����^��q�%םؓv?:y��J��0�H��t4������Ǵ{ZjH��lBR�̪�P��hD�d��V��F7W�w�pYiQY������V��0e���B�
�5��F<��� �4�ͣ�N����?;�J�R�
ibǵc��K�����`0p�Y��Pa�����Nx�eHmR���ێ�2L���k�޴�2=+���y෨ŏ9���9�����=�ģ�\?��t"�r��x�H*T���P_{�u�$��O[�XbH��Ad�v�p�[����B"�g�(FpQkT|�3��
�(M�ӆz����쳄�ˆ�� ��pC���ۜ��D�%dLx�~�Q`�Cy� #��Љ'jwW ��K@�JP��&�eJ�vm�.�\����';��kA�12d��c�{����Es,�g2��o��>.��Ē+.gqlb����o��Pt�V��ˬ�b��� ���G�=d��G�/�����q)����-'�K	��-"�ړ6b��#�@��;'�"�*��h-_�c�f�]`N!������{��|~�?7`M?ϞC�����ݨ�!�Q�ݤ� t�e%��^�ڴ��mJ�o�]�W-g�ˋ�(�~/F/i�@y�P��A@=�El�A��M7��2��ZٳU{d%V�`����rҳ���ӵ��&�Zs2�X��i!�^@��JQ02��ZO���b,;3����F*���W�S��S�����ޢ`��f�
��%�;��D��jسm�/0<ʪ��`���ƖI3cU��5o}WC�����Z���+-���@�S��^�Va�F �Ɔ�1S��>�)���
�{&�S�r��BҢ�����
�(�N������])���%�j8�u}�KV&��Rrpt����^�vҘs����h��6,v����g=`E�h��o�u���H����4W�n���^��:��j� ����pn<�x��R�gk�_�!�N�"x(�� }/��O4����h��-�� � "湥Ƿ��}#�?���:�(�ܲR��S�!vrvJF>���zP"�2���R'u�d��0��R7��;\�=���$7�zTLu�<�r��\�4�&�+(f�D=J�4���F��p>���d��w�'�ݙ�eo��Q��~�V.�����I6��9��ۚ�`�]��"`J�됺����hL/]x�~ʖYޜ� ��#�yČ A�v��%4����[�w����(zy婎�mWr� �3�{>KS�}Ե"��>]a?X	�
�dB���ч����J���""?��4&
>���a0���7-Ŭ�k6�����$k�nݙ�ֽ |s&o�|�����Oə��o=�[?X'�h�nߓ$-s�I�꧁x���{1�����\A�0�]�ԑ(Nh,m��΄�raeZ�l~h���Ej�YYS�Ԭ_̆��'y	�("Z�etp;�'D�C�1�^�6�m�	 ��EЯ�	�u����KNB�,&lK��Pz_m��0l��u�ֱ�sS5	b��y�S�V]غc乵3� �((�;ѻk�r2���ÈK�w�KR �%=	8�2���n��+��eR�=̙�<�-EȊ�Y5cѽ\]�9�2��'k�^��_"i���0�:feA_.��#���H�n���	�RŰ��O��΃J`rL<�)�o����e~l���VH� ����L�^q;L.����t��P�bPM,<\[4�/���|�:�!���A��Xmb���x�������׻"����'��	t-����ϛr�#@�P��������@�r�Xq��	�Rg���2���"r�
�?�g��U���i������]	����2�fRO�d�]�5ʽ�����W�3ˬR���+n�k��o�������æi�	����7�PE�9Y:|=��0b%<ik
`�dj4|wNzC�]@1�>�=���i#{� 8J�NUH-m�A������B�'˝������l�4�P�P��Ԓp�+��zޑ�b��L��CY{�xr ���$Ivi����.��2��n��ќ��E��;Cs��TL��ϰ��U@����*;Q^
}��A�s'�۸�y�q�Ͱ�l��m9�S ��;�	d����u��~q_�9)zN;?��/b������M{�薕��]���cn��m��4I�����e�[��p:�:��kP����3hD��t�2;na�V:5�n}�s��V���G�蟫Tmt����i����r�Wa~_�+�:��@��"q�r�R��c��8��4췃��)���;KZ{s�3J/dҾ��>xE�s�T� z(��!5(}��'y۟@BjX#!;�\,{�%5�<������0;�P�Ih!vݬ�M��8�#{�ģ�6�w�����-�W�Bs�z�a���rbk쀼�C����j��G�dσ!�;'0��L������ p�Z�ˮ|~���|��la_%,��ḟ+�[�8K!, :5����0�1)n"��_���|�t~ԇBb=�/��X*W����>���6�*��WU�{By�l���4��!���@��]��A㼑�����aX�#����zF7����<�]�b����,�	F���/�ɋn6	k6����6���rq�pm��p�ƈjb�r�+�9Y�b�y�%v�iw�<$�m�Z�բ�g����5o�
ny��F*�{g���TX��R��!xz���8"�Ԥ@�/�Lkp�_�����x>�R��L�G�b���"��!��"���!=v�9�s��L���ry6;�o�(��d YP0�+H�osq��j������x}�o��h<Oa�#s���)ܞ=�R�'&��fc�J��	��OH\���<	�D��!3�nm�=�ǐ�6���������w��L�q�2NAZ0����ix�^�k�T2F�:���Y��2yX;2dg�����bv�5d���h�Wpפut�Z�� %�e�T*ll���S���詃 ��p�-��~T���&��K��@�^�K�n�c�@utv�S�೯%��%ӽ���&�]�������=R��TX;8�O��&i��)F�$�2�2�˻� ��/��c'�0ā(�hM%彧�*�-&���W�2�g�6 ����>�(��f�x��W����wv�ct$���N��-�j���D룎禟7��e��f������E+y-*��$c`԰��c�V>��Ej���I��K��.4O�[D���>A
a�,�O�M4K��	w��1�)���9aRsq�XCa��fPZ�<��G�lz�D�+�Z>x6EI�_�<�Š�7cc2/�;����qo)׌1)Q�S����#�����T�V�e��O$죋Q�5�<YV$B��ܕ���v�V_���tɅ$�s�:�pp�N�y��-�_��-'�Z�8u��E��6SE��ߏ���.�1"�ǂ35���K�K?vj"K�n}n�2[E�ע a���{�Ltث�eӵ��C�� 	��Z(Kdb�	��u=�鍊����o��R����zp���kTC��j�R�|$�����o%gӭV�d�Qٴ��tP3ʣ:֯5:�8���X��Ý|�6���G"҃C�gX� )uu;�/2�g(g�!���fh�'�Ueyw�P1�Uzt#HlH ��ތE=G`�>c[TU�T�ʷe0[�8*����u{��3�匓��̐|hw�5��lz�g6�C�*&� ��jH��}Y dDmߝ� T�ǡ��40PN�®��8'<�8{&�_~�3���tN�챐��K���:Ze�9�����m�5�yk1uܘ�q�o�����,�����u�ɬ�lβ!���o��ov�eA)��t%��K���LY���j�Ճ������}8�fy�8>kI�����?�$/;.'_�Ǿ� TF`����pWJs�q|�-��|i|�r��ֳ������Zтf��Q���I�-��_�U�QБ��KoR��� _��� fW��;��c���t
%��l��6�-Vk�2�c�c�Ì��Y�x�:��q:)RM�����0P��V��]�d#�K��������zu�bT�ʞ����eq�B�B�ʺD��#k"G~�A�� x��u1L�[��9���=j��ٲ��<��D ����-����%M�`[~�	��x|ІN����IH$�
1&�9|�r����Ƹϲ]v�rc�v_-j�lF���f���#m:+��#���n4�)�J��E����I�Bۮ�[��R�@2�t�Q�B�����z6�sj1����1��uJ�ِ4�:��T/j���_)@9u�dh���	�) �G�d��
�����2N.��i�����/��vNᒂ ���h� ���S�eV�O$�e��#,,�W{�����C׎�`� "o_���Aΐ�l�.���6�»Q���?,��.����s��Ϛ�+��#�%�o�O����ͫ��0��t�
x����$�z�9kLG+gI���_0���L�qo?%��gU���~�D|0�hZ�uv�J�(�5A��fB������(��mWg<��z���� @Âr���٫J2�^�*��1��4S��2����\M�]� � ߤ�[h�k}��8�i��O0j�vՏ�ۂ?�r�{s��V?͍��nx��,$?t(M�+#%�I��� �LP�M�6�҄����U�#,FhY�N̆g���8TW73�l>�X�a�}V���q9{�uP��ZN��ng���ʌ"��L�f0����d:_'�_��l������6���䇻��jv	�Ӎ��ދ�߃��yd��x4� �S��h<�>�?;�M[�w��8%%=C1S�����݋���,1a��s�����@G��!��x��N�T8h(��|�l�'�Lw�)s�V�Co�C�m�J�͜F���>G$��!�� N�,�J����b��df�j�L�g�(L�b�"�wM𝱟o�r��+���`A��D��Ӳ��4Q[WP����P�Mp|�Kb/�b�_��&{Z�}:����*�X���|�@���CX3%_S���WfNj4rӾH�-U�+F�9���v��� �6VNDE	�~ט�~b�0�o<�8�.��ofXz��+F�����A��I�-mBa4!�p̻��\�\�����\v���[r�q݃kT��P]q�'�f�������b�ePC��Ɛp������]�F���s���k
v"�K)~��q` ���HH,B���	�)�n}Ё��j�d\)ጠ�[�CCX?w������l��/��7��S�dy�q�D`:�ZC�9��x,�K��Q)�׃9Y�B)ǀ�8?�j�����^��;H�5����5��?�Z��a!N$J���,aX�Y�D��N���,y���4�uvi���7�� ��+y�ʼq�r+ޖ��ÍP��H@̈́�r4�H.<NVR\�m	/��`���[A������Qe'��Y��������e��/�~�r�<����I���-��}�Ufq�iRT�K�g���*L<�e������&�4��5z f�������Y���WA�렽� ���,�Ө�_H��y�����CB���h���'|�����N~�#Ĩ����9�&4ui��$�n�e$X*5Z,��g&.Jl��d�]�߇�|��zoiؚ��8�٭���:{��:��.0�Xx?��lP��|Y�F�<��I��0�_	k��#0�'��ç[K����,}3�q���|�5O<�R���z}��E�A<�Х�OB#�����{ �&�����ak�1�|��9L��e��T�T/p�OWb����cS�C��Y�+�4e�64{�d�c/��H���h|�]_������DiL�J�bi�>b�&b�%�{��/"�|l&�̂�[��G�+�Yt��!�ZX�������B�c?b�홎]G*ƛT?f­��Moi2���1���ϥУgb����RpL£R'�dߐ�2��xS�!�	ޤ(�͸�ڰ0���0��k�K�%���������d����V4�[j����t/Ύ�U���9I�d���E�}O�w՘)�ڐ`8�-�i�%DԸQ�6�揄����K��~�~>u�]V([�״ʢ�Ko���]l=�v����[���1��:�Ge�p�؀���[�22�w.��������v��6�W�\&%+�N<oMO�E�C�$b)�H��1�����	�~T�`iV���\�'L韤;\Y���4/B��#qo��Zͺ�B\A{�QCnz�p�0�6�V!�;*V!���s�)�֬UI���$��]M��s �URJW���nzV׷$ s'����WI0y_��Qx�I %� @�z�C�vN��⣩?�1�X�*��!m#��
�ޛ>Z%:��(�֓�8${�M����3�ڰ� ˖1���ޑ�~�R�;�ǽ� �'Ȕ#����J�
2�N5�;��C��������qZ�(�Ba���s�l ��Է�g���3��\��^�ª��:Z�׺Kٸ�Z0]�]?�S>�����{-\lr�����tf����I�+���6?(�tii0�W�<�� �K{�ox]/�a !ўA�g�~�m6��lZ.���|���U��L��u��>Hce����;�Y�A�{8����I?+����6�������_����J���$���/�$%6�BXn�N<�&d�c�l�%Mie��ʊ|�����Z�Q�L{J"THl�[zdo���C���ܤ�d��[�0��0I�[��8�N�k�;���x��������=�u�zy���b�T��e{龦�H�Ŋ�(�ּ�Ϗpշ'K"<�l�}K��zJ����O/Xi�hΪ���K�ҹ|dF������h�҈�s��ҬIwNVWh�A���#%G��2�z!�6��Q^_f��/�^���0yZ�2 �rx ��p�=%���e�6������і�'$�Q�|���fhXvh����Kl�,���F�;�C�X�g�0��n���bqt[!'�O˱�a�@]$��;鑋�!������O7I���XmHr��y:YL
e9�\�D���ɬ�*@)�������O��\�4����sf�;Q�:7�N�c����	N'�خ	�L�2;�3XX�P��F�g��='�+40/���|Z}\�7��K��)��ȑE�j�-;�ᆾ����5�u�0@�t}w΄�:78��rmH�tA�0�o��������`����I��s�����v�kq����l�<���Z��Ɗ0O�el1��8����Pi��*|���_3��;�{Ѷ7���&H~_eT���1z"���e8v+��Cmu�m	1bS)�L+5�ZZ	]�t�.��KG'lw ��E44�������S\�v�R��-:�H��*j��&U��\ v{[����v7��[��F��%k�:_���2ޛ��i1@�:A@�JX�(�TR�� ҧ�G\�x����q����{L��s�P$K�ݳ���qȁ�aBpaGri�=e2��?x4槎eƩ\�euD�<h��K[�l�f��h�I��8��$��q|��TqĮw� ������xV����]��e*�ZR�v���fiX4�M�^^u{�4��*('X�7���@VQ`DZ	t�G<8�m���3Fry2qwc���'���e����M������Y9��>!��[���WX)yW[�E
i:I_�E���?�aK�,���x���<�wO�l�o]�pH%��es	��=T� �M�Q�6�k��a)��ӄ���;>�At��w:��C�-tG�6��n&A�
X� ���L0?#�uJ�F��C�����Y
��o�b�q�/s
�� ��]n�
��ˣ�׏c�d�0���Q�+�p\H�+�T�PՎ�� Ù��3cuv�jk6[f�0U�%;�5mG��A�t�?�����Bv�����z��	�%,(qC�GA���I�};,��q��)C�E�rm���դ?�DX<q*��^��,p�"�����Q����ju������É�O���4��U�YGb�<Rsn��^š�%=��
�Z�ܮ�sM4v��v��XB��"cy��H�d�aސ(΄��\���o'Ls�[^�2�6θdz-ʱk��K2i�v�nezsKW��>�}��Sd5cJ>Z6����6���+�nӗ4$��߿<��j��!��%���W�����HM=).m��a����2�ھ	d��������S�V�I+I�U��r�y�*���,��Ԉ7[_���_u0�H/F�9��JO"��a����dq9xN�j�=����:OE�E��/�Den�?)�sL!Z}YR�,�D@K\��񧆫Kĕ<:��*;�Z�5�V7�1�!�.ȅ(�����3�J:�E�/������Pu�&�z�	*r�?ea�q{�M	d��Da�����'D����`K��,��mqH���ym/�F#���}WQ
^�O����-LŲ�a�i(�ɩs����-��M�"�#�L��JF6�\��J�S{�%��*�}�`QJ���1�� �SIb'�h����Ex�ZƐ��P#El^R|a��g�W����(>�`ϧ�S�>]9��wUd��MЛ��m���O����@��\ĵ��
~ϙ�`r�K�5Ĉ�Ls2+MH��\D����8w�f�Ui[��F��; ��V�K]na���z�pͥJ_�`�xX���N
.��hq��^��C�?����m�2��e�Z��d��=���f��;��_�ed�H�MR#^��C��LS�Zm�Ё�\*��T?ُ~�z��Z��Y�j4;ޱ�������4��V%�������z�6�|�0եde|�+D��㟱���F��%����^	b�M6A�TW���HY}�p��!X�C�E��v�p$����5՚�K��si>̘�L �~7X"�GA����Z}Ӯxg�}�*��8m�ss�oV2�8�t��f�e
{��
��*C�,(
�K�eP�����K�K�8ַi��E�}�?���fE�������D���n8�l\Z����!q���Ԓ�~�+��j�*���Z�p�Y�"���p��"���r����@��֐2��2@\"ߍTVyV�+F����
P���xUq��(kƎ��5ǐ;�QJ�ǈ���9Zv?@2���y�I��D�]��G��b��C�@a����1N���y9��%���f���b���1��6�~W�>Z<%�ͿZ�nOm�7���h�����a';2�s��'��e���-O(J�eZ�(�hN�Z�p��V�|�*�՗��"Kc�1�m�Meb�\�Z��N(���ݬ�;�Ro�8��C�g���H�lQ�ì+�oNRB�y�����:���2z}&7`��jiM���z�$�@OǀT�9�N=����''��J�"e��'^2.%"4_O�����B��H�Y�F�{�c#���k�{�/����a�|Tq�j��nW�d�'�����'��|�T<p���Z�bo=�m�~�~^%.T�fKR�����f.@'�n��!
O2��*��N]�-\�.�Hޕ=&;�ĠiR�3l.����{.+����Zq�:��}�(�"���FEӒ
[o� %�:�$V׫Z ��(�8�'�y�D�?�]ׁ�٦�s��g�jTx|��b�2c��[�b3`e�~�{�����_�B�cB�3/��S��wE�%~���\�P�[xT�/Jp�%ϑ-?-BHe���m�#���]��w�߬_�Y��¤���q��&�-�Z�tw1`��� 	-4��_�-]�tx�7A�� �5�em��$c�`�RQ[Y �s�LV�o����ߡR�V�o�ǲԡ��X��Mn��{��k��`w@�Y@�h�_-�5�_Ͱ��Ӗ7qtxx��d/�CB�gI᭠���"gyR{X�x���а������Mx�<z�!�Ǧמ
����H����-|ȳ�d��c�g7x�9~�v4�]vP�a�p +9�+����F�ڰ߭��)�|�-��kk���1F~�i��y�������'��|i��Q$aNRQ^
��h�{F �:W�EH�#v�����l�V@jT����|�(�4���۴�D+���2�G�/F�޿:Ѡ5�Y���ހc>C/KR�̈́��#��-��~I؝��Zw�"�A�m���ܾ��_)��0�!���L}G(�6OC'�]��}��p�et���J���.��G�vW w<{�{���`22�e3�7�w'�-#;�[��"e��kC�%��2�A_������*+��̀%ٰ�Fޕ�_D}c.���#*ȒA�uw��1�c��\럀H[���3C�w%����Bo��j��&��N!��������E	�6?�j�'��w<�O��d�c&m�KT6:Uy��u�4{�8���g4��[�iu��LH�����0�S՚�1��h��1p�t������C�ci��ywY�9�.�=2J�D.��ðQE�����V�e�qs�������(����rGI&��q��ZE��(n>���և�P[D&�oOF{�Ø��lJ�G�s!ߵ<q�Ŗv(��iZ
?J���'0��VL0��X�&;�Xu>Ծ��ʿ	��O���3i�7b���_�I=�)�/x��9z�uϨ;&D���}lE��減DGxp$�%�/�!���,�I��x!� ���|~�	��1Cz������� :�z�?�5�޾�Nk�Lt��!�
dir�"j��X�p��~׈���[���.��)��N��ӎ�͡��K?����{�JT����\	!�,�!B�WӓI�K�c�y�"I�S�ű������՜�$_��z#�@�^�A-�*�Y�� :�W����[��'̏���v�<%�av�r��_���Ш�H�@� �>n��3eNa5`���R���;��?���i߉`5e ��_61����ti"L*�C�ٰOr��{�B�%���ze$)�P+��XJ�̲z�3��O�F�}��U�6.�6fVѓ�#f�?N�X����_�����4�Ȏ��5�,N8�;�I���ZBKDFI�e�pp��E�s&mn�P�Z�9���D�)���*�V�&s�šgO�G�l�?�r� �ϕ���s�m�k��/�C��RO��~7�~�����K�ԯ֋8�K̆�}�%�1�	��E(���Y=9�����>��>�/|�gh�CP�;�y��!ɏl-�w��է��`3Ǌߌ�"�8����֓�	ہD�Y�\�'�z`�N�t;O%���QӬRDg�%���s��8�R���g��K���V�xV�&�l�˹�V@���t�gB�'��|�2���<
l�@��~1�[��\o-P⺓s�hC�Fyֻ����<9z�q��Â���(�M!wq֎5���ӓrM�l�s�Q��%�MBqΓj��5
0JWz��H���.=7�I�ރjNY+��F���@��,#o��n2PGU%<p��K��돻��$�E�Kl���!�A�#��_+u��= [��	���)g�o��q=<���*.��ɍ���d��b?��ת�$�Wx���K��ƒo���8�g'T��n1�R�Zc�Y9}�>Uc�P���#��1�SG��G���`vb�߽_1��on�_%�ZUي_��_l F�%2��x�ΩI���0kxvu4y�����V1��Gc��#�z���wJ��ѥ5'�@ɞ�#l�^[��;���:W��L�-n��+�)(o݃�O���B��v�юp�8�6c]F|�)�"��Dk�m����>��7ؾf��y�_����ڼ�ƩX���J`5"_��I��ZK���Qr�Ro�ɝV��tX���G+à��f2t��Jd�� ������{1��u{��{2vz8�yt�h>�&[C�vM�
������xs�\���$�xPMʿ �p.��:�FV-55J&��PV촢5t�$��(�^r�8���}kj�>����0f�4p+�z�����x���T��x��Ȓ�yL�����L�\�[�5ԝ 7?\�}?��|���l����K-�Tʂ(��I�0(�oO��V�K�&E����~�n1��� ��B�W��}�7�N-���ޟ��\�ҺƋ��L��d���G�a:�F��Rg���}��ǆ�J|���U6�SǇ?'\�0ժ#�+�@�.\U@�dc�Rfv]��(V�<F�)l��r�q�eG��f�f ���E���J+=T����úg�T��`jN������ؔzXT�:S: G�$�}��^'�t�-���t�d�'t��łNDWx��1���N�
#`��ԗ�ڼgsȡ�61�`��i)
�Eĥ���ur��@Z�uo\xt�@ڑ��`�:�q��@�'J)���8����0
B�W��6���? �o�Z�����O����}~�>����i�dO��X4�1���"�{��-:<P�8?�v����Z�R��R��՗V��.
x����xfH��jK�\�yj���;	�M��b�� ��x�6Ԇ-�R��O@KF�+����&	g��M��^�x7���5G����"��ڻsа�T�%ц�c/��X�s�Y�te;~�ؼ�7�{��Ӑ�� ɹ���@Up�����|U��[�;|~�aY.�����n�0KB`��.�ȋ��:�[Ȇ/���Q�դ<�g�!���a��S���} �;��.�)��1�i��E�R[r��G��*�d��A�HtgA�Q=�	L����W�e~e}�?b~(����lw]�*-��F7��Y��#WQ�ϒ�j�h����(^6��B�j�]��f�6r����&1k&��օ���1�+.���kY�<]�'$�dh\����WAF���4~����E���_� ���Ԛ�;�D���I�Jϑ2[���>l�O���'���J�U���=���պ�plp��΋�zӢ.��Y~^��Yr̒\���}�f���=Ȳh `�r>E>��8)og9 ��T7},%��
>�����ȝxi��q�j�g&�����L����R��a�^UC�7(�o��s�H�`�;Z,�!N@jVW��z#�����P�>Xn�M���M�$���vNU�#7�~��Wv����*~K�I���Nz����;��]璎lh+����|����<���'_�X��>/�g��RA��۳~?	�����q)1@�`���.	��E���A?��B��,5Fbx1��o�~G�{<To�����:ح�w�)#��0>��$34*�!vuJ)��,���b�Tehܰ�t�&ϻc�Ӗ!�2xq骟�jA,�xFsrqQɪ[���Kl�1�Q���>w�1	cx;�Pȕ�q"�
w���o�5�)�����:<�+����st +�ʪ�e�b�;*�M�M ԣ���xz�8��~�?��L=��7%��|�����S�G��p�]h43��q���6B��h?�5����S�l 7ɩ�I��<��ȍ��*
���q�f��"��kF�W'�����g$�xI��K��N�o@'|�ĵ��X�m�S���!Ąke|ձ
�.�̾���#��MǇ��7oA��n���)b}]Fw�#'%N~e��(P��+�A��Е�����ri=\�x���ѽ(�0��nP,���idM��x�c�Nrg<�nV�ZM�Q��K(	��u�S�:v�o��]����~q��G�2�b�yւ-v�*7����ͮ�
����h�2��1,���Tz�q}^?�l� z�7n��F+u�FV��t�p�?�� ��n�"��j���"��,�b�ֈҬ]N]�OL�Kz	e;t�%��f��4(��7_�=��x8���K����6y2���L���؞n��"sS�}�����`
ɛS�uI>8�vjTn���2"Y�	��eBh�d�㶸���qH�#�ak�v�U��e�ך�H�㫁1�4��4�v���¥	c���L���1}����jД��HS&!��5��p�s)J�S�F�z�y'�S�;zD�m�#]es��D��f����I] �ϳ}x0	�����[�v 3�ڠ��`Ϫ_x�t��R�\\��)7�Ё��Q���n�ļ-��W�˭~q�NЖ���Z:( �JJ�Q`�h��ى+6��L�=��*�0��+����ZOx�	�Dg�*��@s{7O����%�.-lT�8�$�B<p��/�+bm"�1�t��\���b� p�ԇj�am$l'�;����S�;^�KYي�;:mpJ���sV_}�Ͽ� �� ҽ�A�9���$�f�*��CC��N��v�	����E����:�%�������2�@@��h^��e�YWoCX��I�0��pDC�nV�C?�X�_�����S���xݣ�Ļ�d�CSGz���,FP5Rk�2����U�>�f;Z�S���qI赦�"C7���9��̮���s|�ckNɇ���k�i�l�('C��~�;�����5�����!a�Q��+bl�d�{} ��t���VH��AwȇfQ�"����w���*�m� D�Dmv+��"���.B:�
I�R�M��Q����(���e�I<��?\�� $����D*g�b�}Yi�9����g�늿A��C�*���r��x�3;�q�H�3�Kb8��,TeܬPg]�`��r�u���u(PQl* ��C��.!0��ϋ��v��45���ep�O��6U>�`�[\��C#D��FW��FXu���u&��ׇ�A(>�Zh�j֠�YD�%F�w��t��$�+=�&�p7�>W��Y��Ҋ����(p�o�K�,���W�z�@;�J���z�Q4%���+y/�-���֬e��tě]ݞ�n[jf�?�ꪚ���qǍ�۾�ܗ(0iMԂ�
��h?(^��"�OM�~T��i2S,CT~!5��;��d _�H�&j�3�b���<����q�8�,M�v�d�k$�y'N4@b����_�݆Z����4����9+^F�@���]����^��^��I���!��<a�]��t�0��IzB�C��$A�����/���7z�P+�hfs_p�9pD�N��~#�Ռ~S�s��&9'�q�Ym���1�=�K��,���Pu�AM1���7��
�+᳨
GQ`�n�b��cT����F1��E\�V�<߯\'{qs��Q�73���(a�C&�c�Һ��J뤹\q��8�v��[U�{X�=vLXN��u�H�Y���=�N:9�9A
�����2Dz|���c^��h�}S�Y����f�o����kYX�<�Mpq�Y"Rc=�i����d)�z[=#��*v��u���#f=9T��u��~�~��ym�^B|қeL����K+"���&�
 ��6�V�gw��Q&�Aaq�%OZx�qУ ~�ZIf���c�'{Ҝ���tG��4d����eO��c��d�2��ӝ��! ��('�}�a�F�4��#p��-J ��ԑ�J4z��0�3CӕL�
r��&U��Z��<z{��^�=e�%��ZO��'Z��yJ۪͝�|tf�-�w���Q�b!;��i���]��@^�c�r,C��N��j���*���8�P�gR�Ew�_��&l�(�dTUb���Sp���)�Ⱥ�Mm佦=�;�0�j�\�1NT�w)�m�_lg�r��Z�����g� E���6)⟣��7B�Yt�m��	[�PP�p�hk�k}�:��DE�ao�����O'=�	л��e�@P]/�aL�{�F�^���TZ �S�a�Uޖ�-Wj�d����/����c�D��z(�;��xh��!�� )>���:�s��t�&���ɪ^��� p<`�� ����G�7�z��%���./υ����"w~K�����~�;�9	�+�U�wAd(oA����k�����>�[9dEN!����y`<�}�������G�x������p-¼��N�x��xWUe3�"������Ō�>��M�7^�(����ބ�j͎,Պ���h_���m5Zsй)H�}1\��X4#���i�/7�y�����~h�9��wď�G�7���x�v����rƍ.h�vD�H� 9B��zͪ3ފ%���+jH	���1;���ɻ��ޭ�|#Dܜ���������u%�K̏��k3Xt���\H${� ��W��k��#G,��`-�7N�����Ct����2�B��0�yC�#����.�A3��(��^s��N�B��:6�89�L�ƒ�YYk'gsт|�%�Ua}��0��/p�Ӑ�D>7�-L���O�TE ��d�l5��8%�jꍐ	u�3Y���b&:����o�����M�_�z�}�^����޽9H�ه%�H<XS¼�ն��E
�:����Bbs/��`�!�2^I�/��=�Pe�.��"E'�|���Y T�qPya��?Y�/_��+��O���+�s��k�4����aR}tb�E��W��G�Ke�r�B����7�k�L��]��m����	�8Bd���`7�4|^�1�DS�N��k�pO8�Q{��n�L���k�K0�s�ύ�/��� $m�գ	��ꮎF�Y��'mY{e#��H��Ò�a3�wL�U�U�����X��^���\��7˘�&C�&D��p^{n��u�]���a���t�9i+�X�w�q��陶����" �\�
�����t5Rh{��F��	
���<P ��e��]�~����4V�aR��H-`GL5�$�$��uT����#q�!�H��f�=��Ί��������?8���n����A9~ZM�-o�
A�����亶!tW��2w�a�0\\�0&\x�oS���Y��/�"���L�EK{ϳ���K���ϯw�)/QtSoQP��O���B*�r2���}�$YgU���g�!~�+�n��n�_	��Y�c c�A_��L8�;ZN��q¼���i雎��6e�'e")����+\`hT-&D�$��!�f���O���R�GOd噗�6�������Zjb2����=�>�UZ� w��]Ԫ,��D����w�Qg��hv���:0��6�v�|���
��-%f1�&��,8��}��l�B�[O��,,�g�ڮJ�$�"�����/��_��i�ð��÷�Q����#"z�+C�̓���8l��tX���G��i%��2K$&�]�Q}]�?�����Y��k�7��^���h&gt�h.Ġl�_�G�p�����..�c׊��_[@4⮖|}5x��oגf��n�Λ�Y 6�mk^rm2�|}����B���"+�ǒ�AM��$t�
j�Õ�yF� ��&���&JR�`�as1�~p�n��ϓ�j�qɀ�d����D_'e"jJ���n���.?n�KuRl�G����:�E�ʃ�=����j9���d4#S�m?���}؍���1��)I�Ŀ�bjK�����(g��\��h
�Wb��<4W_)�m$�ׄ;V��?�d�ViZ9#~j7��q>��v���]�Rf�S&^��;\\�sA��\�Y���Z�)���>�r���x�
RsD�y!S�صL*�k��9޾����ZP�aD���lf���{ר��U�L��>�b�v�A7��'|���Ᏼ�܈٤����� w��v���;�ˎ)�և_�x�} g��iɊ���(�I?�����&5@�90���B�gY��-��0h��(8�E�W���Y��~7'j�:!eύ�wM��,�V���n���?I�(���BtJȌ'�r"�l����J��d�t3��;7�ͥ"�Ĺ��=L;�kCg�(T$�>��*r�E_-4~$j�C�@i�k�@�jY�b��~�R?z�)�XH�~7!׮)��TvY�r}���$f`N�&2������=�rn��7J͉^<k��!
�+�C1��ZA9�tI���f����C�s�t��d�Sv�v�rz2ae�̵pW�-���7��#'����+��m�~����0�M��wd�[J��+z���&c�=�f1y���зZ�j�d]/N���=����eA7�v�
�+��]"�36⻤�QX`]�l;Rcv�j�e�V���X	�?{��?��ܢ��N�k�jCu�6]�0�zy�yPX�Ӫ�E�Д��K͡���(���h_ley���U)6�$�.��[�l���6���n|�h��>�ŉ��F� *�5/�C�*�3���Y�����Kݙ���&��_��T\�9��ތ3+sͬ�ěm�����r�>��H0?6ůhffp��Qm��
���'곖�&���%�o�~:N~�3CO�U��a�Jn�v���N� ��4ZR�k��&�*���,�+�j�iM�̍Ƥ���c����gGDc}Zi�9�1� �h� �:�@�k<�j5?e����>�v�P��[<���HN���Hn۫����e.���NL��2o9� '8�]�*�h����<���uS�{��Yz~���{[��3,��G�������H�W�ID��ϻk�F�3Q`x}�7�-��t3���*(O$�(=�k;���}E��KM���;��A��R������k��S��B�Pj��וxqo��q��)�CKw���ا1��ڨ8T�U�W�q�P;�N��3����Pm�c�g��Էٸg�7�����ʈ��:�Օkݨ��`�f�9�I�{���gN��Ds�%�Wݬ"�4۔���I�ed��I�~@'#Q���~�n��1�x31p?�Q|rR����k���)a�A�@L�YQ�9�X�z��`1.�B�q�sD
��T�ao�O`1�r��*0����'�i�_4�B:�F���;��7�O�����k��u�O��X=;��	*/3�c��J�ͅ�5x�ԗn?q��
��zr�+�>\�hq]u�~�멂�]D*&��/K\8�E�d�k���!�H�������8�~�#/��aF�sh�o�}�L�M�^y�Q�$^j�������-�s�|O!@��黎��i�8,�1IK{�>�Q���q�*����C��h�/IV&��؇��{��Q�z^�Ʈ�@CbVǶ!��˫��l��,|�X�Ş��v��U���6��^.!O{����s�;�dpY;gj���_߬�XrS����/�w�R�Km*d�s>�T�b��)��R+��,�K����J��Kw�{��)#�i ��@����>5y#��'�?��r	���R��h��3��P�� KR]�����6�Wh���9�\�^���{��D��-v&Y�``-��ۧ���V@/�����Bh�S��Y�":�-¶�!p��	)Zj$K���+�k�C�?4�,ϲw�v������ֆqې�C��<�JGr���=T��]��v��+��h�׎����7T��w�B�b1�k�����	���o�W!��<j���Υ�藃L��ֳd(>�Q����׷2ʁY�M��t�
�F�YWޚ	p�t�3I��^��G�*�q�C��A�y�=]�^"�����j>��|���3�lVLျ�������*���s�t	�ǂY@�D$�������eÃ�V����ZJ`A�#?0����H$x��G�q�+��L%T9-|�C��$���NH�������mY�ti���7N\�YI�ӓu�����3	_���n�j`����5�}a���&
g��%�	0�#�&��i]��<�B��nY?���m�g_�]��Q�v[���YYw]Z�����03��h�0~�җ������1|��s*�,cl8�i �D��qk�m>N>I�Mc7�G� 	-���P4w�M7�h^�
i)��J� GS��	��G���cK�)y�+3�\c|��ftp�P TtG�j��@y�V�����A�� ���dSf0�A�SS˳ʌ��m�Q�G���1�*~F=�����9�k^�ʀ�#nUcS�IS$�x��B$6l��O���ea�ڇF&��0��0>�A'n�wi�?&�⣹�ɪ�i�5�C�1���3ۤb���U��
��3�1�˪�.�j?����۰�� :�k"�4
�s����j��Ǖ��L\R����5�I��R��)A2�y�)�|�6���RVJw�uE�"@�8�O} �Yqd�2�Y���޿&d'ax����'�|���s���$s�I#
�#�m�oؘJ���`d�z�zHut�?������i5�b_O�UsC6vcE�롻�K]�"cX�ae�k�k��^�jD��M٦y˫5�F���F�E����l)�m0��r����mwdF��v;���7>�+'f��^�m����b�����M� ����]
AR5"�z�W:�\��e� j��o���I�
R?qo��/������]�<����a�gҎ˟���q�+"�5o��)�o;�tKj�G1m@��iA��=K���N����+x<�(�^�oI�0;�����5��r6r�Y�t���i}�*��k��tUv�S6��q{4���]*b�*��F c��qV�(Cm9 ����P*��	B��M��+1������z�ޫF�EM�Ґ !%D��*�R�8~h&�d%e��`2掜kP�������)�$������A*�%YXI��)v�䳳�� :;�+�d�1�$��G��̱<6��[��L!��ͬ���Ǒ7���Q�_n�^��jy(F%BG0�c�����H�n@ �;��zv�.��DkO��`�g!�9qT�����v��{Sb�9��@��O�����[�Z�6�a���
d��{��<ߞu	anT���j�����/؆���o�Š�8ہ+R�*�G�O��>C9�h4�����<�,e|G�
����'`Y_�nMf��ux��l�"�1�mR�(�Z�'D���-�US��|����unH�"H�v���W���VYgQl4p}ٱs�/b���m_Hш���K���F$�|P��̳�ɦR�����)Ca�i{b�/ia��$���B���LFa���C��Y���#�8�X�@p[ ��\�+Y^B�B��U��w:�ِ:�rm�@�~>-�3���?�fs����.��ӴP��&�o<D3�cE�0�7�+�hǌ����Z�hGZO�CD�Y� ����&���I����xS��}�M5��WS�>�AX�BŞ%�:��� �`�㶰��V$�5�?�B�bZ�"�T@�*���+��O�O�8��i{� r���5fy�u��D��#�������-��==g�A�����ֻq���S����Q`ic��3�M�?����A���f�.K	�c����7O�+���_ �끚ʺn#/�b�oMY0�c޺���[&+h�D_������m$>�r�W��~?s� ���cz2LUL�"X9��cX$�?.����}¤���B/ڐ�Ú�'S�g���6-��|#+5�Џ-G�-zư@pf(�<erdL��V�(�蕅�϶ę��)e�̪��G<���!]I���+������� 5q��3���K�[JR�tN�@/�O�m��w���kdǺ0�DX�>�ש^�� peLX�V���D3�E*�ZX�ǫ<?4>��EVX�fq]ʢ ((>k��Jj���A9�|����Ѭ� a�0T<�7tF��Z��%��h-�����n\����~�`����_*�%��^�t8d��<�	��
�:ߪآ)�OL�?
=�A��|�(*����]���fk�Q������;������W/�Nz7���^���|-��s�XŮ
G�4V�$�S-�t%Nz<+J�sr嫒���R��]�l���f&�9X�&~��ȳ�8㷒�c�"� M�}pA�f%Ѱ䯜������t���^B>�ȷ������<�.&�F��6w����;uD��ʂ�up�x��K��Yhik�������4`;����t_�Be�U�A�s����E��C�oʣ�*�ty�z��Z��,����_#�	6;�Y,��u��y���R20�+ږ���n��"{�;(=��v��7I(XOzp��\�������oY��S�r(OW�l�G�$����[�藞�&�q7D&3�=�_ ��@�w.�(�� Hn �^���)�8�$�Q�eپ�.���{*A��A���T�Z<K�H~�r/�{��p�Fc;d1�V�\�]d #�F�	��3��,�o�L7Z������hs>�7bS�=���xH\d,_�c��j��	�9�J�KJF�������,D��Z}?dK] :���s܌�j,C�!֏����Q���ڙ�K��"Rv��!����վU�h�}d�sx�PY��۠�m��B)!/G�5���w�@�&�{�
��­_b}?�N�@�]�?P�w��[W��>TΖ7mWڃ�5hŒM��R5\�ӈ�I�4�uYϴ�[ie���^���������_�������s�4�,*��\LB�!�)�b����@�G�w�ͤ�]Y �L�����EX"~�S0�!An�j�w����gT��X���:����klxX�)+|)!�R�ZMa��W�s2<Y�?�w8�����9��6��_�w(l@2������If�<�;�(�c��s��x��|�Nk�1j>,��m	��4�>!�������峲����!6��C��?��r�;'q}x����r���h��p�o{�:�I�@��:Q5c�~������~���Q���p5¸>��n�4�J�QD��ǑH��nZj�e��b���^��e�R\�z;�j���s.0���ۃX/��[����L4��a�{�(�.l�b�TC^����P�Q�>��%����#�ܟ���;�P�	MT�z��-kTt�Q]Z�Wᷣ(Ⱌ� }��M�����+�s�K��_w�lo��E����jp�A{ɖZy�"Λ,�|�_���g�Ȯ�d���4�H��{I���ʨw���U��g!�I"��ޮ�W�f�-�r���Lٯ���IV��&��q�R���e��l�O+�ɋ%�b4���isB�O�ݺ����s�.v��+�V��N�:*��(�����"R_�'����406BQҎ: ���
a�Oױ޼���i�>�[5n�jG��}���x�#>~�s����⟟��Q�U	���p�m�Rd���@3~$'��Vv-f��J�%v�������z����/:',�?PĻg3�_�[HQ,Lp��?���z͖�_�Z�;�c�5F�I9�QW]�q�D����.�F�=4����
��DS�gq��C�ѓx�c��h�=N��U�!�)�XN��`�L�c�������F`쿊�@'�ٍ�^�'f�B�v��Ӯtu�о�0Ŕ2����<��a���/|<q������-�o.3��D�s�h�_nB�o/��bUojU~��Z�+whb�$;Z�� l�0�!���R}C��������S]�q>�p� ֽ�Zk<<��}��b����m�uZ���i��ޢ����6�_��;��1N�`��L;�2.����j��nҐ{OЂ}�n�u;��6V��J/�&��KR�Υ������q#�Rv�ƩO�`�+#��g�6줩[�����30kŬ����V������?�v�j 3�R��<}���+�};�M���!�v��"/����߭Ժq��+���*��sոխW�NY5������jn�^;��o�\��E/qH�f�%`µ�i���qP.��w+��(݀d/3��v���2�Z�#���(�D�2�f(�h�[�j�=(I��W\Ȗ������w�YsM�{��1/�!&V^�{R��w�a�<hP����B��@4=��gj��~�9Q�z�C`�ҮyM��
���P��;���c�DΆ�H�@��Ъ��vHQ�z7ЯtBԓ�oFZEd��8�Vyup�K2�%a��]K[����q�����3�t*�Ic,�+��X1�vg�}G՚x&N��t���5�3IWʿ�a������6 �))vP+
Ŝf���8�g���HpB<�u0H��� 	����s��e�8s�!_�(���\GUx������Ӕ�9r�������S\��
��!q�C�l�5*q�U	����ʾQyn0�{�T��<��!a�_e�VZtP�e$D��kI	���b������֦���p���H�ɏ5�I]-�ק��7����gh��*FnJUq6��~	��-�.?��bC���io �$"��I
�@��Xs�@���	�I}BRo9_�����V|�Е5�F
�,a��4_�ޣ}���<��-G�yO)��<<�#!k��.��11m짲"3��N�{����[�b��B;�E48���Ţ�\�(^$i_lE�Z��QhM��֑���E��V��`ϥ���R�eN�(��%��$8j�Az|�h�Ho/�qn�����r��(/��o��,Dy&��Ĵ��JN��J��+��z�#��ݫXq8�� f�̖A���r�=�1dAx��%�S��a����͐zJ������Kk���_�b�STAMq�9��Q^D_/����k���2�'�.������]�N]*��j�#�v>��2j-����g�s����}0��8>ޛ�n��3גo�q���]����H�k��&ޜ�w�qF���G��ul�k%^�x.�zZ��]6�� ƈ'T7�B�&�{S9����-:��%o΂+������R�����|PHq��
������,��Ԏ����_����?L�dd�l�r���u�t(05��̲U�}K�@������^��0����ܓ�����7+�l�K�J½�Z�}��מ�$��@�.g�J�F [֛�����`죀Ǚk�􍄊m�OjȌ	��I�G�����-/�O=�?��GWmf�)+y�7����޿o�ILD��ٓ����L&��U����T@%�%^KУq�=Zt�Aj!W��q۔�'3��~\�L�1�-��s��ڪ�H�m@#CJtLkS����q�6D������>�	ק�p�(�ͤ[���I}~r������g����h?@|�	R=�U��c�ԅ/K�9P����ZR���w.&��j���(��@pMKV�i2�R�}1��g���&<I|{�moo�2c`@��k�r�ہJ�	�A� �\���w�O����_����K�L]S�t4�S\�[� wݰ[�o6�^k?ɑr�r�S��O�+��L��O_1�o��V,ޫo�hGj�������&RA�W�}��-v�M�F�Ŏ�N��同���f�x�V����ON�G�a�O��U?v�0�����M怺��#��Y�x�Yc���Na�qF������{��J{a��|��0�����H�P:�
fZ,�Ps��-��Q���&~}�ߘv�/��'���D-�u�r�ƨت��z��	��<�y~"'�j��n>�Գ�q��=��!>`�Ż�I�Xxh�ui=J �&�Jb+�D���]-P�(���d#P߃nX��E
��bt�8�:5�����m?���붛.���z��Acg4#�ۡ��y�'��ڰl�]N��%��3JV��^�i���j_8�D�װT!���A{��XĘ����~�[�_eN��a���	�~��,���THnɗ���)���L�Ѿ��ܱ�u�Ǘ�]�i%Ruד�t.�,���&U��Y���e���7m�y(9C�C��Ik�+XW7��yR/T���jئ����b�2@��_�yX�vN��7����p����p��iG0ʙ@P ��WXM�i���#y���+�e �|'������%�?*B��ǡk�G5!��]���¯+-��d��o�YJ��9�!�q�:q��1eP��-r�n��}&@���^�2X_0pI�גB��MxoB2����h��f|�%��٬��`��B�@T�֩�����G��Kr.�����l�x�]����>@��i�&Pl����1P �e��t�gy*l��I�R���Zٗ�i��"��Ő:��)m:�g�Ԫzv�|l�����\h9�G9���7����� C���S� c`c҉{��r`���f���ʮRyR�2��.[,|nNW���x� Q�|�Qʹ��A"���.r����E�R5}�ƃ�.�ә_���&SF�P�U)�2#2�%�h.�o�A�d���&lmr�,�����=�v]|�+��Ef��;��r�-q�I��y���^"������{��E�t���I�T��A��w��&T��tyyh��p����CH+���������8޴�6�ԏ���*CMU}%���Aיx���G���n^V��b����\̒	"��c���p���T�؃�q�#U�P RN5�-��Sk#�P��7ٴ��?�80�4���4Aא ����/�\�����cZ��J�@<�79�� :ʠ�k��IL>U��Q@�5�'�,�= N�W#��3��I*���I�us ��͝��V�P��Z��젭�j`XR�ag��#��%�N�a�e��� ���+�Er�T�͂$s��<}���!C�Z����˯ ��ۆ�F��M��]�	�q��ťy^o��(�O��P=5_���	�`�Cp}���6����o�ܻ��ǈ��O��V���/�u�xxO�WS���oX_9��q�٩UJ��߃�u��_��{+rt Vk�K=�����T#���N�������86�,�씸�A�ai�3�v��K�C+��%������/���3ܤM�����Mש�R�kZ A��E����n�*"rSC���C��򥄦h�*�j�:���j��D_00E�r�A��]����9���@����������WC�AHn�Բ���P�bV����T��a���]&C���5��Cf[� �&`��1FX�Fk��v��:O�#�`Ϧ6�Xi����穬;��ޯ��`G
�Ɵ^VN��Ra��#�OH�MګQ��t�M�7�sL�0de��ܸP�ʔr���>T�.���d��u�h�����+y���Ȗ?��&��x��|�9�ٲ�����8r]n�f�g��3~��2���'��M�	h��s��|�NI�&Z
��!�Gp���y_�=�?`�]���2����ԩ^�O�2�KNK��·����Ll>�z�>�+��-Xy�k��ςKA~A:]h�u�.�u�V�-�K�,�W �@<ˤ�Mκx�ڝ.B��GB�!�M���;�#�d�XY�{G�@Pq����N��ArA��ٶ�F��7j��|��P��T�����8��&s��� ;��>ZО�ߌǱ��ӧ�L鴭=��H3����OK��IB�����Y]AW�Wح���_�Z�����ެ38�}�kz�l|�/���h�����U�s���xJ��n�OE4Ux!eYt�I\�~UD1��B�.��`��9��-dR��ҵ@�����%�p�l �r���W����)�qT�̩�#ѝ�:�c
�x��i`��zl]k1�ca6�"�~L����o�A�+jY"0���+0�{`����<�->Z�k�/�Tq��$�$Mف�8��@/���E�%��A#�]d2�Q�#�Q�Ƿ5P3�˰�'EF����?�b�mB�;	�=c� zKh��s����/���M�"h����j��3��A��G�}IBР��Is��_��)�CG�J�g�����}Կ�+�O\mLsx@��a�>j/Y	1���]�z1�(Zq�?M�pFxp��yW(Tr�Ǝ�?�B�ڸ��ј�|5	���CL�ߟ��)�ɞ]�u��"��X����s!�� ORM&A�؟X���H���#�:��������cvM1�ƉU_�,TG�K�iD�+�b�h�e�ֵ���ݚZ3~�l�������7qe���a�N˲z��t���;�u[��:�FQޯ��E$��N���p��p�k�1���迵B���[�?o/ّ�66;sȲ4:��!s9~݈D����w}��<x�6��`�ڒt·�i�VR�\^�"ϰc߁�e�����_)�G����줚�ȉ̂�A���$3/
8T���i���{璔����?k�[&������ba��|{[@��/����9]���`��9��� P��(�N1���#,�#(w<~g�5+�,�Y�]�Kΰ�oDd��Ig������>,�l8�����s������M<��K��=-SQw�/���͹��r�zU���Z�J�5[ft�x6a���x�Hɯ(x�0|_���0<��:�6�=$�x��r)V��B�K|^�`|��L|'d�P7���P�N����\��VQ����n��.�6$/���,hlji.�JiQt�Ǒ(u���kh���)�H��!�-��X@�hn��n�s��v8l��@_(��3�^�G��OY�t��M����A�SJ�]������.=n_���v���+��(�#�o�� <il�G= tԫ�Z���Xt\���v�@~S�Z|�X_h�������C���ҭw�P��9+�����D����(M��KtP��g=�����$0�+zt���@ζ���M�waG7�l���*�my�=�|��з�fjđl��HŁ|�љ���� �C
�W!�|�k���:C����kM�C*���b
LJ�?��J��j*G쏥r�'��1%W[�t��XD6$"*��b:��z2��\1
�9���<�ra-1�qcoɭ���<��]���$r�9S��&�ۭw˙A�.;��6�,�k� �ޖߺ�4�|���|t{�L2��������SZ�%C�C8+>��܋Fl��EO>H+����|�u#SS<G�V�gN[�9`_`*�~J^��M�]ܬ���R��?�iD�d��m�@ŏ}��Gf,_��U�&~�(�B$]iS���oq�����c��Ts܂������]㺽0F��&K�wf�s'�˪[pm��h��5c�W��l'��P뒲o��YY�Z��;V��׺�Ё�~�G��[]|�73�B�:dͷ��e|������{�lA�k˂P�B�A	Ů�w�l�*6o^��D�SxD�",���LkI��߉6�l�`����o���
gx/��>�Q?�=����m�z�iw��pQ!�H�K�hP�y��̢�M���K
��:w�x)&���_�q����Y{m�TU5�|��:��O��@��׋����'�a{���b"�*ݖ���zB��3���n����M8s[��U�����æ&s�6r���R�u���(���'X��ZX���'2s\>;�ܬS語�T9���˕f�s�VOɶb����yoe��4�G�ѫ��n�m��$[�����h`�w�X���g6#���4���/n~t%i���N�Z�����~�QQam��*�2��T_=���̗�jBv�� ���S�����`�m�N?��aG��	fõ�����F�TvfTP��8�U(��CI���qF�p-
���nBQ�+�FT0��������,���\�V��ݶ����T�&\�H�2����W�#��p(���pG�[M�N�Hŵ�6��7�	�N������c{��	��e��P ۑ[�#������yv�WB��W�_����inXd�C�7��x���ʗՅ1ső��G
_���H�ٝ�:�	^yʮZbp�t#�3���:	wm�ݒZ��zMp��O8X
<YQ�[�3:X���E�v,�ƪ����_��p<��o�X�%�sr~���p�PX�\a	�3� ?ݧ��>�;_Xu�(�%r��+�yJ�����I���m}�%�B�h���Y��9�%y�Y�6+.��dȬ��Ԋk�iR٪�'�4���s�Ԟf��.�<�����72�����ʼ���J��Y��8rf�=f���)t����ǌ65�
����F�X֎�!�*�}�ּ!�$�=�C)�vn^��nmKŠE�����t3W�z�j���i	�8��&XR�A"���C�C��ʈ�H�
���8�'�?��u9�������G(�O6�HK���W��E�Uy�e�Gn��;˿��-�#Mc�߇��!�p��T=F������g\,��
v=��~O�
SZ��XL�Փ�Cb3xX+Lo�qh��r	�&k#���n��KBN��8��%#�l���T�|\��|"�-cN�-���%�ʉM�o�ML0��1�����˦��_P_B(�N��"��đ���
����yx�y���춮̌?=�N�l��؁���3�}ϡ�z���7׬3Ԍ΁S8�fJ��p�/�����j
�n����q?���/�Y�-(�1��{
���c���Tݒw$�	,�W����ZI�y����Y�ClB*���uhS�ġ3Q&�L�� �/^�����-i�������\:�Q@��u)�Ǳ��ilQ���<c�p"̶"ȑX�Z�N������@��,Z����N�~��mK����b���kU%-NӴ��g�0Gt-<ڦ�s���/h�St�%��Q.T�<���In<�*�@��7�_�����_����羉�����"��M��$�#�(�W��\��3�[�nP�j���	t���F�O�өQ���[��N:��&��[0)����X��D~�]P���m�5��kCZȲp�/Y���bhD?�H��hJ�P��X;?��N���'�y�`���`�AN��^�f i��Z��4�����[$(؟FbiE6��g����)HI	�W��3i3�O�:P}�'k~|]��V�3�{��'L�T�>]1�"кfd����Gy
 2�m�>�h�}��u�T����0w��zC!(g�SEi�s�ܤ)����z�Q����d���>w��_P�T�QZt��ƳH�켆ْ����v�Tg\�����(n;�E�2b��^����%X�3�I�oT1X&QJ�9���^��q{����p�1�$����6��ʶ��;�F����e<+����:��I슪3[��2�k�N<ԩ,�;�q��yd�ƈ��1S�D�F���!8��4��.��g��Dؼ>]�$H4�<Įj�3HH�w`��.�����P*��� �_�#M��v�R�h|J��=KR�(��"H��(�z��Nt�\�}��q��5������E6/�M5"�rm���wā�T��ǟ��M�{����6r	۪!����2�e�E��XzpWN�!ZNl&X"�}]����V���O���7�ß�)ʜ����a��0���P�� ǢsNy�M�(����d�y��>��(�m,<q�׉]���i����#�ړU�]�"3�\H�S��}Ç�d��.���f��2��~x�`i]�w��N��k�ÿ�%'ԃ��;��D���$�%�! �F�ŶPh�n��o�*{���+��J��i	�!��!v7���s�AS-�giQ-/�_��r�s0N��V�hUĞ�Kh4͏��ΜZ}�0Rz��$暃�E��[��>7�Z���'��*�MY�c�M$�u3n/���5a�<%ד�����$�|�f(2�M��P�ѽ0�G�і����7��%�Z�=����;&���]nX������<�ǉ����2Җ7�GH:%%'�HE���d[�`v��6�b��[a��87U���oM )�h�Rt�(�n�(���F�˟ƕ�Q���V��64��%�`�5#�4FN��2@��u������|2la0�M͑������BHy|d�6NTj4��w��M�r)C|c���j8G����/�|��tdwyσU܊��U�i��q����	&�c�ة�D�;���ѐ�G���6CX<�`�0r�O�a���C��O�.b.����3���ǅ�-��&k���;l��NBv)�F<���m�xI`�	�D�[ƾT5(����ʌH})�|������9�{����D5�r}�0^ʭU�y��G�mV��]�,��Qbr��3�95��s�:�g�֋��xfs$lD9��0:gK.�g�(V=��ਐm�]g�u��3s:�k�'��-��$�K�țJ�I]Ċ�bE����ccY��)�9�(�i�����N���xXvmN�1�?�^����g�(I�>�(���h���A�#,w@����f��hhM�����1���@�g�Ԉ�^r�����~�
}�q�t��D��6��	$b����X���}�)Eq���!2 &��ywaC�}|�����h��lM;�pZ^x������l��դ���Z�z>t�C�n]� �EIP&�����1���F�۷*^C��X�v�*u|���b 򗓌�sg���)�����un��`J ,��c�m����C��=n��TH�:�T���� K�;��br9JѤѿu�[���p:!����=Ca����Էn������=���+�»M��|�Q鲂���A��j����2����)d:X����B蔚x �k�Ϫ� ��ϏG5Z��_p�DI'��:dT��ۛn�'K��hs�����Ϗ�ѹ��� �DW���#j�s1q4Όy_��H�7������'��kA�0�����ek.��O�B�f� �B��&"vS+��!��`�Z�Y6���P	&@�P�=����|����p1�26��Ȏ��A%;����W�>YmK��?]l�7ٛښǨ܅e������H�MD3����ᎦC'�����Nv!n���̥�lv�N����.��%���W��[�J�/�&�l��-�XSxXC�P��oF "9v���w�F4 ��4wD�[�
[�5L �y���W�7�D��{�N6s�t�Lv�����G�9t���	X�X���^�F
����nh]�}���5B��3lp�ނj2�Ujw�HC7m@gM>��������g�3��U�+�xN�F�e�`�C c�{\`�ͭ�?C? ^��T
T�-$:2���,����ڸ�F� d蚁,�@�g�Ԉ9�Ǔ2�f��j���dfoj���L5��E�/�;̅�b�¦͂��=;�m��]�Z@�i�O����4ܘ.��o�}j�ӏ�)���&1�vn�S M��MhH�x~������s�T�*<�Tr�zM<���h� {���,��3�[��ze�;��b�Es�k���T�-bŀ^�c[�@t�>0���"4v�WЩ�9 �Ev��M�k����Up*^Ϩ@M����Wy����zo��lpJ3����tG�`Ha}��CG9�@��y>�)�����w��;�C��h<Z���Eg�&y�.�y�98���"8�j��w���g�JI�W���$�^���	�s�BwK��z]+�����T!>]�ު�uu-9qL��w�+��LU�#��m
i��u���H@��BHWI�db���re/��+�U����BW��s�uɉ��ҿ}VIf� �>��� SP�:q�1�Dg"�}�1���-��ځ)=Y�árB~��Z��Bd?�P�3 {('cCh��}��i����K��N�rީ�ﺻJs�P�K?�WgT���D3�s�3���B+^���}Ҙ���~*�Sås�~'��</�짪gȕ��``h�gp��R�����2����f@'u}����+�9�D�{�<)��Ăr��\ʳ�6�1�,�m9h��!�R�	j}|�25%8J[Kt}�U�+����W ԑ��…��f����:�cA�m�$à~���5�v���m� �;�1���MN[���;���Æ��=��v���0��[���+���F�/���[a�w��Ԕ��}RP��~4�6hr�m�u(~o�JA�p5�]�鞓��k�R(:�!�)հ;��TŠ�Rz�A�������`�R��#N��	7�^96�>���1=ʺ
�C�hA�.�y�v�ޣ:�x����@�����z�A�����@�|u�'�s����"�C�̀F����g-�=���ؼ�{�3ެ���aG%̫��	�s���u�o�Kg�#���L: ���z"�� ������~�C�r�9#L�P�by��/���:�~�➐wh�+���j�8g�
�Jy$-ފh�{eʘ
�WCn`���0���I)7Ȗ�pls�0G|�b��pg�{m4~L���P���T��A��b�4-#���R:��6�.�
��$�熅�.@�����+cs�{MO��Ѵ	3���ωL�-����*��g���wїе�<jV/B�����]��M�7�
]_���<8�ȋȔ��R��DP��3<����>hnB�np0]�@��c�$)4��B�Eg�P7����u�d��J�k�7	���d�yna.��C�%��&�+��%��&Z�{n1�H�	�a����kƙH_ƶe"[��T�
�PY�y�� �����Ҹ�B|�����W_���«[w���=C��e�y���ʱ��Ʋےg>VPS������8,
�Q0t�6�2x/aC��zV~�KV7����~��y����M�e�0�:Hc�킹��ͽ����'��`����J@�r++� ��m�m}�q���$=���YAq�`�X����V��y͵�z�6��},_o_jL����	<̻���t�?z��t<8D��BY9m�e<�(�E����zF���L'}��د^W��/0^�4.QK� +�����K���*�	J��P��ppL�7�Xt�X�Og��>���,{'���l��
���H�֝iٳ��t�)8��g���Jy�g�>��r��E���{��z��Rݾe�Uϊ	孬�":��g�ND�w�Z{ߩ�� z�x{�[9T^>��
���Rع�r�����v#F��0�����d�S��|%��������`���s"⠛Y+�m�o�ӡZ�=G8FpmQ=U���:顝C��s�Q��j`Ö[9�S��rWx�ɼ)S������[3�X��I���].7��q�ت���(eH���9����e�c*��O���#(-�g��nx�oU�&�ܼ�B��N��e��p+U���EcL�]��U��;�"�3����UV�&ny����@S^�9ԋ�8*i����b�K��bQ,D	�I�A64"*�����J���]�`�3q�-�92����0ܴ�wD>�H�K]����kRL��o��hk�K��d��|�su��L�. ����9����wk�sPd���xξ��I	�T�6��RC�"-��/ːDˎ�i�D�[C ��ջ
pv���Q�:���B���6�R��dX�^��]��%�t���+ ��p ��|c����r��c��N�&�ҝ�B�����8�~�п2%�$Vq�s��U��'U?��X�\M�N�.�`�B�~f__���n�����k�Z�6������X�olP���]>��]���!xG2�=��z�$R�{k"��f��G(��3�u�IE��C��#���Ǹ7Q?I�q�;! ȧ��;o�9���A�Ő�!itr��Eʙ?��v���&(�L�*\WfR]��H��d�$������ٷ�^�ۻ�w�v�a�,-��J��:�B���ֳ*25��Ԛ%[�uѠ��D�꾎�[�zw�o���<c"8cr��p�Wc���?�l����6��IvZ�t�C��?P�l�Wl�DC�o���-��T��øL�7�aZ͘�w99���~M��ӰLDj�9c�֦9�u�ʍX�)��;�������%k�|��n�%X�i�5VX_E��8X
�Z�Y(&S��KOI"[m��T�RT-�U)�i�む��"h���n�(��W��g <4�)s��'G�Azn>�r�n�i�P3����l���W�D=0L7`����:Gx��-!(�o����hR8������ꔒ�0�@�b$/5�}d�/��-�@NR\���H�8V-}㬛�H��o<��-�Ƃ#:��x�?[�qo�ʍV�"`���_{�K^=��U��*�pWzc[I�n5z0�=u�fv"P=��P���|?k��w�*������zо�l�Vv�
F����v@HJ����Q�m�����Б��7c�ƈY]��.�8J�vR�p�!��Φ�q����e��b�V^ۮ�w!m0�	9&�Q
��]i�5W��8�fh)/"R����+R�"�������"S��I�2���|����A���]<�����<$�����2�9([�F����<[F���4dH��^-�i�+��U+ti�+ȉ��նm��X�U���s�߭�k�)��S6&�Fp�V�B�j�}ذ�|3�z�3�l��tT9�b8���E�fG�<h����}W���V���FE6��
Q�v� I��J���0r	f0y
��n���*�����e�>C~�-��R�2<d��}����?^�ڔ�E�l��l�a}YH��Ზ1c���$�7p�N�|���E�����Q�Å����ҵs�@6�%#+gw�v��K^TO����i~�u��cӢ�z�j��keR�FlX��ՊV��Կd�|R�<��e)�ޒ��e1�
�Wc�Pcq��K��^z%� 礘���Y�:�lM�P���oo+g:�x�����r��Zf�]U�I��N�l��NV�/�	(���ʭܝ�����p��҈b0�E���X��aR��Rf؀�S���ƥ�d�A����[̪�1s<Ǟ0
�����@��S<5�gJ�ak$4��C�ڒ�������pҤ���+s���]� �˥0`s!H��r[��Y5p��WB�S8�`������A��U������<_ؒǭ-���@���y��o�|Zc슈2���&M`�(�\�M��>Z:���r�% =ۥF�ܻ�&QhCE��&Ar@����e�J�O31�Q#��<1m��&@�Y�!ԶB�� �#����C��������8�0	@,�P*�J8p����O���UE�rP�(�b�9�β�t����4i�X�Q�C�.���+OE�V�W,��܈G�
==��o�GW�tF���{d� W,�e�Dlu�e�K'����h��t]cӃX#@�Ġ� X �!��۶�'HrK�H�-�������kʨ_{w���[��[�]�U���[�=-�D{�Auix��7�h�y,�`�x���p��!.S1��s�z�y���bш��A	ڦ�<�x�(C���}L�����)� 3������Hp�t ���6pU��	B8>����w=��6k1�Fц\���Y�O�G�Q���	��^��z��]�/�n��5/����]W���#���b�'5O��& �py��,�O�.��7@������Y2��.��]i�VPR�@ȥ��|3*wf�J�!L���7G��;k��ݐ~JJ\��6��A�O�H�I\�'h̹<��Y`|�/�2��Z'\��hT cR@P�Njs#����~B�?/7N�Dn��"Е�4�~D���@��!M�>�4/�㻰1*�� ���S��z��0p;�}*�9�@;��7AP%<��M���]i�-ZI�w�6�Fq�(�)��O���1����i=oa��+��8����/������-w�x�̮������]8�r�=�F��(�IVb��2�|&$���W��[�lf�2� ~*��|W���M��C�x6N��cRՕy��Ba�x�Oރ#�9�z{������ƃG�3����E���T.�ΐPÌ��Y�iE�곴�aw(����~���g�*UP�q��Ey�/�)X�8hZ�F�?�~�ΰU�V�����R�YDS��u�.3�|�ya&�i�
�����6;�h!^
MR�v�Qr�@ہ�!=�QEJeB��n�8��i��+��8�Y�?@3wb���>	yjkE�ߋ�pB���T�a�ؕ�A`���I�l�p ֜u�B(�I3�H�$t2%уXX�: �0��(jf�%9�k��	J	h�\Ȑ�y똌s�ޝ�����{`��w��~bc�R���T�w���Ԯ
X'fO��k!Ho��U�V;r1���%�C����n�^��.ޱ���o�j~ι�8p�d��f(�;i�)xI���8�����Ա#�a��1X�.S���b
|���C�G��T7�q�!�����P��@G!�O��њ�s��t��#$S�{i��!�eA�tf�T��R"�-��
������'C���k>���@) @!~���7�s�7[��Q��D�1=�D]��jSK'(�q�]����3�Q����
�I�'�Gv> � 2�D�F�c����IQR����`J'��V�p�������y˳uu���{	:�]����n=U;��3��s����	�Y3�1�̓=J���)�崯c��oh=Jp���3K��<�й�Ms��Gj�-����%�F��:#�o����`�G�g7�dH�B~7���rۍ^l�|j䐢UHC�7^ZcZF��뎚&_�+������B��r��y���t��5r��`F@��V� 0����LL��
���a�HSγ&gog��v3;c�1�r�K+&#\K�t#��t>�ެ���4;�f�Z�b1�^�l���,=��x�Nz���ykSO/XЯ�ww���&�� ,붥5��_�*1�;��k�|�
����Rn���ſP�N�.9�z����(�i��o�O��(�����?�(�}$>�	��	�Xb�u�[i�<Y s��a�\�c
ё�v����qOO2�C*�[��ƨ�q*I�P�%�Sd���C�^GU~uѢ\$�+��/V�O:�BP���d�ư�Ud�d?G�=���$�^�'�I��6�#�G?�ʘ%���C�S�HY�����nU��Ǎn h�5#.�<���}��#T��ɴ�S�6�Pd ���!?rmm������>d[	%*S�Jq ݕ�*�G�֚/�6!�1�&R_�*�8���ع\��d�ܒ�)�}ơ����mT:]`��f@��d<�"��ʙxW��� '��l��e<��EHX`�mb��(���X7��S�٧�,P��2k~���X)�_���Z�#��V�]�$���%_�'!��,f�S�#�\CM����m�Ըq�i��v�;�Ȋj�~�U��#��y{�@�@���4@yŎ1j�UkX�i�'�N��MO��@�ճi�� pO*F��(A��}�SS�CJ\���YN;��M�Z�"N�N�m���C�`\���z\����
�ީ���?,l���	��{���G�+(�h��
R�/�]D�������O�#�mϭg�i�]�~���0e�GJ�"�C���[Ԁ����ߨ_��$s�<���n���/��'Uð�����9���^$�zw��A�K[1�`�d����;]_d�Oz��/��lZҮ��@�v>Fq��KZM�e���.�o�l� u&���*��'<���=�8N�H���T�����usTf�n�a�)��v�J���g�*��n��d�r��'63x�����?B�6�$H'�K����*EW^h�k��M�_3W����Mp�g�u	��\z�rW-K+�is�+�2�����a�-{���Z�k{��x�oV�\�I�%��5%���Ł�A�(��`�����`��w�`��߄�du׾��_x���
�nXk��Jm�h|=lX�Z]�]N�h��Q-��[a��tJ�+Xe=���E� ��t�̟ټ�ۂH���c�� �ba}�!(}�L2$�c�u�QQ������Y�ZyJ�!����j�]a[V���u6��d���
aR�T���D��R����eK�U#N�ɼ��Rx� �I��3@�4�ú����\ϱ}��8�Ñw�y��*|�-����/�C���U7	5D/c�5�M��5�iH�J�tHaT��{�,W���(Pb�`���IS{��P���@��YL�]�����w��&����呜ffőU��?PhLj/I��a��mV����b��Yc��ЀQ�����e�s�t4���.dg*ᒖ�g;���\�d������5&���0�t�n�	�Kͺ�>wa{�t]>���6�N��0~��Z2?��˼ֱ�<�r_�I���2���ư���-���d�G ��^J#��J(�L=��
�Ap�.I�3QsR �G�3ާD&FH��KAs=U��5����~؂!iP��B6�L�c���܍9�����;7��赺��l��#G&����q��g�]�� ,bm���_ː_~%��@p_̽�4�cY06L;Ȏ����������:G�36i�l�����~־Kҷ���;���dgi�C�\1�0�::"�����v�ݓS�m��t��������?u�V|5��۟���[���2���r�6H�y##�_�I������~疕)S;ڗ�6�X��x��
9�*M�QMܟ���\�1�#��-T��hX¢�E�,�S���4˅|��*��=����+v�֓1!R"�ȱ��F����l&���s,����X�A��Z2�.̮��E�!�y�qA�G�]��5%�ga��X��5�+P�R	HŏT��[ #��W1�[���D�a"Wd���厂���?��,�t�93���m�C8�Q�o�~�-tz��_��� ~(�?�w&>[s�-:\
���BTW�8׸C׿�Z#��#)��;�q�	^�¯Y�Q��W����`a*�\��M��Q�4�dn%�۵<p&�*�^\�58��t	v����J
����d!���z�cq�ʵS��|9Q��7�bma��j�\E��o��8\�&�_t�6��_as|*��1�h���~��W�j�a��g�"���^؛�X,����Un��&���H������D��e\�8��$b��崬�k�֙��}M��p;K��'��mCr��3�A�*������6�Gĝ�i�sIv�r���R�B��@��2�\�
�q�qW�L@lm� ���d��n��>,�:H�ŘHE�&����)�(�Al�:���M��ת�qw��U����*x�\��K�q��`�5��x�ԪC0������=9;f@�����	�x�lk���|f�-�����o�\)�f�b��9R��S����_�R�t��C�h}8&�_e%��y

>�������i��PM7^�<��(CR�^�r��c���nZ���^	S�J�x�j�E��Y���M,��.U�$��������N7��	�:����s���={��%b�:�!�%�C7�د�p����I�#�+N�e3��7=c>�|qnK��{������AGW�D��|�P�r;��~A4Y ���'��;�x6��6�x��b~�D2�#y�.̍�V~�����xi%I��P&�&�)^0[�ꦰpG��>F2��( |b�R�>�k���Gu��_��k�w���z�4'דc?���98�E/��ٗ��#^s�Ӛ;{+�r��n�~���ݙ:��v�q�����\�)N�Y��3	[����ds��;�p�wbe�Qp��t� tN�]�x�/Xvӿ{AG��^u�03 Z�g�|��.�.L�!���]. -��_b�_L��bj�üXE`P�K���0Mb;��)��>�Vgn���\�~3�I�d��}�LQ�I8W��������f�!b����֙P#,?H
T+���0x�2)
��P�X'~g+�~,�6���u���;^���Vc�Q�CQx�e�4��ԢFE���$�(<H���@gb��/q@������QI�e��Z��C��VӪ�֬� �щ��PW�kpo���ހ���D�tc՗�ɶ�PiE�;c�K��6�5<~E,�$@lSƫF1qZ���|��+���z�`�G"��/��gJ�@�k���i.��EC��#C�~��iY�#4���l[2
(��aq�{�)k��_�ٶ���t)E9I�ԚQ0��ܠ�ga�3���V���_��(�ՠ!]i�H�b�q�y5�/��՝I��lM@"�M��Ih��14��y�X�jdZ��h"&�'��&�x���
��|�#���'� �XU�MOTH0g�e ���?�O�7���ԓp�h��8"��g͒t�U¢Gq����24������᭄�ѐYS�gB�[i���,%���t#Fhh�xz�����uڅ�.�G�*�+�ڬ��7�e��p�}����S1�H���<���.��F�3w�����
~.o�^��b��Ow!\h4^�U�˱��@#�q�eG���z�6֙pk�֓���K�pbFX\؍Q�����������N���<��q�i��N&)��c� '^��CE�+ԥ&���b��"MX��:��3�&�/U~���nx?�|�FdēƳL�@�N�,1U9�lГ�Y�-��B��N�g���V�L\:��AC-����Ts����}LBs=� ��,N��./z�@�`�j�'6az$�73<���=����2�q��Jd��ŕ1^�����%�4f�H*ᷞ)4��D��1ֻ��$`,���a�s�(t�V?m,;�.7: c�Z�jۋK�Tr�:P'Uv���@4F�n����M�èP�iFe�ϭ11̣:��x��^]���f1��hѱ��x�?%rϒ�8p	�����9|�P��3��a��!��z�L�Z%C�ھ��x�&�ߜ���#.�T��C�}X�C��𲾁��Y�� ��,_�{@|'�2�q����4�aq���,���XzVC ǘf�O�ѩF����Fr��4�ѧV�J?�. m���h�K���1��:�>��;��3�����U�t]��� 4��Gx��U�k�q�Er�=y#g��l���{��`��+�Ⱦ@��0Ǧ1�";�Y�~�Ė7�J*9�L����Z�C&cz�BQ"��<3�:}3[Z?&��8��~�gJ���T��(t-��u3����ї�}�1��X"Nh�{�L��݅�s�ٯ &qt/�3b +<C�sE	UN�*�tȒ K	�fF�4�9�r��Mv�J�ҝ�Վ��ߔC�4ڸHz�� x��c��a���έ�gVK*�I���Z��9{B��_[���k�f��x^nVb�n�F�z��e��F�}٦S	Y�}0�n�~���)F��qd����=̊�Zl����6��$�����k���D��c���^oخ4P���yphr�l�_|Z�enGn�+�LW��WҼn��)�7���<[�F:�s��������.q6f��6&��p1-��2���9$���k�l-hPN�1�� ��	�-�5��s�R�g�\�:��1���n�UNJ=Y�^ծ%�#ê�O0��k�~Fl��V�?շ���o�1�n��A��!��o�!����o�j�����;��&e$	��?�Q�r���0��m��g�P��l�x�$C����F�W�2ffm�=��u6G��*'k(�QE��U��0(��}�]�� )oŅ,�0^M�Gvq���Op�S��C��<�X7��ץ�!�
�h��#�<ғ���\��L��eJ't��Z̢?�ɘ��3 ��2�(���Sͥm"($2�	!ꂓ1�I�.K�F�n���O��jխ� ��{�\@VF���3Y�I�9ә�mn���x��."�	g%��A�s�RB��;��_�M��5(y�%�Z�u�I�m=�m�S���l�jّF�x���;��qYĭ&�	�3�9QW9^|(��ZlB��Y'l��=�����ĳ����#�����Q���7���pŐ�s"������%~So}���4�`���k�+��� ,��4�Q�����lw�]�z��ŋ�c�Wjȿp��$L.��V�Q��}�t@�:��+�i�2d&>�ɕ�5�U.�4��g�Z�TB���Ӝyِ��]Ǭ�؈vو<0��̏	q4�z�����_ߊ J��y�
�:�"��ЙZ������+��{�VuXr��\[)�&;e9���U}Sݛ�!�|�u�NUPE���I�ajF��]���]{�!N6� �9(A�R��`�H�������;�}��cÉ��iV<V��^q-�2B�)hv���׮3�a4iu������K-���<�"�#��{S'��C�����������f�ݝ�O��,�}�ľ�ul��H��M�A�.N�f�Ti���(����^5�맀絟��ԗ���i��	<�ⱷI��<�!Z_�fi8'��
���QWCT�}A�?<^3/ U.[<X<��
ܒ}�Uxo�0r��}{V�㝸�f�qz�dg=s߀��q,t���6�~��:)�����yk��.~[���l�R�M�w���+��b��� a�j@�H9߁�x����������(�{0�]�!�%q��%����ĵXD/q��2S���������l�aH	J��!CU	5ϓt�|W#t���@������,'�cffu��N�`�O���>LO$��	�G�-�	��Z�+����:�|����T��vES����ieR�?=@m��b����2�A"����07tɢ�w�����������f*9U��H���Z�n��F���N�jrþ�f9|5R����<�0�p�t�r�
�������T O�7������A(��R�Sv�/1
�0"E/���< �����4��&����%-�:WU'�[��(�9m��k���vTo�;�q�E����N�e�8�_< ��LPWH|d���n��[uLg/�����	}��~��'�.LJ��������65M�@��7;������˄8w)}��Pv=��x�v��[F��8�i�"�~O8:�a�^h7�w�A��C��f�b!�|}�1��!�U4����ɥ�̰�����*�$�]<Km=�~)�M�-��Z/s)T6�G� (�����~��ҦG.��P��W��Ƥ,��c�<4^��p��M���VD����!��ܲ�,9蟈����A���/���uy�!�db����;/(N����C�~noȬ�zEc<��	�9e �7�B��;U�|u�|�N�@9�fdX�MaԘM���<�~=�S�t��>�T]����C�A  ��^t[3�C��� D�9HC�/7�j�[�ˡ�+���g�ms��_<�Yt�yf�'	x�ŏ#��S���|X�'X��,�
��Vw�+��-�H��2�����~v��_���͕2��U�K���v�O����!�Q�lj��O@OK@��o/G��vY�:~Ò�ڕ�XR�,�ѫߊ�W|q��F����_�Q��ä+�J�Su$��p�.�~	���|�t��@�	}o�U�ٶ�� C�zf���f:sL4��M�-xow�(�/,��X�S�e�Q���'��
V3s���p�|�ˌљQ��9�7��3	?��o^b�o#=��ndO�d�. \����i`���֌:��#(72l`��SD&ѨT��R�N���n�ݢj����?��^:�߲��Q�u��|�( S;���=�Y�"VyIc�"������L}I���]";�;���,���Q\�[�5<p��!R���
(���xx����j<dBk�Ac���$�SRHyfS�?����TAB��.��W �%���c>���+���|={Kۀ�Т���K�<F����A���X��2+/%O8.��j�dMp~
��z��"�_A ���v�Z������O�Y�H}W�[��{|��|Nk�p=c4B�����e����U����������bBi%� u2�v7�@���[�1?�qUWLk��;/��"���51U4��H]�i�%U�zE�}�H}���	m��I`�;���L60z�К���lz�048d&�2��u�x���QoLmf�����ٓ����~7X��(�z<VtY���>�g�	�׶�NC��p�ypfS�����<�Y��Ϧ��p�sk���A�\S���7}t-M~�юX� ��]�&C�ɶh��4{�k�#e���	eָ�壻dMv��=R��0E��	����^(�0�UB�	,8�����.�y��P�
C4���e��JĈ����C*��:��p����_o1}%Fz���-c�S�+8��}Ͽ#d���ز�c��m���&�x?�U���$hk�v����K�3H�g0Q���b����T����o3��C�vY���+�Q�b���M�ヵ9�(�S��l��s�2h����WH�,�s�[�U�4���-T ]���V��p�	��O���  ����8�QTW�E���!���q�y�=@�ɚ^�q"Y<�$>����1U�i�������_v����ѱ�ףq�*�I|�]��ɐ��Y��
[6�E�5��.�M��M�^� ��d�1�|��v
�����)�g���q��N,#]i��pqʱ�]h&ulT�%�צ4�6����e�g����YrYr�f�(Sq�5(~iu���]0E3������w�c�{w�n�D���f�WjTp���&���c�7�d{�>�\�[/)��W�T4u1'J!�)fH[ޥ���l�_	�p*+�Ol�Df��3zЯ��"�.�a�Y+%�����bO�����U��}�LP�|3ײ�c��8��V�;?-a�V�B����kb�)II�K�ɨ���'V�ٷM Jt�ǈS�m�g�����J�C��jo�Ź�j�YԮS($ө�������ğ����� 6b}���y����^28�*M��-y'w	�n�.�~��|Ȼ�O$���A����D��UA��Gou�4#�_�am�K<򊬹�U�����b�9�ދvn�7�|�B���A�{˨����V�>Zx�����\z5\.����*��v^����7�Y���TR|X��:�F����O�����E�a��[4�Kǡ;��"dtN��pmI@r�/;}OI��ɑVWXF�����Q<�,��}FB��)Kբ�bK�]>�1�!s�#2nx!�%%���t��z��|�gax�#�l�^�ϣz��m�@�&���� ���#�4-���>f�0>݆t8qT�I���s~\w2��;�JveP�8�oT�-+R�|<z6FԞ�F1Xb�N�\���_��A�'b)r�Wت0�8?qc�O�r��L���N�=|^O� ے���ɺk.o@�ٶ�N��=뎼q����՟E�+&��͡X�sU�Xb��D��X4_x��~��؍�w�yH�d҆e�h�QR�2a�)>�$�؈]�VdV%���W�L��5��ҧK���EV!�pq/j�4�_��J���^�m�·�H���#�p]����\p�W�>�;Y%�������>�T��&��⹟j� �fj�?K�� ��DKA�Kt��W���b"�~�۹uѽrB���S�K�,�r$Gl�i��d�c�5�-e�1L+Y�hm��t���*,.��N!I�������=��>�NJ]��g��e-�fĎ�Ȭ~����Xs�I�Q5\����o��+3S%�
Q��{�S�e��ҖWx�	��	d�j���\����]vG��B�Ё� �gA�X;8��܉�矕�o'�˞LM%}l(��$)��>
�Sx�`��_kH��41���grj$���t߰�Դ�t�W�|�Bz�9��R���\���n)���%�oo��3�"��Y���q�! ?���;$�S�_f��08����?��*�5�˻��XǙF�	6
�5]C�_^f��ƎoTRh�'��Lr�2�% ��mi��R���6#�^.=�5=�=qh��F��I��x}h��3oh=��Km5���΂�_�M�U B*���w���I$���=~\LxHu�8�vc��J�@Bt�W+�QE'�_��i�����1|1�w�j�8��J�m ��9��yX�'��{1z��!�:��(�:z�;k$9ɲ��R|w��� �ϩuMr;#!�.w���E�z�F*��V*��D�O�or'�0�A�]&�ʭz's���8��
��L<��Ψ�"��>�{X1E�S�q:D��N}ȵ|N�:�3:w�����1ُ�A�d1����Q�t@yha��a&�V�������x��D[�p���X]Յ��&�8fغ_�32�$�a�-kTN/��.�8���މ�K���A&O�4��4�	DC�7�u����'�H�+��`'��-�ĀG�����(�6%�dLc�,#��yw��3���>k�ӫp}�}x�S�#҆l��f��A��y�S�zJ�7�
�,�T-"��wTV�2ˬ&�z"�r��K	�c5[n^1�AK��_�o�
�B���g�5���?�^=kK�����۩Ӡ�y���~y��D���D����e��G,�,���H{���54m}��1�i�b�h�-�"	�-�I�Y��AD )z�H���������I2$K�S����2�9|�`�:u��r�n8�IϺҲ���I^�+%V����0 ��z
���a]��3	�/��Cc@yb�J󿒈g��sSh����X=��幦�@��W$��Vg�x��I��+3�wЪ�n�0�x��y&#0�_ߕ)I
�]�_�?(&%eQ��k呼y�m�yzL�����$��}H��mi��Y:��)݇ �x�o��t,�<�#����9�ʪ{�@�S��.p���"�[ڪj�M��)���QT6�3������ٽg9�)�P18��dh��W:,� .�à�o`3D�����XP�b;r��4�!A'��0��J�=�M�%%��x������P���J̔������^Ίi9�"������d�-̤���r�����!}��e���"a�0�sW��(�H C*T��ԛ�'�" ����,��uH��>���B��/>���Ac�X㵶�4 YbFmh4[x"&��7��*�c:C�a-c�S޸�P&���*%���N��@�a?H,nR�����1}�=H�s��	MV����CH�B2��`�G�_l�n��xq��8e�:x���.�bk$�6A�A�N���L!�ޘg����2!�����^Fʷǽ&f9�ӂ٥�\JjƠ�_|�mi2�ϖow;̆T���b�9��aL�-�2E��je��O�i�(�������I3ȵ�X�觑�
ÀM� �je� ���k0�-�疶�(Y�\�����ׂ�aмԍ�Ft���2��)��-I�&M�Tg�DF�OR��A���{,��ƴ蟷uY|z
�N#��Y�xp�42�� ;� X�N t.�n*_ T���*2V���UM� ����Iʷ1k����[6��Ms��j����[��~��x@ ���R _�3j�@����ۑ��p�9ps�;���@���&i+��Wa*@� �N���NG��t�Ai2x7�e9!+O��G�s��A�ؾ��t�:��@�4�����<���Y=�����;�6��%�+ּ�ض� 9��0X��Y��f���Nh��ŝ�Z���h:=D����[�r�n�z���[a��� 9E��v	�t�h�i�g�κ�i�u{r�r��I�Q̰�^��8��Α_�F9g����G�oҩ%��A`rK�V����Y�|��5䥏*:U秳���h�-m�$�M��ɼ��w@b���wJ(T�&��nYz�q��+�|/��P�<�0���_��h��/#�H�����]��+5�nV>��=>�`��Q�O�⪜����b�W\q����ՂN`=wz���Ҫ-�ᰎ[Ӄq�vهe?�p�p�!F�oW���;�����WR)�	n�Doz����Yč�zs+�i�(K�3�:�q��*kd�Bɞ0�֗�^g{#�qW��Hwn-��~sQ���z"/�*p���ںhO��>��v�ߠ p����3ʜ��4�;aqǝdf�n<�8-f@s�D�ƈ,�aO�e���5
V�����3#|��n�I�c�]j8�_^����v����L����c;O��$��7�a0�y�K����L$�BOV�<�A<i�Ix�,OC��,���cX�k.�Ζ�ύ�?�G:��e�bB+ʩA��	����'>J��l�k�v���a���A���Լ��B�ꜣI�y��rf:��X����x�u�Q����e�ԾF���\J��M �䤇��Z"WX���!���'і�FU.g��T����X�'.�E���H)�F�+&���p�h� �����cQpg"����j��wۥ�V��hH�-�b�Gs.k���y���VQ��K���u�Ա>�K�J�����IvwE+ō�H��2`�SN��h�>�_�����*���nb��+�tJ���kv?��Ҿwl	�L�~�T$Ob�ɨ"�Cd^;���������1�����s�$L\=Y|h2�[���b�.M}Pܢ�݄Y�����6� SE����F�
� 8�ې��m��Sa��,rӟ$��!%A+�C��o΀�Ӂ74�� �j\!�դl/�M��V���:��C�|�_kD�!��<ͦ��j���!w��;����ʑ��U��xi,��b��ɇA��B�6�y2erհ�4l�@|�Ѻ��ɾ��ɐ
N���_w;Ҥ�&���:[�%�6�������o��a&9jMj�D�&�o�i	ֽ�&!�yϔ����}�+����0e2��a�r�u�H�2��E�������fw�Bb~;�.B�`�fh�J�d���f���3�g�Oe4&kW�ⰷ�E��Æ�r��.���l�l��7Z�W�'&�P|#���6k�f��#��?Uh�;��	�3Ú>��T�E�x!����gg�[����9���@ݟř� �oc�&|nI<�>�m]%�;@�Y����)+�IW���	�c�Bc�Ȇ��EK��?�)����iP��z�P�?N��ش�|��,�)�����^���.��9-E9�t�jL���u��R���b%*�1eLU�Lʴ	gٝm�}&�Q��j�a*��@1i��F�F�CW�"�8*O��y� �]e��!��ke�bk_� �C�<�-F@�.������:
�'�4[��2&{��I��{jW�]틯.�H@B�/��
wSn�z��a(j��R�����r��t䭗�5��A��^`a �r`Ys4�S��\��IC�ܓ$ ,�a�a�ZJ@���JP��z��gL��Nr�C[�V������X�����y��;
��������}8`��I��=5�=�ĲK��@
��!q�<�-O(o�ɝ�}�5������_M:��ы;T�
eA�_!��3�P���~6;p�x� �9W`6�i�4�w7���[+�?�	����7��V��	��'�"i��iy2<�J�~����LI��;��#Qi;s�O�䪣�ъ�K��K/����6:Z-뒲�ϊ;�;̺��!14!U��8&ţ?ߖKN��"Vgic_W��y�T�M�%mU%�	k��!�ϣ�ı�8�E�+C^����^�mM�xJ�3ѳXA:�j��p���+�bv���s�[�o�$W����[�w<p���c	�����U��o������٭��9�S�/L�$:���K�R�����b�e 3�Fz��R �)��h�X.�,?���W�E[�; /�l��:�d�1@�"	{���
����@m.�d�u�9��Q�W��܏����`�q��;�&��Pt)"M���DBZ���*�vL}<���5ai���Ⴁ1=�}��k�)����<��y{�e�(\�flC�-2�*���uC]G&c%��g���/��D��锂�F��<%d�qWU�GT.��&�Pl��{b̠VMO丱���@� b��q 7�M��}\t�&������$J4 U�^p�/+^)�Bڭu媖ц'�B��Fm,���������I����Sl�f.5f�����,��<��@c�blw�lNo�}mƀ�Tϛ)�f
����Z���Ar��5���a��JBh��H����T*s���
��$?�)�Z}Y�qg�\j}�$�sT6�`��]�ᨌ�рՈL*�lv����[���{M���Q�IӀ110^^ܯ�q�p�J[��sĲ���U��ݟHs���e?:X�v!e����t�)�����\�R�Ω^A��9�j)(lFEb�^IIH�ӈ#o�P���O���F�3�\Ӆu9f����.`��0V����؆:��9һ��۟��{�oKP	u�x�QPmH@��f���Ccu{���K:���ڭ�i�_ɗT;]8���`�L�i��'�SS���>�a�#�����͂��8Vh��LS1���r����\z|�ۜ�!�\%����o�������w�h����q�u��3��R��8�3X3%v��_c�����R|.3�1m���Z��2j	
�+<�{��3+��*jC�M�_\���?H��&�Jտ�ݰq(����N��Em�L��(1y��Y�k�승�M���[�L+�F�]�m)̩
&�����#n�a�"��b|P��ar�L���%gɂ��P~�w�cp8y|�5e���P�$,���{|�j6K_������p#E�i�?�8W`b��!�_�pS�_&��+�3Jհ��I�o��(?P��|D����	%���6��\���c�՝\� E��%�d���!$ ���W2O�P��͓�du�Ϧ�����M4�ѵzb��Si�@_�Kmq��qE�C��B*����,�)�/?�h��	 `1�Q���L!\;"��P;�
zI��p��0ͬ������G���.^����C���|���=������|y��7��.kf*j`~�f�b��I{��'/H8*Ծ���z)�i�!Y�a.|Fzg����Sa�R�B�y
�p� �w�0i��2�A�����Z��qo��Hٹ1�����D��>�\��SN�r���ců���D�%�Qu[�x�bk�E���,�Z.�z���.�-�-qX���~h-
��sO��*���μI�P[��g�N��6,~��)�3o6�t��JE\u�FI�+�����[KoJ�G'����x�8�kq�.�f��ڛ��O�Y��@���������VtQ�&,Xqm�/9vz��g�^" �(v�bTHR� A:7l��	����L�T�bZ��Oj��1�檜�6!�J��N�J�`-�ٗ���MtL��f�5������὾�fU���}�F��4�%��v�B���6����1��d�2�D����G��N�w�`�A�n�ܝ��I�����e̤��(�h�8���օ/����v����Ae^�R�n��T���Z�����[��r^�
��%bL�v;I#T��Xv�������-N�y6^�n�r+2�SE�A7�>Y���I�*���_�N��Uh��a���#�ڤ�y���>K�6���w�����0�r�֎������҈�$	f���= ?��Nß�� �� �և[!��p�ϐ;����z+u���]Jc!���Z4�!C3&p�h��=�Rm�߱�u'~��L����1�ڪz��>C&#��R����-�|q���@h�j�78hh���IA
��+�ƿY�_�{^�ˌ��%'ݾG�.��Z����J�b^��S/�����aś4I��px]��*�͓d��.i�8y�L��x{8�C��sTc��-�=����[7=����-��Ww-���n!:�F����o-)�ɰ�&3���vD�'K}i�.ŔchlE'�0�$�;|̾CNt��$��Ud���Y/I#����$�7R�Vx4md�� �k���1agń�ߡ3�Z�E����� ܰ%�	���w<�&������� ��!�K�x�?Pxl�3=n�Ej�;H.Ild�b�d�����'&��	�D��g)��+�j�g2Ca��Ey`��"1��W�p�S;K���u�R��x��6L�����n�ڣ�\�t�U�,W(��"�}Ӥ1��$c��JdRQ}����0��NM|ҘP]�lӐ��%�l#�x	�:����[�Zo�����Ќ��p�̿��Dw�!�&��9�+1�� �1��yy_+.`#
�r[��~�{qZ�U���O����?�7��y`97��8������s����49|t�%����R|.��\����f���|�������u+�$(�ډ� Vk*
nF����o�H1O�6.��0/#oLy�Z�bk�՟&,-�v�'��E&H�$��e�X�$���u�e���cǑ]y��W��y�b��(���,r������hC�'��2�\��҂��}/;~II���"��61)�޹�b͊������JW�g� �O�ÿ�2v��������}"9�p�ɯ��#�CC���*o�'@��L��2S�?_Lb���c��l�fu��(�R�ș�Q��X�[+&$,��CG��>��5�y��̨|�I{�8G���Y�L���s�����n7ۅ}���OL��Q�a��"�-����Bp�a�;Q:V��cA�n��`�H�Xں���SKQt�𽴬�W��%Y����@��8<s���
�kj�=��I�m��9��#��#�BTr�F���s^U$�����x�(��	�l^�݌y��ҽGlw{�}5�pG�����	ZaP��G,q�[���`)��Ձ50 �a}'�$��9�ڤ��|P�[t�������yE�M��I"�X�-ء�|WlzέRK4�l��P'��=SȆٚ?�ܶ�{(���Ia`��K�+��������\v�������-�Z�r%�����̽u.XU��K�U�TKM�t	��-d�$���k�l����|P%ƚ���!-��V���l	�u��sd��x`�N�>'8�+�;a*~�8��k��R������ �|����z�6�x��\/Z]J;(�� ǘ��:#�a�.,i:��t{��'a���B��2l��������\�Wjt���d���!g���� ����f��ڕ�`�[�iNM1?���[�8[�aCua���������Q�J��D�?�i��XʎUd�Pi�ü9M0�DM8��+�<u.�뼰��ja�#`U1���C�ǋ���l�`L�P��M2��刹#5vN��Y����0��͎3�6�q(B�s?�	y��Q���-���+G<SICˆ:�U˚�.N�<�W�X_g��(WO{�#yf�P�Z2(1��e��%�ՠ�>Y%/��`�k�jB�&��+j�U�Gx����&�s���EO9Ԧ�}�q�M�KC7]�>��Y3��_rx2�����F^��j���b��q��f���� �FTRj-��(���Z^R�/�;m�)& ��D�P����Qv�}M�<�b���	�n%,��nʊ��=`g>OLz*QC|&�
����+4����SD�3���E����P��<Ȇ���[�x�cbڗ,�kea�<銽yS�/��X�'%�5J�5[g�.2��:��d��6^�.e�bS�Zp/EW��9ʊJ̗{����{����}��x�c��;���D� �X��S������꧜�������� ��������͔Ó,���7r�^>>F8ي�-�8֮Q4,�=���� ��-���X��oԆC� ��t�I.7r��N�%�K�Mn��ǅ�e����)p��/4�b�HT㝤�1_�'�ߚX����7�F��]}m�,7� �W��.VzN����8��}��R,��I��2��LF��d�u�ui����O���{���j�f��&I�1c1�u����='1E)�`i����B��6i���;~=����[=��� �<�Qxi���в�u��<���!��*��͕p�?{��p��GZ��sGh�BHafX���"��vS3J-\ƃ�!m�C����ԡ+�3;e�"֕�\��(j
a���ro�i�o�e�[z��]��~�ao<6<��� ��Rg	 �k_������4M��@(^��u`p�}�
��Sjk��r���>hcR���!z���Q���<��,#,Ǥ],��2�\�w�Uw�hA��=�>���T��IΏ;���!�=o��|��F�#�FL�`r�q��ce��c_�{���4=5�0�T�����]a��~
c���=f�Lv��-�HLa�ڠ����6�Ary���ߴ�l]��_�s��6h��6[���N�ʈI��X����p�t�Iם�aQ�)^)���&��gәFY���G���Z�DEF����eFմ��J^:�����i�I�F�E��L�{���N�p��G�k̢t�Ǩ!'H�M��`T�O���$��m�>Ω�B�.�A���c�H�i�}�W���@@3V�ʉ؊v�����y�E\�Ω���%�>�0/J�vlC�oo"�wޯu� ��P(����p�T�t�3x�;,>S�N?6�5qP��.�7'�`fc�6YНK�^L��~�́�f���	�rX�qĪJ��o�cdj���m����*>e�@�iw��eF��<y��?�	�=���cMw�Cŷ�N�޵�WKΖ�Zo��-�P�����gJP�t�]mW��4L�9�"V�\�[����I�nt6��G��[����vJ_>iv��q�z��p+a�&�X��-���'��N:�~�I� �[�Di9'*Cx.�3ʈ�"dЗ�P�?56���8��'�UEZ�QUS{Ay��n���P��)����>�(�0ڰ[\fV&�t��2�]{�S���7�s�N�h�Y���G�\���A��xE��:�
��W�[������Sz��嘠B��幻6_	�[����k�?+��<K9����h�;�
�~��f��N�$
#&�&Q���Z)\���X0����I7��1�rBa�ףl��>l#��?�W�;���5E�C�͚��f{6��pכ^�2��z���L�C�k��hu샱�ٝ��N�Do_2y1|���>jO����A����sw$�#�cH��OUx.�p�拮��<��%ȄF��yt��r�� 9��%A�w���#7gCxg�[@,je�Hev�d�c�Tz�ҥ�k��*��Re�g(�X�s���Ut\�5$�����d�6&3d��AC8U�IM�Z2�1Z?&�lS���o�Y�H��
Q�i����)<·�5���O�����Ў��=���:M�W�!i�b�2�nJ��8�@���m$��w���gu�s:!:��&���s�B��ZF�F�?�����.���)�&{)~�%A��K�s��7�R��{���W��a��m[�$��{F7�^�7A��̋2# G�C�C_w s�CHFo�j��=��*ɍ��9�?ٯe4z63i'T����C�}]tc8*l��^8p�<%M�,�D���p׆�����C��`ws��,&��|~��M>䶑��%�9p���*ˇY^2�"���a�|�h��þ�AhJ��jv�f�5��@�b�����ȣdĊ�Z�����+�gH�f��΁�Q���� ��n�a�|�ZB�x�bK,��\!�X���mb�Tx�@� ^���K;5�q�����@'��a�U�}������l��4�0��`ǔZ����V@T(��I�73���GF�����ҥ�B鵡u��k/�p-)+)T����񿰠�2�H�����#fM�[�L
[BL(ԙ�P�<װ�A���:}�^l�{��O��&�#�X��)XU	,����t�q�$v���_NQq�g�@�4��YZ�����vkE"Rʀ̃�����LP���|���bO٤n4b�[���ˠ%���HQi靬_\��5�
��2T"��"��fd	W2��b�H{L!�CN��������^��� ��kJ�|v�á�H�������	m��/�I ����u\`"�1��?:Ci}��J�+�%���ʣ��5j�QJ`B6����DXѾ��z�'\�̴h�Bw:κO�
�4����g�㴥����(���ʔ�a����QKp���I]c
/!Q��œ�|>�-!HZ?t�>�-mA�l�5�&3����7c/�ڜH�J�D��\&��a�!��0L�&����IT��Ŋ�i��T�$�0khK�&�hHf��3Cڪ������V��&�w!d6�O^?�I�+n��0���	�_�(^g�x�2�3�ۚ�[?v�Fn�iZ|�f�p�Aq4X�TTM�+l0'i����,Ƣ�s��JU���1 �h��@������3 Y�Y��U�Hn��Ti��i��w�+�<�g}���$���ǳ?���l� p4-�o���X@��3��N��c]n���q0�ᖶ�
ĕk�%�*��h�":�$Q�����m�M��Cn]��]�hB�YZ��wA��b_�HjZri^a�K��q�����k!^��>v���R�����F��f�3x�d�b>q�<�Ln-��QMD��~H_�Bl-pIhk$9>>M
l�PQM� $8v��djP�����ly{ʟwK��d���
�H=�U��wD{
�W-mY�&~h���^e�>r�,wJ�D	���#�V?1������l��X��.�g��{�G�"M��	@��>���a�Z����l���V{p�������i��98{+�[9�
��O��J� �����2��j�?jYi�{�T��Rҵ<�zI*�����uNJ:�*���y����q���Df]}���C�(1����<��>I}�� �sk����8�3A����N�}%>*���x�����@E�XU��h�B�&/��� ����|@�z����Q{�?� �1�����n�mf�"�r��j ��� W��r��RO���|���,���]L���s/<�[���8[�7�V�q���^���IN�K���D& ;�I�aEh�� jU�q�k����-�!>.f�jL�jw��Ϛ�S�W',!�ӎx�^�o`�]�LM$��А��|�jD���2���(@���S�I�ӗ(t�Z���h&��_�; :�X�E�ᱡϣ%C� �� �[f��B]#>�Y��y̥���2�A�B_h6������m���J��6),����/<[\�п�$Mb��������� N�G�t�?�/�0i�������a5��hQ*=j��$�P�}�!Z�<TD֖#��W��a�.rwX�0!M�b;��'��S3Yg�a�Y&�*k�U0JҧE��֍�|5}�v�]x��RI� � �"��}�(wg�s�7ȫ���"�Ě<�?&���s�2ciӬQn��wԄ_=1��6��<'i��Eؽ_-�>Z]<��b�t�p�=��p�v�����R��R��D��OP̓��=?�,��on�����Ľ���������Z���>���u�k�|�N��"���?Ę!p܋��i��E���\yR�K�0X;�
HO�]�a+U�#(��4*:x�+�P��L"I.!��z��˿&~�k�}�K�B�����cH˗En� ����9���^������2,�A��>rJ���a�WA��I���$	x��'r��4gx��JS�����+�s����۩���}D�	�婘��36��˃�"[���q�xM��V~P���h����W�'w���j��WR�<N�M���0m)g��$����A�ZM���~�)�tA�a��6�7����p��~��2���_
�Qގ�LH�5�6/�`�h+&�
t�W���2h*J�2n��x~#��-m�������j��ma�����k��dK�VF�y�	$l�A˼u���x�=�(��K��v?���g�mgԱf�>h�W�	}�=/��f�q�_��.��2�f����f:#�r��������u�����#nv����{�[�ل ,����m�T���g�f����>k� �cZV�!��]��x��A|k�Y1]`Y�<4�I���-�r��p�XY�*���P��Pp�/��6y����ik��Pin��b�$|�ȉɴ�]՜2�5�"������d����lkC�ۚa���}#�����p�yq� ۼ�f���+�Az�h$����Dj<�����Q#,�9Qo���d_�\��A}�o���	&�q��h��$��ܙG���/�:�Y�r�'��[Oش�wFBLO�\K���č�~�/C���壵�Dp�1�U7v�w!ܤ;���i]�?�^�a���H�'J�9m�NCA��i�`�(	�40�x*���m/&����G�����l���X��@U'��,��<��!e��%�.�P3��)#p/�k�&6x�\��H��Ɉs�
�ni��<�y�G��:*�!g���+�+B��g��#�$o0W�?��97��O�4q��O��6�M��)�Ϋd%
]n�Q���!�����m�8�`jZ����uJf��A\��e��#4��;r�OM���_�h��w�Ƽ�[�9.�$$~��I��X뵥���3:\����u'54�D��\�.�L��4��t�<��G�ƙMx�U"��=��"ZAO�Y1���S|�S���Ӷ�K�Jy�3�%����c5�M�wF�
�t��f.wcW)j`@�Q�V����Nc�&FJ����ꖼ��˗�c���ͫx�P���_��o�f�s�`�6�+Ő��I�Vçtlϓ�(kE�?������
ػ��G4-����W8سL	c�Y�H�=!C�$�~'ŕ��u}����~LC�c��.զ1I�O�b�5E��T��(�p��d�������LW�|�< ��̕p��Qb�d��6X������y^�����:6]�o �M�ۋ�lyj�}�6���.��n��^�1���� [�*�6\�pd���*�z6Q/v���O�$���1��4���=s�d2W���~W�=ǳ/N�4�x'��\��4�jt#�u��k����Z0���t^�Ǿ�@���}6;�C`-�����]m��S=�#�
a�~k^m��}��J*�>ޖ�=+���ou�t���O�k!�j*I�PQ	���l�:����Y�5\�U`-��-t�A���৓������cۊ�ɪ��RL�.^���D�v�����_����*#�b4��/�%�x=k�±0tj��=�"E�s\-}Y$�-F0��$�!�o�1��a�d���,=5�uM��A$��eCw�����c�U�$���<3�	Z'<��怷��]5
<68>c�᪻M,lA���|�����Zny����BJ3\4��O6��J�[N^a)	��eo�B�4��?��h�#TYn�ݤ�!5I6�,/����z�J7��1yq|t�_�H�=XD I NF�m�U�X��ά����#�,'_��&�,�`$ELF-ݪe*�cYQ�]����I��ڂڬ��<5��/1�Pܻ�H ��wXՊIߎf*�T�}�~�V�	Ofx���u�ӻ��H@��3�px��^����B��`�6�_��f��gM�i�Pe�M�8ze��p��#^BE��)k1��;�KB�k��z��;�N�L@�ov��U�=��6��� !o7���4�h���|�F샜zƚvޝk�
����A�@��T�X������Ѱo�������J�tU	�D�q���6x''�RY��j������`�^��΍<�Ѧ���{���/ Y�?�O(K8�)0�~r()}L��i��e����c���f	Xi��G��%��Ğc�AuR��F���D�x7�L��P��ǫ����<�B������q���;歔=�*�`�r�,u>:n�馓�3��܋D
Y|t`�6C�\�gS�{�!�C�q�9�I�Oe���~ZiK%���J��`"��
�!��IF_uH�6���"L@��u��	��	�b�q�b��:��P�Dm�5d� ڌ�P.�c�$����E����2�5�چXJ���;��ǵ�l7��ѩ�
7�~|�'
�m�a��ܐA��2�´ނ�G�C�~1��2�q����!	 6�˪D�M/Y���G@�=�KC���X�+��V�f��5�ؗ��ҧ�`v�qJZ�
$U8�!+���'C	���&P�md7.\�/Xo37. i�ɨu�nV>�!�K��c�lB��u�%i�)��A�!O�����Ԗ�) ��	�ݢ)��'σwQL�"��Xi��t"*��N�eq�u�s��l�4~E�{㣀��  ӥA��|]����uF��q5�"��߶E�g�Dz�LB|��<���4֐o4"V�2��y�A��O����e��t+��}��yvr��l�_�����2޼R�7*R呙'@���33�Ih>�CԘ��mKO���Y�P�-�J���5��_C��_x�I�@ Yl���w/�Ba#?�C��ork]'��}x{r۪�!*	k4� 0�@�dD6�n�(�p荐�֗ш�/<�p�gM��g��nI{,#ܣN�<w�f�EP������T{{�# ��B�C٥�
1)-	���Ω�$->x��{��Wdr�����R�u����p��e`� ��&��Q�L���I��	T�뚖Q�/�'���3�F]	�<�o���`�	Z�#(���uʝLMw��' tۣ_�Ї�^d���J���/��<�P2�N3��]-X��ˈ�Ғ45�U��_J �0ȀL������ �xŁ�Ӭ���m$.�$�(�3^uO�˦!�,��L��k�K�s�t��!���E�g�(zp4��݆=TP]���lH�R��5�Co��+�t��h��{e_֏-���p�L���� %�>�� �I���]���۸��[�(�~�>�5F�윱.e_�G���"�5�*)��Q���_�g��
/���k��h��o�Fo{|��B��Ko}���(���36�$+��Lg�pw��H�P�bߧY8�齳��� ~��^��S<(��Ϻ�2��Ȃ�R!��Q�&�:�S<5��Z ��;`��C!�jms�{�7vG��#�YFS��zD�ùt6Uiv��M'�c����Q�,���ǍJT��BH��m9�h�y,����H��v/o��'�c�-a�$�p�jք���8�=c@I�f�ԫ�7ҥ^���J�[�X>&�[�FU�?�ؓ�(�k�}e���>ԕ�]��h���?\�)�y�CE�\?�V��p�.�|��gUӆ
����V�.;Xts��aE�Y�� Ju�/��a���P5c��]q�R0�7^��Q��(�>/�J�}�)�^�RL��mYy�{� �ʡ�|#
����0����i�1x��9;(�(>��ܿXۏ�
�%/3Fe}�����I�o{μ"�d��x���g$5G,�K�N�Cg��MZo�ˉ�N;&5�:�&�h���-��+B7�t��LT~�[C:`�d�� �=(��Y��%Li�_���Xo��.("�5�)�v↽l�5w����&T�!�#����Y�(�^�������@��O�[{���kiA[+b��U�X	'P�UA��xz�O�� ��[f~�Du�5)�p���?]��ۋ�뾫�f1�C.�g�/���6,�m�p:�``�a�r	��[����PҤ������Bx�oz՞���@�����^)r(�)�r#3��A鸗�/�)bN�>��
�������4�s�^���f[̤|^�3�7����g�)�L� ���G����nʹ-���H%�{q]�_�~F]�93}�pP*�\��Z�";[u�Q�!�a�8LNz�D$�Π�ȵi<Žn稔Ir��l�p��`��������b�I�{;�F@�#��|��Ͱ���6y��Jr�i��� NҘ���	�1�3�E�Ԧa������bs��'���f���*E����_�4��_����x��¢ax!n�k�y��1��`q���Q`�xv��:��k��J�ܡ�6
 �Irh� ��O�ǲ<�*B;Uf����)�4� ���2nX*��;
��Up�����_�Jt����������M^2tj�e�p��]�C�KB6@�v��_d�x)C��
.G�q�\�qRʡq�����#!Ǜ��R��ꔍwG�Ǧ��8��Y;�9�;���KV����A!ah���Y!��B���~��U��K���C�&T5w�ᔯc��w�Fszلa~Aߴ��D7��d������2�/}�J��i�#��DίY��a��$�F�ѐ\K'8ݓ�d�Π��U)��^�K �AK����Z��C˰&^�GLēX��+Wԅ<i�R1Tڎ�Ze�Vu� �;����Zj���uO���n��6ߖ{��d/3Z�+��&m��@rCFm\K�Y��j�e�,��v���l���g2���H��F�d�/I[�Ys2�t�lr�m����]?�U��1�"��!1�KPp�\�s�p�\|je�X��uW ��Ot��j'.ђ]d�gA�r��oblF��V��g[W2��GA�Ÿ��:�����'X)�/���@�,�+��/�[Lж�2yk*���ӵ:׫�o9�t�Z������LO>9��a�J(������D��$١� w?���l�w�����~~|y�E�;P��@���[fS�~��x6:����5�4��~�
��e嬵<j��8�O�#���WmA�3��B$P����Ŭ��س���ˤ�N	R��2z��*����)_#]tk����k��Ї �Γߏ��3D;�<���n�3����e!��X� j|��]X+H�� �lK�%�yO�w�3�r�u4璥u=Ŀ�H%��Z1��&+�j�H�ݚ�����D����:5L�EC�G-���V��2b�yq���a�4�E���p��e���-�E��zB�`��i�,~G V:��\g�2�1?�u����$sbL�rW���}`?מ*�����qwpm�E��p��lI=�dQi��B�;۷��Q�^3K�v"�+2|d~�i��2�*WX5�N	��9ǌiq-�}�H?2ɿ,4TdWu-���"��i�f���V�I�9��cE5h�^I�������q9u�==��ޖ�]�� ��V���x���}�� �o�y��XK�r\@摂Hƿ/E�ԦR�IFɾ�J/'��I��"w�FBR)�sR$����A�Md����aM�ƃ㭘���),�#i�Hעe�Ć|���T���c1θ*�ew�гU~zWF�j��@����2�ھ�d�}���g*3F%�]S�i��o���A�Kh"~����Ocq�������ON�c�Mpu��|#G0HM劃���'��6%��m�,����3��S<����g��ҋX�|�����4�W/�ժz*M�ٷ�R��V�#�F�!+��9�����Ϸ�߂�� 0�Y=���sOԿ?���u_��|��~��=�Q"��ڂ�xPd�]�t�&��Oҍ�]�a�a���B���Y��_ns�F��c����aL�-� �Y���hS������A;����8�J0��d<��,�!�Di��5�Hl��yts��4v�Ig:D�*gƓ��V�4F޷��9;Y�����k��a�!�|���*��K:7E�bOH
C�`s�u{�NI�h�������N�5��C�bzs�e��y�h}t����r������<�N�}�R5m�:�Y�na�P��J��t:��h�ʃ��y���h��m@RV��Ysy�J���Hy���8�=��y�Mn�F��K�����wc�a���E�Y!h�-**!j*�Wbk!�HI�w�#}6ʓ�]��%�8_z\j��W΅�E�/d����ãr���IAD�_�|u���؍�7gO蚃n�ߵ��i�0c�L�i�$��bR�2P�d�C��}鴥�b�v<�j�n�IM$��(�useUX�SuY����k�O�����5�x�Ǜ�i��YE B�� kR��*}&�

���uIYEAI�-���V��5Y{^f1��������j��Xڈ�lvA��WeU}q��l�O�|���bn�\����i��	L ���-<����uN���d�Mӕ-I�	�kp}!�M-(?.t�(�1�Dz������<pD���< fE��K�@k����?��6L)�}������-�V����h4ϧA�ןf�7��c�IHO��� �pgbȡK�x2c͠_*%��G�w�k��.UdZ�G�}�J?�E��m��|h{�(��/,ux/�V��(��Ǯ�e�Q�D�1���0 E�Z�e��(��s�.�<-�foI�|��_>�������x�#����PS���s%���7`�İ�P�g0�g�/�p��}���K�i4�t����$-(��}q|(*���JO47c����:�Ǜ�����*7��#+�����Y�+Bfv�9t8�[��0c�t�U����-QN컃�|{�"����u/?�_W��d��
���0��dѐ�ҽ��<.�T�NQx����BBC��\�a{�L~g�DVF7<$�,8��;BNm��WV�\p�d���"��03J��@<�!���n�UK�8#Z�]����C$�,D�4�td�U�姤�o�^�Q��,~B�ԪH:��為��5��/���]��:!Z%��� ���Z+b����*�D�">&�GЮ'4��u��T�)hU���NJj5�@f>L4�PQ�����r7�r��t�| ���+�t%)W���ܳ�-�#�9ڣd���g�H��w�K|%�l:&��B��j�4\���2�"h碦��!8,6���_\����XR��O{OJ�o��V��,,�xޞjw��d�]?��emAQZ�;�"���n	6+?l������dmh�����������mh���pyTo'���6Ԥӡ�U��	�������c:��u�D|�����q�9������&4����I������?�����H������G�)�A��H�����!.ތ��EH#"?�DeEy�����~ �^悄*2J�Si�Z��g���kc�����N��*�?i�g� ���� ��2�[�aY��r�k�U��H�L�3�������ߧݖ�~�M>y3Q�����[%[pLw�(�0µ]�)N��k�O��@�X��B��SW��bk�_fy��!�j��K:JBKT�F�Tv4��}��TT�]~��S��J|�9���/��a�2O���
Uih�7����H�$y#��'�Y�η%[��&]���_��} x9DR�'1nk��<� ��K���xr�/�!�'d%:��Y9�B��� Y���&�}#D�����|����t7�
��������e������o�mq�Ȋ|�5$��O��&� �d�7>Q�{.�C��R����g���{�b�ְ8w�;��+��;��HN�[�� �V�Z��D�J�=[F@��K�{���}x������Ċ���)�1�_4�x�2�� �y�l=�`Dw��R� <kP��ƹN$N{�'fLS�Qʥ��M;����4��h��C>�9{$h2`�܁E���]$84�Q!�ލ�vD�'��`1�$^p��\��>�(�|���3���p;ԇ#�+�g��'w$/}�&��^�1<�t{���j��2@��Af6'����`�t���\^>CHm>�;��l+�����.a3-��S
C��#�u��BfG��ZY-	�����a��+��e?n����������ٌ~����:�z��#�l�o@}c���ٛ.᜽��B�}����勥�F�3�C��YY"w5���]��"��xnx�������� k�ƀ�B���m�x�T��E�Y"Ҵ�l��\�`��ѣ&�K�~�;�9����.�o�h=�ުjv'��o�qt]��&�z�	mt� �����`A�
�~�F6�q���+�,�I��ݪ�Me�~a����l< R���5:Y2�u��]��
�<(#^eR-�H�r���V���%��l�Բ��h@Wе�'��ͩ\r�N��Ɗ�iN0�)���Ɗ1�Wݛ��9�t���
�<$�,�6����䯰�x����ۨ�סx���]h�}�	��EV1eG��%�$6��C�ud/h��䣏}w<^m�t�p��yo�H:�Vx��~Y�����6�����>�J;e�'����Qa�`^����=�,�5CR&��қ@ʼb��Ӓ���Ly���=(r�Fvr�Ϻ�=�S�MGV��ӗ`q�
]J����Mg��ݎ�On���8��3���M��a����cy`@jG��$��?�E�)DB~�S������?�_����h�Y���8q��I�T|�sg�-��pݪz�hN4Y��O"���S�F��T�u��j�eyP���9��ͼ���Wį�)p!�!'�ˍ���B��1�R���V��^FV��;�?N=5J�U6��Q�&X�,=��;x�n��
A�����a�9�U��4�y���W�uڥpO»��:7��슗�6�Ċ+�5����[v��!&z������"`|���6z
�P�4♖�M�h,���6O-���dl���	�E�b�N>Ӵ),cs�dD�a�r�F1�m?�C�Z4����$�TO���7ܟG�0�Sh[�t�2��-5�0�ޜw�x�&x��莶۞q��3w|厡Y+z��;�⑉6��\#H�Q0_�2���@!ڏG���-�Vv�E̒��0"�ۃ*�N\᪜GYRe���"������
SnL?�1�q��O�TvV�]8�+S29+�A�DT"	�p���0*��ip�I+�H�����
tqɥ��(�qS��51���o�_���]���VҤ7�H�&��٢�p��'�}�%{�|�:Ij��K�,5.�{��\U���=����q� �����Ac% �H�(�	Eq&�vUv���^�'�6�<����Az��Y?a,&D�޿KY�xV�T��&s(�ŷ���cs�0&��Y�-����|�MҪ��Bqs�4?\�$]9����8�g��频y�N��B@N�pm\�u��ݷ��]0�5rV_��.�\]��H���'�a�,�/�a��������df�q���X��(���g'�dō0��.�j�p���
=-	�j���x�CmΩ�2�χk|�d��[�d����޷��!�P85pAg��0��k���v@V�%쏬�p�V������tw�ƿ�)o����a��sVV�T���l��/H�fR�
1>�Ė��*�e�Ӧ֫L������u`8�g���9ua���w����a�Xz%w���!�V�j g.9���uSa/�h����	|�	��Бm�����8oj�x��H�ϞJ�;����W�YmR!��!��s���k��%Kce(�~�UdX*�L��I��2���!��D��W�bPz�T0��������$ȕޠ����N�ӆv�%:�`u�����J�]wF�` ��"SK��)�`��d[��M���mẉL�gbB?����Ub�c�M�Qp�KkCVi�����}���g�Y���y���<����1smG'��ͅ�}�#�{��!PC7���iagO�ZDo5��<Li��D`s�����8m���="3�v68�/��J��e�(�U,��e�tB�e)ċ5�r���N�.��.��8�e*PZ��(aMȜD��R��ú���Z)����[!E���n@�g:�j��4��o�����i�3|
�*�(R��@A�7�2rT�[�*D��oXk�(x�i�:r�L;��7�ڦ�U��u~������Vy�R�2i"f�ݜ�6��I�K��:����6)�U ���=�E��ɩv�\��k�d��X(2�_dq,u|���K;�Eذ�������h+��.�<�n��)���i�VD��:�)|��+�P!t$�Z��;�Tq���Ƿ��V���8i��,/�so}���~�l�K��ԽcM�i�?q�Ps̺��6?a�ʶ(��$����Bb�i"���9��f)0�Hp���V�'3GS�%?�i��^u-��1��dY�B8a��n̕ܝ(���YXb�$Ⴚ~ �'�j���ɲ6�T����é���\���X~�;d�-t@渋�<Q�'��X��xD51���1�o�Ԙc���I�G�Vg2	����u�m�ܥ7�\�Jom�ͿZva$�?�F^T�[�����L��#�	gnǙ9_�U�E�;PiI%P"�%�dY���{��V��1��
Υꏚ�Ƌ��*T:�PİK�t��ӑ�o�=� wG��#8p���^��|f�=5�kS�q>����|����6�>��Q<@䮧	� ��m�"��F����90#����/�:�?E��[(�͚���Z�-X�j�A�Ka��~՜7Ļ��z(��B �p�nG��Ks�1*6��>oy
�e��V`@���B�>��I��N�3�iv0Ga����(K��o]8t�U"ϧ�-�.�.�R�uBk�)���w;^�М��(�4�Cj1�_$��9�q]_Z�o�xvv�%>�>�MG�Q:rD\4,�i�rB��-zfDH=`u�;O|dw����(�ZUz@o=L�!c����}u�TQ��X�j���
yɱ/ehSE@%���j����@��qٶ��GA!�h���c�d����>���@L���{Wi���E������:9��QH�t�-Q�Pϼ3�-�d��Eɐ��A3�6򚚷|w�'���0�F;�N)�Ї%��|O n �>oHD 6Yb2Rk�U��/R ��s�I�'��[8TV�&nxb����R$E�1/�����G��Đ�w�ഩ�*N���p7Q��.������܋)B
̑a[���j���l}���R\�7�E0�0���k&�/�W�^�sU�85���6��ӈA4=/(W���-��C-SU��.n�^f���@9�殊kN��14���s��ϴE�hڬ*t�[eLs��|���o@�j��hz���Q��eG����d�}fȅ�B�|e��~&��
r�~�mh��	=�&ԍ�A� ���$;Zh�ܲ���BXt�Y�(e8��S�c���㈩Q`ҷhM�}�6����m1��0I'���'�'+*�}�&3���il��^޳�K�V��\�g�paN�m��^���L[�ļ�q��xo�{T�
�;^B�/���_y)A�0�CP�T��z�2y�g���}��7�8���8m�V�{w���>�p
��/���5�9��%�cٯ
�?2� f�,����F�{`Ż����T5x��b3�ߧ�=�\"p�<�Uғ8�x;*j �p���{|*HI�o�O���ōG�>�@N��R&{K�|<|�.�c�הu�`�������B�3@���ʪU�!64�S��]u���L���T���tT��aW��U���8�ɔjrG%�7{� ćvtr�}�|�I�!�yS���M�t&���4�	嬱oWPIl���/8�"�s��0M��`~K�a�]s=E����߬l~]���K�I�A@�4#bĜ�`�ƃC}B��/W�(�Zp3>L2bI�r�V z��5\4F3��{��9����{�v��^HY��oU:J�.��2�wS��D|H�_��9�O�7����L0K�k��l>䥒�6�P.�Yq�d�����<~�"?6�H]6���n�؀E���~�� �?ױ[�}�Ad04��J��P��,F��]:�h~E#!�a$������]?��Y�k��?i�� �,ɾ�� ,l=(N
�b��J)�i��S7ЫtП^�$BK4�m�W�?2T��4[-|�4�S��|0.���*�Q?I1�d�Сje�G��5���R"�l��"��,���N�B@oվ{���w�����y��;�*ǛT����-p�$߇�Fu&�o�'�A� �o���dOm�ߜ�-�����y/\R_�I�s���	�����`^�:B9�3���>� 9���ް0H��p��tМ��U����|m���kq�?	V�鏰uSLT�`?�2 ��wY�#�Y�-�Sq%^]Gu��8f��PN ��@��m|����3��R)O;˙]᥻$T�m��\�n#�`0$9��*e��\@D�VS|
�pL�8W.&_1M�~ke�/M E͙F(���l�Bb�i!�ߦU�ީ*Z�ұ�ڃ�	|�J �T�9��-E٪�/M��{~`�%�Kɩj�=QS�鷖M�l~������lf�1�V�g{�K��o'��	�6l��n �a����!��;|x$G�0iJY���s�z��bU�oїM���u����+��.ı�C
W���|u�L�������\�T�L�s1���{_��*ز�~��c�4 D�[���)��G/�����>���
:D�M^\�AH:j}dtH�V^k:��)Z[���U����
�Rw�j�f�Jk	�1ڞ��f��V.wr���qz�*�^y�����Q�VY2EK��5�2^�{�Y���a��Aq�$]v.���)k�I������[B�ŷ~'-�����\�u���4"�X	�[@�N뛧{���=�d�ᢝ(�?�Bg��wW+{��:mLCK5���e�Z���N ٍ`��Eݧu��H!-�Y���q���W��h�+*a�8X`�Se"���j����l	�\��#P�'��0懤���a��Y��b|e�a��i��K]���pls�1��j��S׳�\�~�7H"XN�2��{~Q��U��"�9f<��vN����#�B���Eyfu��i�I~&%��w��a�4(�y�}f$m�P���.w^�^ڪ����Q}:��A�U���:�c��x���2f�.6����C �5�:�bL�s�30� �zن�,th��r�k�o�x�g���q�� �d�L�A��vd�_�Hr� �E� ��T]�	 ��XY̴&rů>Uο�q~JB�oZZ��2��.U�G5�%�ۋ���3f�ؔ`�$����'�Dd�M����. ��]�ߋ��;��~/i���؋h�xd�Pqb<m�������ܠ}��";�2}�@��(�3VP-��Zk~L��f�#O����W�$22�Lڡ}�r����u�����lt�y���]}� �ֲ�(��̷�w���9X���!��M��,g; J���v��]o~lCZY-JpD�����I5%��%Q׶��e�a�<G�� �ݷ_ `�g�d���S�P��%�rѳ#�:5^���eB��X�,;����X"��@{���V.Lb�ʜS���nW��dHyAM`5�.��'!���r�M q�'Ȗl�QEǔ63��.3<ߢN�.Y�Bj~�7�(�y�S=	�s*�%��=U�ՀK������
�=�sڮ�K�խ_3���i%�P�����gk�{�۩(�~�+�#�|@�D^��>�mJ�+��1}�����P(��\���/���ny�NbI;��4��<����ڬE�9׀��3��\�`G5�{#E�|\�6@D��|�60�3��o��zI�y�5�l8n�63EkKqs�H��ĝ�D�>����VoH0M�;�*D�9NF�^%�㋵ޝ�����@B������'
����ãV-�7x�F#��F��D�h_��4�ڱ�I.z
z	��PI.���R;�A��)��!� ������YM$*_�
�x��J�0��h�v�4�	�15<������d���}���RQ�=Ԋ,ykQw�e8M}�zu�WE�ߏ-Bd�� ?�jv���%P�Wt��Q�M��V��@���>��M�3�w�U`.t�l=6F�W7�Q���N�O!��.kɻ��h�b��!]��Jj�>�$X^Uqz�H�ද/u�o�����N*f�Q�˼��>���sS�7�l s����Du��P�×�S!��0���������\g�7���rGt���9(�i�ת�`�5�dK��!�ܽ[�X��9q�6�,�kAX3�M��E��*�����2n�����s&�(_�'��MIB!d��|���3��i��#^��y˫̖L���oX����ͫ�h��?��. �ww�Z�?��ae��+�2�S�}ߥ��$�si��J"����� N+�ƚ�������ї�'�T�nw��:#�����I'Sft鹰��/#��\s塵��)�DQ����CY��z^�� ���Z�w�0�|��I~�P��)�=@M��*� V����ڪO��qzʼ[p+���|�!��+��h/�S��@�N'K/!�x��@��9��T���n!��r
C��̙߃�����?��5���e�h�$��Q��E@3�䊥G�0ֶ���׭�#�Ogwq��C���<?�4�E�ļ���9�X����)H��e5^�Q���pouɐ8h�Q40���4��W��-�(}7RJѤT��y�o �A��<����Q���Eч��m�&82�}�~hK�o�DBcU�H���W��*��D;4z�Y��Z����F�\��o������{�*��5�cg�{������e�{�i������ö{����\��/���f@��Ϻ���f��%U�*Z�HY�D(�|��.R#�Z���9���tY��vZ(k�6�&	���V	].]��^�g<�6�b��l+Ec�7T��q��(��Q�N��6�$��ݫ�9m�R��)��UJ��
�e�t��U'�S�F��ִ:NB���*�&6���{gLJU�?��Y������o��C1����R+��\��3{�]������C����ֿعQZ��lH±�O���(���'?�Y'����/�RyF���L4�PT��1�OR���Vt�.c4�f|�S�^�7��qz����'�آ�)��@��5ǔ�����Xշ���A���F�F)��U��;;7k��X=^_кU�F�EϦ�S������ri�3Y��\�x�������t�u��$�o���<ucVu�3�0��#/_6k�ɘ�n��RhkPN��`�v1���#*��{�7�Bh��O84�`�V��p}vFv�Z+x�*C�8���ʻ���kuL�jP�c|�o/;��Ϸ��uZ��A)�@ �f�8��ɵ���\-nj�}�jkQd��*ɗ���,HZ�q��1�q�a���9O �gR=4�6j�x��Q�.H^�-�`z�r�G�f��|��हH�Kbw��Q߂�d�Xo4�BC>�{i����6iv�$y=2"Qĸh#L���G��%V�J����,�R�a�AZ�.�ڦ�ř�< ��yr_�t��h����{P�Ht�e[�v���$������n�%��ˮ �_;��o�?Xo�_14��EΠollf�$�_c���k[*<���<dLB��t獻�EV��ѐ��a�p�z�t���bn��̦�\W��aɜF̫=d0B�i�.�:��n��p����St����f��<+c�OT��	k����`���؟�.�!ZeB���u�f)8��όH�`ݙ��i�a�o�J���O��OΝ���Ť$pg�3�R�MID���}���[݄yWm%1���"�=ǳ��~%(̶=���z�9m2����ns�D����4v�(�Y�� �A1�pMϛه��7�^����-%l��;��s��lɮ�B�����������j���6G�`��߈�%C�^��I�1��c��E�O&l]�VXR�7��Ɓ�os��0��\�����wd3@jJP E�H2�)�kٍ՝;��<��p8I={�k���F�/�y�iL�_<`b*P��R�)�ԌtP�Y��鞶E��>6J�t�r{3'g�?�������aF��h�x�#{�j6\W���+�{E12����m�C�VGh�������|�(Ok��/�$]�4���H�Gٰ�(k�պw��c���N��O�]�9�u�6E�؀��x��nhm�
M���ƒ���9�6i�����}����ƃa��B�( ��SxJX�M���b����ʖ�y
ame����w��>D��A=N�]�!.c��#�P�-1���g��^�ŷ�h���d�9��s��.�7.j��JY#9��R��5O��^40+�#�|��X۹���s�.Mr�_�R�]\��(��Fb�'��\o^S���b�M�i��C��&ms���ʑ㭳��c�� ��.�E���_��&X�9�]�v�|��е�b�XVB��3�*d۬ad�(_VH��dgan
�N$�t&�%3��� �u���$ᱟH`��M��5��
#����z�8�s��{���e4���;�D�C��w*np�T�U�cXļ&`]c���_�5���~d�Jp{�"}��.�q���I���Ѐ��v-(���<��Ļh ��Z��ҥb����V�Qqx۲�SFt%�d^����7��XJ�ab�`4Θ\`�J�A�B_jjC���I�� �c��tCt�T��g�	﷽Z^�R�J�k� ��_#Q1fW��0����(8��X�.�$H��n���z%y0Ԗ��0��֭%��U�&���fv�rM��,���bd4C��ouʇ��lq�w���Je(0y��� �ScD��D�vYO��	cU�F�#ԝ�����Crȷ�$(!����¡��pR�k�.��<�h�ql�Tvt�X�\�[�Uڧkl������r��a%��;֥OB�<0���Kք�C�M�%�ۀ�h�W�cc,��hHAy�;����#��|�����ԩbg(h=ӭӐ�4��/�{F�6��J@��v9��vxk{F!��+i�k�7h����Or$�u����q��2�8y�>
<��~~K����]d�X��M˙�a�0hM9�'�W7�.t�ueq��6>���,�[C,s1��\�gP�%!4�M�������m�Y�D��?hW��=�eMCW�d�b�u�n�gś�2ˀ��І�zx�q���#���U��Y�C�E�����v3��X�eLF��}y��ZA\+z=#ǭU6D̶ef�OԺ�n�nFڲ((�?��b��t`s��Z�FP­�%�{k��}^XL';���� Qwd�s��j� �J�4���M�oH�+=��JC��T�u���E'6',>��<b^[YTn�"��a�ȮO'Jb�,�Qr�h5fr�3�4f���Uڗ֍���=��)���~}����s��?ٓ�]�CG�� koů�"#=��e����H�'N?lC�D~����2���1���D�T_���a��|�l���$�9�$���/ W�k��2?�g!NO#a�\!������"��8������F�[��ܙ"���;:}i���n'�JJIx�<��=���ϛ��q[K ���Lh�%1Q�\�����|.�nm�����0v0���Z�
.����fv�!���0F���t�:�uLf����܎��M�ĥxy�u\n�ZQ	�9�f�����*��\T�Y���	t����	��FVY���o5]QS^W�������}���,�y��5�#o�t1�$�xF�����9"�	����r���cET�P���H�^Io�ԁ�.{lC@��o&e�~#v/V����A�=fCU���+m��F����_��n����m,ѶY�Q��[ŝ����ֲk��2�?��+����,W�Tf*��jSh*�8���/8%8��$kr+�:Z��[ Y�~�+�aOQ��"�7�ø\��ǻ��e
�^����~�L��U��[&w���q�i*-)9Q���=����"
��a��)F(�M��2F&��l,W!}⳶�s	��ѫ��R��=1�9Ć�,v��"I_�RH�����34�<O�Y�v�?�z��͓��P��!}�`F�ڼN�����>��}1��{X��w�#�� ��D\ ��YUs��A��C���T}�.�������^*�3���|�m U�e��Oe��N+�QED���6��E*u.Y���Z+���= d�ZW��c�b�+h�d^&	]ZQb�-:���7oϹ!�|�?�>:��͙�e���:竦�A$��5���?�y��X��C�#���V  nq��v��D�3(⋟8;<^�
a� G`��d�_lf:���a�~	�WeP�����t(��h�T��s:�`6Z�ҔD�S7-mձ�aK��d���
#�G�2�����LN��A$u���+�������V��
H�g2JՎ���6�����<N��! 	t���_Fͽ�L;�؆�O�%��%+���6@3�[̀�c㸏�Of��H$c;�Q<D�G�C�U�dC��Z��b����X�z�D�G�!��u�檁be���Q�s\��C�l�5�6�)x��rQ/���e��F��:<�S���� �ׁ\�VeK /��͖�8�W����+��䮍-�_ �g�:��@�����doz�����P˛�,ڮq�3M��ven/]*5fʹĵsaEj��zD�o��a1��}��^TC�̲A/�9��Q)��0��=	�3B��u\FEYm�be'�S�bsA�.5�
�� 0���i�&�B(�BND�>tÒ��� ��huX�Ӱ��@TY巿6�8e��w��h��K�>�ڿ�\U��G���1X���1>�($IV�A�oKP���W;�f&QvI�c�����V�7���f���*H�����U��-$!UU��F�
�ϼz�Y5dD���E��X5-:�x6I����<r?Ɖ��n Kfᢦ��!w`v�H�Lv �c��^�3���d]nξ_�ku2��d��f��0�vE�A�z-Dbٿ�G�W�V�G��i0HV#2?]U8/�����
q���4 V�4t(����e�Ld�Q��A`b2z���L����ve��{�uu����}�Z.�����p�N!���\ ��b�}������?N�[b"�]��<����0D��P8�/G��`(��4���
�kj&��daA�K�\�=O7x �8(U?L<������_��z��1Y��h���)�9l�	���Gxu����J��y+ף y������wzH*ѓF�U�i
1��ǡ�E�1{��%�C�T^��z�@_��K鴞�����^q��#怂�r�@^1���������,�&v1�j�v�Goa-��1�>����jq{>f����H0֘��J���b����kU��B�����ݕh=�Rd���`�}):$N/��дqF����&p�F�t���:�O��|l��C�g��U٭aZt�z���I���{aC�T��L�-KK @�@p	�gdĊ�@̆�7o�V����L�,�ي{�N�"[�[9��@��)�l�r�6��V�Ӆ�ZNX$>5�&=��u�4q�E���vO�m!}X��ny,;|�r�`��no>�� V�r�GT��*�=	�P���7�V�d�
���n=��7h�N��dwkb0�b�:=��`DRP�y`N��u*�~���N�n���5m&���R���՚��B��0�O���6���7�;�����"�]��C��2����R,�_$�ID�����]��I�=��	�W��r"c�l�Mۮ_���ܷ��>nz����l̷���.?��������?욹]�xBT���n�������t%�@[����n⾪����"��"Ԩ8���һBqA����;���g��Ġ�;�. 5Q˿i�����/����pZ-�%}+��3�&_����	����)��G�73�<�` �WU�F�̶R�<CϴSc)qs�\�&��&�5��/�I��H�뷧v����P���\��d!ةf�F�D�u����Ƣ��+�vH!���r��ӹhe��Si�a��".9҉���^D�d:g�d�dei;wcu�9�YeV���wx���U�|&H�"76-��)! �*��>$�L(�K�j��r�̢ڏ���84�1�p�10S�P����������,[�ݐ��v��&��O�8���'��TUD�h���t[�[7k�grfo���`n�����c=U��az�t����OJ ��"<���S�!�K�4k"+������Oe����r 4:��ȩ�	+����G���hp�͋�wO�SM�Q��-d��6��V��Waz�=����C,:�`s��ț�r:�?�+��m9]Zӏ�Ct#�9�Wg�#S�р�U"p����[�Tu�(��y�>@8�/d�I[���\9Oޗ��4w����.����!W���-�6�����ˇ�Tm�W��Kq�i����4S{�8��ļ-��$n�o��j	��U��K�+G��tl��:!�� �@����&B4���:Z�rc\�
z���Ԣl�g��4�N�o�,��-YɰҺ�h����A�5d���;��7�XyQd��v���&v���h��Cr��	����an�ɸ����+mʩ��S.qKt�_�J�l'��iд_~p��Yv��F}��ڻ�R�|C�óڭ�E*|?��Ɓ��D����7L`���A���'f#]&���ؽ��g�"�x�ay�Z P����ؼ��x�t����r$l~��!��|�_h�veD|.�ᳱ��)`��"T��3�^</*�ed��󑚯�u4�6K耎!�)�͹<�:��z_@PF�����*�AɃ��W�-Yg��]��!����}�f��[��f5�N���{������_J}�Q�P�4�7�C��0F�@*/��)x��g�wja�𭵉?���gG�ؗvc�;?�QYQ�F����n`�@��|cĂeX�Xk	�B���r���0Q�H��\l[��Gٹ��o�A�^��na�("��w�wO斀��<L���.9y�6����{zE%ɀ���*P����-�6��)c�����6J6~���M!P{}�s�
�N�d����ͻ�nz�z�����wjB��d�ݾ��{sx�ܝ�(h=�&fS��1��3�N��k5���fQ����oD�2���Q�,h����R��3 ���\�� �FPiiI��}ʽ�P��A�p������]!�|@�4�<,�\�@�p��]i�C�sƈ�uB�����p-�OL�����B���xd������ց@	��=��Cg�)��_)�؝.��"�!�,��o��G:2�U�ch�ۭ�-	�s 6ƨb�{��8��n��o������*�����|N�d�=�����hJ0��D"5D:����w�.��{��xru�
�}��铧X�媰t����f(�e�����2B����/+��E�B뽚>o%"���ˌKb�h�Eұ|f��� +���&Ώ�?�c�Tb�|�V��ZE�%�Y�4	�xK��K�p�s���_�,m�@��\�^xj���I��wtX>�P��)2̨R�������w�����vU�!��☳����F��0Bk%]E@���dj������Dӷ�:�9"�Q�ꃐ��Q���'p��cv���J��<%nU(���qL"Һ���	U����<�� �p��XLd6{m����V���+ZdO�����0�债�H�KN4���눪%�����=0�7YZ�Am#B�2��]6��H�e@��@�10�a]��:hH����LO��y�jM!G�ͨ킴��,$LM��K�[�j�/�X�ZG�	�uq�¬`�'s'�w��R�p��sq������Q�d&@�%0&IUAq��	<o��O�𝧨��v+=2�{q����Hk4������2I���,��/y��;/����������d� y˵MA�cұbG��E����o3˶�QI
����;�?��Հ��\��Ű���i\�o�O��䪸���DJY��\�:w��=��9���D��j0���
��n+b(	ev���U�Js���p�g����� u9by ��IO+%i�>�g�Fds�L�"��&3x_���ϓ���H��;���u�Y���ϩB��u�W������8;�vsN�Y�~��ML��H{�*<��>��e
-!�p;�:a��W�v�=xc��ա�Z����#��H#M2��qK�K�:�XՇ��H\tQ�����/�[(07Yv'��ȵ�"�2*ڣt%�F�r(̽,�Hz%o�3p�Օ2���:��/��=3���kՄ��l,AB����7ˌ���;B�[R0�=x��b��&��+4(~a%�`�yqk:����Ӵv����4R�{�۩�&�^����'������ы��\���3J���A/�L��Σ�*u�b�vWV�#�n�Ra?O~���b=�� �_h�9ެ%�[�ؗ����?S������ww5Yg�&{:��/�}�Oy� e����+/��o�uV�X��8��.�or�9	���p��<Q�'ݠ�.�.�0HJ+_L�9`���Km��Wܧ��E/�=y�����2�"@˪D�Fj*��hGlyV���ޱ��_���7ପ��Z����AN����ޠ�jY]�g���	i���� ld;��{�g)�*ei٩���cCK���2�i�X/���ӹΥr�������YY�ǩ�tT���,h���r-�DXh*4y5
��}E��T����6�0���tk7�ӓ�o�x���Y���`RQ63G���V.�AޙH}�-��ǫ��
cJ!���	|B�jwtǬI�M�SiU��?�E>�n�	������H���-z$���d��5-q�Yc&4�̭O�Ri�mXm|=����
������z��Z�8�M��J�<��R�a���7\�[��6�ܔr�AT�: �P�)���:���p#fX �ս��w2�����d�=}9s踄Ԝ
g3��w��|�
׏��h[�=��L�R[a��-�P��,~��29)h?�M��N�O*R�B�n�����I ���u��F.9� ��>����D�UI����#�,�TH ņ�r��{�\jOc&�y�#�|�Bbã{�t�r%������Oj�zkn.F�2��%�⠬��?�q}ʁ_^�l�W.V��OR�a/�Е��`N������"x�Is;�&5�?f�;/X�:R�@�
F�$X��O@Zú|<���φTJ��)C���d�b[�	_*I8còC�AB�<�������5Ԕ�R��\y8xeo�� @p:��*
�y�Gt�(��5D����:��Ɗh�����5������_3O��{t��́������(��X�>��+���(:ϳ�OJ3�3&�+���4�K	���^u�����U�P��_U��7��j��a���{����ʙ�1��[�nk\���p�Ii��tr�q�~�)9���~�w���c|
_���|u�r8#	�0�bqF5P�5i�x��^Z��$>x�E-�Y�: ק��k�1e�Q
�P`�Ą[�~�\��G9o��[my�=g�4��If��*��#���{m_jBk*���{� ���d�7�s��܌-�����˞�K_f�0*�e`�������~�c뷌ĵ`g���@* �
�Ӿ�<������$��l�P3��(��u���9H�Ғ��X#�����-7�*9��/AAU7�p�&�����h�r`t(�$����Sc�K����vGh��drh��O� �Y��|�?n��"�j��;X�4 *��B�CH�9��T����R�óD���E�'_�����@(�|9K�h =��[���T�T���#@����Wq���Tr_6��+�oMi��'ϕ�\eqV8�� ������aCI�N�𖱄1���`g���0G1�1�9�	ă8�qlb7B��P�]0������l֏��%Wĵ�O�u*>�C�}�$<HNH[�������59��R>�᭮�ʪROI��*�J��S�U��ӵ�x
3bީx��W�����(��?��4�|�����������G��hW�2OZ;���������֥<�3�d+�!1��
��sw��g�8S��Zi\v�z9�l4X���}��I���*"G�p"1��:3md�e3��!vWu��M�- ��u1_���&v��i�<e96��(QᶱF�۟���WRt�A�]������Zh�j��M�P��n�v��tӔY��ӱk1�Ծ�
�7��r�{�qƃT�Q�^�G��I���e$�7��W�3 o~��sk�������ۍe�@ؓ�R�.��@±	ydOZ���R�'�6�Q$��y�dL��-ԐX,&��?6��FH�,�^�[���/��-��7��Sˮn��0?�
ᇅwY���SI9�����Jb)����l8�h#�J�&F�?�Q>s�b��gᯜY��KG�Lp�s�S�^�<������i]� .Ow�j��>.�^Ð���=��Y��|�iU�E�9�Xd����	Z��x�a�g.L��ƴ_�;`��N=7c�:0P�@�����o���"]yiI��^���#�۝��[�T�uw�?���ڄжl�ư�Ꮊ�?'I���עr�r��F= �sg�8���\d�hw�FD�V�<���s�C�V>S����s�9|3�5J^�?zS��@wI!��ξŸ�?����*�,,�L�5��h�����F��K�q���Ff��O��b�M�^.�Sh�թ'��ZkW	dA�>׺P�a`TdT��`V�y�m�_Ϩ$��x�_�lA����K�Ï�s�e5!�87sK��! Mb�`Sc�������\x0+ߩ�)� T0Y��#����f��/o{�[!ݶ	�AhXDX�ܨoV�Q����2�N�P19z\#�i���)ї����
���|�rZ�ј�����\\`R���Y�H�O^��V£M����]��*��{�qr�^�	�|w�b�L�<�����<:��'1��ڢ./���8�/�:�cI́�����/F�ni�-1eS�/��w1[8%�f�~[��ឱ'�������lb�k���4���v�u�*�{jOd(c��*��=a(��ӣ�+�a��3�����(��LM�%�ACT"�e Yu7�]B��/���
�y����NJI��T��������xG�(&Ώ���&��/�$T�P���k��)�&N�?�P�+� ��/?�c�.�:+2�?���Y��s~G��v�\�B�0o8���s|t�S]!�ށ��N�M�'ͩ���trtFVC���d�����H�\�-vU�7�XsxG ��̫�Z����mMK_�;�
�٭D�?�Ot_�<|��{
��e��<0������=����tv�s��X!t��av�(C���mt��h����n�Y��d���Gū��p�`q� ��I6-H�P�+ٮ�<zs7U��:�x}��f eM���"�C	��9 �u8Մ��&����v�������L��ҷ�������>i�(�t�]��J���1iB`!�X��;�^������Θ�mB�~�C��W9b'ԅ������&�4�b��{X�D	����F���.X:�R����E^�Ӕt�ղ.u�|��S���⧊z�.�ּ�ۡ��r�0w߬�������ÎiD�Rc��7��^�'�$�5��ێ�a���)<�:�8��c�B�d$�6�er�Yk��X4�g��]���"�d��=�s
<�0�E�m�w���(�q�2H��R$�jr��st������،�&Q�bDx@]%z��*-z�\�Jvp)���\%+�<G�a�q���P���b��������zD�������*�*/�����#�VUZ%�=�u�S5�YF0K:�\�{�GO�+	J�V�4���~į�J3���b�p��mC$�l�[���F_�^�JХgf���;��N'O��	���scR.{�� ]M�p*{���X_MA�!z	f���f�/��i�oC�֓�0#-�F5F7�5��]J��n:�I����]Đj�}�T��U����E$�V��W��r�`�U��*��2��i=կi�}�R��G��*�L!��@���=���T��C։�h�b+n�#gT�`� {���ET���\a=�h��o�NW��&���"d�4�),Dy��M���|��/�a|<����(*7��!�g�m��q�����#����3����U��%jNN윀�� �L��r��഑h\��jû#�?6$-��:�1�L����}
�kz�s-�~G;��A�2���w��S!J[1dh+��cې&L`�8y׷�dR1�J	�R;gae�P��=m�L����ZӦ2��0V��ă���I���2��_ݦݵY{�t�,��{�Q1��V+�;{X��Ϋ���i� ���̤_B��6�F%T�ھ\��E��[���@p��'��hM�dB����%�����=�@o�����:�b;�xER�����Fh�6�e�T! '�om_'�R`*z����mW1����������`����{�)�+v}OV�"b�n� W�=��P�z����_(k�_��J|M�ŕk��d�oo�p:0�&�S����c�vp��Z�>��0���J"3������O��K?�3���,�W����� ��^�����\��Rd�#�J�a�����}�<j���&�P��-M���S�I���lu2�AK%U���i�x�;Ex�-�H���<�N��2�P=�E�ʮ9	g�x}��f��ۚ0�kW'	��k�m2��CP�HW���OGgzP)�	������voά�{|M����*��N�w/��= ���$�������\,<�&E���&����l~�dȸ��	@)*F&y��T��}k�'����!.T��� PA0b�`���X���@7m��!���2�
�Xu����6TH�B��h����|����ߩ�5�9��V�>U�@�B����E���S�h[zHw!��a��� ?V�+��#�;?�j�����!�}m�D ��B��PW7L���c�T�|�����D�.��J�<T�LA�5��K䨅����\Z�7�5nVx�ԝ�����X��+r��R2q��;�Ϊ�iH��Pf����33��p#�[�CA|�EF�S�i�u�����Az����0����g.��!��^D���_G*��\�ڐP/g ���E�L����P��/�sJ@B�r�{�6v_�{�9Ϋ�� wVa_�@�)L=N;Z"Ċ�JA,�)�+Ζ���7�'g�h�e"9/$�PQ�8�vn�/\�u�B����*,�O��֖�ER��C�Em��w�7�S�Rr�H�ز�I_uY2Bv`j>M�2��"�!=��?/O��+uP�a?��܊I *<s
las�'�V�X�<��q,�A.8a��8mJ���U��v4��{4L�2�P�~���W �u��O:�Ŏ�` a����E��@T4���'�u=�����I�ls�N'_o�][��)�?�#�d�I���X��M�G[btY(Z�������l�"������֩N��|L�$��y@�сgԆx��^BhTw�S+r
�ӈ44/䊂bX�S.��.���n*���Z'��?���G� ��Ɇs>JR�o�	3���&u�0�ŊC��
����no�-ف�Ha�/hq�����dv��U&��n;�us����ڼ�^��LlC��b�|�3������<{OB:݌�.���q�y�*�E�b;(�F�E�;�)]��s$�������~��-��$I���j׊(nM�^;�_Wlϥ�$���;������|-����gU{x�U�߰i[O�P�(��Q������E���ܘذ3�|xs����T?����7�V�)Z�=��ӷ���>O�C�r$p�?	ę������8B|�E~5����:+��n&(�SF�S���ǂ{�1A������f��#B��il�.���x�:�ֺ7��H��N��j���Kg��,�����5���� �����Lx?�X�ZO[C|n��DE�� 6��d�k@���G�"q�W�M�T�vN9��+�<�z[���3A����&����#gyQ�~L���^�B+i��mA#l��i,����o�fN)�a���Zl��nRqx���\9�lne����@�EL`�>�:)`Q���u�;�9i!?��ח�Q�� 7ɝ�����0�������.���U�56�O�5̱�f��j��I84�FѳLg��$�[�k��&I�TB����$7���-	�C{���g��E�|`z����ӝ5޵T�~'c���қֺ�B�sB�y[��D���*J`0�ck�~�fr� $��d������� ��t$Ö|5�&P��������7�B��� �2D�[����CA��@t��S6Ӧ�����Y�o���uR�pv�b�ߔ���u*6�4˦q����׭8޿?�n�(p�8ya��b������[8��B��Ø�Y͗��Ia�} �ks�~�{���@(��9�$A�Ν�aSI`�Ȥ��s��Ӑ{pY�[ٽ�r+�~�^���	%oDϚ	��\p,�6=�}�5f��ZRXZ2�|&y�֮�������͈�I!.{����"�HN�ˏc���R�4�̏H�ER,�o��,���I�]��w��1�/�Ŗw+�����9ﲔ�X[�w�5�lb\������ٽb�hq;�/F_{e�j)��(aiS���ލ�i$/=�Q�n3[}c�,�6+��zīY�0Q��H�-�	����� ~+����-;��k1Y<�f�pȡy����ڛ����}M���Ξ�C�}���9��1�4�H���n���C�8?��e�a��&���҂ew��i�R����Xl.ex��C$��E��*����}�`��d�c�Yv[b�f~I�BG�N�����}�_!��B�B�Xif���%�|�`��Ei=��2������*�P˾(���겲�v�#D�x�#~T=��G�E��U�}@�� �_�F%�ď��r.8n9��c{�ݯȍ�7�L>�?�L���J5��mL��C	'Yi������1v���L����G�޹~����S.ֱ�C����^j��B���G`�XAc��6/�H�	�L���u�O���b� ��?ղb�EO�.?�(���V�"x�N|�(�/�U�D�f7���͇�k��l�����W�}B������@�SNlA�����h_T'b�g.����bpE= 6��P�l��.A�;5jb)�
�S�R���4qZ:7{emT��g�!N��0��b�Pk��=��j�N���C�����"����k��b蠧!��R��Ǡ��t��9�BT��@B������P������W)��;�
�=�C�h��
]U6�_(��/_o��N���'ks��|y��4����j[���)��s��I�l!X��;7D���E��V��PI��NJ"�j�>�7�_��&�
���ԧ�P'��>�s%�v�V�/ϥ�&9�E���v!����ז`�!��b_��ia�ۆ���,V錫��<?|
h/�yZ�J��#6�R4�ay���C�|��L�(��e��v��h�5����?N �ZP^�|&�F������-�Ym�8��伫Z����V�Z��3V�T��B�X��}O���M��%�KAcM��~�o�*�O�h6���Y�� ׸U$Z�z�}|��#�� �Mpe<^��r�C3EI���B�CHP��F�,j�a���%s����ML�8���>@	��Kw�yrA|?)�
N��n�$��Ү����ՠu�<��Il�YV�C�	n�[�����O*�D˚�S���-��AG頵|�lJ<u-��S�./�+�<|[�R�<�1��P����6��Vb�����t~�g�g���@�&���}��FA����kHЫdUև��zAN8�w#n��{j&=c�іB�l_M����
x[�`N_��)�,ΈFE��ׂ�-kW?�1�ՙLp-]ܮ��)��M]���fM��se��"(~zO�4,}B���V��jS� _�P~A�o��Uq{5}�@W��ؙ��WHc�aF��\�J��/9ɺw�_�j���X}��%��e�W�~�J[�2�4Hq@F���ܣ$���p3���w�v��ݬc�`�H(�E?�=%����˷
7�z�Y�!%���wiTʕ.�?y���44Ϳ÷��rIh�1z�)�����֝�����@r�> 7�1�Z�<P��v�{��U3�J���g�m�gZ}�
0灥:�� ƶ�췂����)C�C�/��/��r�M��W��_��A�P����3�fEmy�H:����4P[��R��I�5�&�Dt�eg2ͭ�#_~ݸ�\��&ZzL?��.�%���{��&��*b�O�7=� 1��o��˵�$�w����Hv8�e���-!3�
��mL�H	��3��@���;��*%�,y?��n�\���}�!(�e2���?5ܸDv��c�3�f�A�v_��V��Ll���MA@�5O��cX;���7
�k�Bre���:�8��xo��-�un��=�wb�6<�CKU��G��-h'/��8�H'^Zg�.�W�v��S�Bw�6��uh9���j14uW��L�sBO�+���/|�/��Pb��P�7O��������|�<7�j}���m���=��ۿɡѻ*���"��O\���`k�1�1�[WY���c�$�!l��	�"7J�m)�"�"U#��W������T�t�j�X����q��yX8.�1 �ZP4E;��X�r�"�%ʅA���ɋ��v �uR����H�>U�< ��qJ�d�>�g�L�+��w�٨t,L����z��/���*C��(��BZd5_,>�����F�Vx>&�W+(6�'���NI�s<V�멿4��_�O��'�0LHԿƗ�y���(���!��c7��=������܆}b�6^h)�FC�=�U�����:J�!�m�	��9|*%Ї�֌�5[��	�Z����0gAp�:���jR{��KT�k�ua�P�șT��ȃ��
��B� *�\�3�e)��!/�p�|����f�l��I��"{|_�ߚ�N��҈="�t�؉Eߩ�$t����eǠ"�����ͯ�ρ�j�\u��X�;KS"!�����}��Μ<�F���A���=�l@t�-������L���ov�zӨ�AB,���=�<HL>���g��J�A�F+Ec�rv[�d��!��a��[dd�Ɋ.�6�vϚ��yሕ,)���d�&������0�~P?��	�RХ���~��tӑ#�M�IE|ѥ!5��,jxLw3b���'�.?X�QļDtp�B�8�)���.QƳ��;��;8�]tEl�fY����Y�3�8i��Y�o5B�>��l��o�G���E��
Ǹtxb��w���s*�c�QC}���9�R�!��m2��%O�^ �،&��g�Ɔ3����,���MءU1�3�����܉0��i��0�������P4*h;��,J�H4{H*�]��=Y+�T����C��ʳ���=ٚ~�� (]���<���S���W@���T:���N�3l���5zb��K�Kv�h{����/���L��2b6Fs�hR��|�v��J0_�����Q����� �j�׾5�\fV�hw�T̫8P(UB܇���IF��|�\��1ϓ�B�H����8���I�~5g�6���pA��u:K3@�H8����� *��f��\�8�˵���N�fJ�Bte�BO��&4���M|6�TN�E�I����K�����y�W i-z��|S�&V��v���L#]�@˘�Z=�T�(��0lC%h�S�F���]�t(9Ɩ&�<8��Z �x�O����z�y��P�Z� �I�{��Z�����cV
.���O�t?	ˤB�R�]��?�N�r�h@�#x���=�+`�8'9��[���;a=�fy#���*D ��3ROK���Z�8n@�ҦGr�k���8��]���ƌ��������)o��ỹ�w����l�!t;EN�H�2�oO���3<@�����&���h'��ls>�'I�1ը����x�8��A{�|��>�Ǣ�"N[)�/�t}(�rB&�+4T�Q S�P��&}7g�,[�2/i�t&a��"�C+r�4�4cjڡkT�u���Mث^S�_iC�ƁivڑkBWm鳣5� XfbUh���-:���$s�Q��2�4��lԇ�HO�2�,,� �O����ϺK/a� �r!x������ۅd/j��i�Ǚ���1r�]�O���tdY6u���^$����Z�nx��b�}w}7�N<�E�,}yao��;���Z�C6��b�����M��g��O����n�����j��{�!���wȉ$��<��X��J~�;Mb+g��k�5�����B���ʀ]�`�N�$�5e�9x�
�/1����v�4)���9Oj�v�o<��g�F�pڎ$�v�~�g�,1ϟY�e������� �7yo� �"��ao��c��Ҟ��Kɟ�?I֘z�����a���1�WF�ݙ�#鲐kU�8�������·B�XÁ�3�d�m��~�%���N���y���+�$��QV�{�ٶ�r���F��Sl�z~�H�!� :���DL8�����?ȴO v2��NG�����V�gMy���̈˚]w>J�}Nю	q�Vcҋ�c��L.��e�ʹ{�EX��&-a_�,p��)��+�1�e�;�O�e�1���7)�c#;T$��/�� �2-�?h�I��8��g!9ٵCx��8�A�_��V���u�3���hU.�o�!q%o�m�g�O���7C�!-Rr �$�?U�!"K�^��Z�,�� �?�U�J�A���Z��/���S��~^Ф�@Ȫ����q�����~%E�9U�i��9lc!{˻�L^�e`��{�}�z�z҉��ԑv����~,��WV`X�d83J,Ih�f�X����o~\�,(�������C�r\��"4�Yt��Ae3��0��REqs��0MZs6�<�	���k*�ɡ	���������#\�	�p��@�nNk~9�'`�4�&վ��m�����h]�31�W����z��w��֪1���_��UcH֢�����Aw��)�����WGY!�ѭZ�<����h�)� ���+�w�%^a�=-�%����)��ِ���^��Ь�9����Mg٤�4��O۪�{����R$4a�e�Zus6��w�fM���%�&��bm�;�[��Cgq<	�o����%��i1éZ?�a���O��-+Ey.�7W߽)l	+2��epV���P��.t"���1��<����	5���+� �c���X����V��s����/*ǟ���{�y/��@rl!��o<G?�ξ�tC>h&Ӑ��p�{���MvɆ�ZS�ud�v�>�lH�Ca�>�â��;���A���~�_�J1�%���a[,Yu ����'T�f���'K^�������`M�谀;&/�%3��r�:s���sZ�R�
�f��,m�m����̾��uN�k�7�#�:c�G���	AR���j�� m�)\� �^e��R�q���Ⱥ1��!n�{n	���)9�܍�/ui?
4vc�� �&��{.��n
������V��~K��;q1��$.�[�Ft����JҌ䡨0��E�O��27U���w��&��X��)(zӒd��GӇTH ��p����<�gE�6j����#�8Ȧ���|M^�����F��J��v8��8��=�o=V25tu,�1�\9�KR%�]U,��J���� pW��}.�U��v�����+I��4�$R�݋(�6��eI&]�.<au3��7�� ��9vF� ӧǣ�̚Wyͳ�┾��t��IS��{;�_�J�Y��T�d�w�s�]�y�IU+���H^�)�Rw`�]��U�H���~���V��B})[�:8×��'�9����+y��t1}pMD�v+d��!�6J`�d�~�!����� ��঱\�y��.���8��U+or`��x� ��`��]l<37,���alb��e��h�L�����'m�4.k��e�cO�%���Hw������Ԥ"�%�����E(y!�K;;425JJ"�F�~������B���k�4����~��]r�+]�����ŕ"D���V�7ޞ��Qz�	�V�24$]M��aH�E�/��E��f��RY��I ��웒�f~9O�P3����M�H��>�UWݴ��U���Fꏒ��_t��0EM;���XQ]�W�Z��5���e����W���;�!�mO�]~ǚpnr�}w�]Vr~��|�YCjc�$�2�Jg�".��cW�&��H�6�1�O0bY:��=�S�)�4�O3a�\��[�M�{?EaN�:�x�
��,&�};��y�Ÿ��0�DlȪ�:}�H�>;�)�I�b}��8�C�`\��`��2��C@<�5|9Io��� ;�c��
���q��8�A���(�OWp�͵f�NR��
~���%*'��]mw��O7�M��F����,	�
�W R_7���W�jt�}U<5��0\z��&��)��h��?.��Q��J#�;��ފ���yp���7n�B�8�C�B$Z��ht0��<�M��9V�����5���{�&訃��u)Zi0����6R����?7���pl�������V�}J-x��bqf2��f�`�F�X%"��vI�&V*�ᮍf�o��.u����9�~�1����� 
�껢�F��+�r�2�7lc��Њr+����`�=��h�:[�vm��|"���.�7|�jXÿt*hnUI/�a��>a/��m"�?�:����f���/ՑJ������a0�ʂ�@�� �  f��E��J�7#a���PL�H���w
�j�Wӑqp.�u@���������~�E�X���}0Jo����Z��=OXJ9B�,�����o@n�p ID�#9~��=w��^�k4�2>x7S^�k��I�}��2&�z ��ǳ<�?���������	M鉽ب����#V��t�k�3#a~�x��V�{���;:�`m����X6㐰��c�b��7Xnm_���Yx�"����������_�M�@P��&��3��տN[
9Ur�	��$��җq��X%��T���b�<Ȓ�|2Ymuu��C�\�D}�R���m3��=�u-�5��P��S`,M���O\4�x?� �D�����|�?Y�Ӊ��7$��dG��d��]�8��Qѝ��[ĵ��PT���ʦ�~2�����%��|s�������x�EX4�O��(E�ÿ=�V�(H�N:�u�^TUyĆ����Ϯ��&�EZN-�Z���3���.��E�k��Vs�@R��ʏD��S��/qC��.��?��'���`b�Ǯ�;/��/�MĢc��M(an�c=������׹鎥����uy��� �Z. ��|�M��f���m��x].�8�/�z·��Ƚ=PÆ�<x����we�JԘ�B�i4'&"+��xe��� k�CG)逹�ڦ��J�^[Ȏ\�̺��Fin�6�;5f��Eׄ:k"\pv5z/�&�Ҹ���	+W�hc*��~�H�pvV��?e�fCqbT����&9������&���![�aʂ��ɕ:�U�'��hS�2�-Z�v�����Zۻo��1�C�m�\;��]^;�_t=h�����<B�G�C>j�UNA��*�i�А�\@UMFv-l�3�"H��>F�'��@� 
`�A�*���hX;�1J6T^Ȋ�����D9�8�RB=?�o�C6�	ٰ���qU�� tCmպ���߷�!Hؚ#Sg���e ��jW#�I�&S2/|�El���T�NЈ�~�j�+Q"���#Az�MH�%�Ơ��`r�Mf�H23�w�M�F��2����#؏د�˹�)4n;E�#Ǡj�	�KMrql��(o�Y�(|��y��ႴBlCc�B� g@h��TԨ�v�g,L����^
uN��.Q���As��p�᪗�#"�Y5⢗z�Z��H<NnI�њЂ<�1��-4(o[&}y�(�X��#�;2���܋2v�z��nK�U�������k͖�SesL�PT�׆"A�6�$*���?Ok�:b���>��q@u�����H��0�h���|�j��������߸˳��B���~�X6��GKFik�K���p\��zhM���͡��n��=t�OgG�$
��I�0(e��7�r�ͺ�Pwʓf�����d�գ��v.S���Ȇ�o�_�aÌ�%y)~S7UoJvaٺ����[	��VxC�M�<��I&�ٽ> Tn_�4�6ڃ+&cm�ڻ�*cy4��c��D�4V�(�R6 {
���M����5���0r��$��V�.�Wx�-����s�펫�w����Ү��J	j)���f��K^c��ߦ���X[B��F�6���[BKF�i�Wj�3CG��9rX:��y���H�kL{5L�27/�7��]�3s�g��=�����pE�C��}貨f��!�ջ5Ch)��T�z�Y�F�Z�Z��K�����:)0����["�p�\1ODn.���Z*N��@cj�-~�o��9[���q���Y����xJA�[�m�h�x�FА'�p��c�c�2L��>9�J�2�!��d��&��M���N�`�h�p��o��b6���8���ڦR��9�/�b_WF�RPb��Q�+���h�Z��H��=�?�
i���R��w�^@� !ǅ�T mG"�ߦ32�E��[2z�Xە8���+�>�|� ��{T����n�I_���'b�����G��1��#��r3ڜ($�G�rY��݁׭����Ɍ�&E��P��ʽcb���7�3R���1��ӏ�n�<&����q!���դIJO&�x.gC�;Y�~B�9 o�k�i�+VRc/�����0^F��(�<�@s+ZJ�-TI�>(��4�T[�sslf�Q�3S T�a�[%�m��R`x�J
�ؘ���Ƿ��+����W#����3��;��p{X����[o�^hN,O�=�b��5��J�-�u���7&���bL��Bcu����r�c}0��r,�����o��-_�EG�.���J� �6	����5q��9A���f|gR����Īj�qG0��qyF_.���9��g���V�v�p��'��>��� g��<ߨk(ol��Q�8�<2+\
g�����r1���8ӕt8f���
���$�k���]�{�Q�w6��wcJ9��i�p��Zrr)w!N�g��fy�D|��3�:u���h��h�
�8 ��/~�3H��:kz������Cm�%i�jR�#�kLx<�L��a#6�:�yxFx���{?�]�+���4"*��li�!�N�:	ډ�5k@�������i�I�EW�3�nN�סJ�L0_߻S�4��R u�P���eb���R���c�C�A�,��#��Q�&�p�tXۃ�#�����<\&d.A����d߽t�v�SR�,�Ǻj��͡Uu�p3:О�(>g���;�XfD��ޜ����Q�"���l��Կ�B��(}�Fs��S����g�_
s(di�|��_������f�6e8��RJk<��8�:A�^5d��J�<����2��� �����b��T�_\2��) \�����Ae��1��������'����ʼ��y����8�n�kE^���j�����V�>Q�@0��ҧ'�
Qu�ڥ�{�ڹ����?�AF���֜�O�ku�Sw�����;qJ����Dc6*o��}���x��~�J��ĕ��C._��>%�eZU7�/�sMy��!:�26��u��P_!r��*��^k)�O'V�$�lU���UT��C{d����-[��j[�8'�z�ݯ�$y�e*��(���25@vf��9gϣTQ.ZPY?�j�f,�v�YG�S�����A�^_c�Ԅ$��B�g��S۩D�X�r�}ޮ�ش����w�S	�G$1|t5��>Ac�ӣʥ�Ax�}(yѷх�Ų�Nn}EL�
ߑ$]ҍ�9'e�� ��"�jŤ�Yc#4��r�K�B
��աwj��mH���:_a��'��eR��(��SE��?�n�#N����Y.�HQі�X�1I
T��ӵ�N��-��?5�*FD��k�)���O90c؍��dyT(�$�g����^�J3�~�����Rk��x�@sN��w�?����<�]_�K{$)K�Ǭ�._��/�� T&�G�/�y�5S_���<�[��d֥
�=�]��j�# ����H�T�	:�}#�� I�����E�!e��1��/���$h���H�mƟ������L*tMN,
b��OG��I�*�l`&�d>����P։v�vQ��kQ��S�xg7�t��!����,�v�d߽-9�GC|J�-� =~�L�N��"����іT���U�����L��݊h�����\�{�9���r�S{+�Q[!>kG헜��u�+e�7mv��oSy���.�|v��zM�.�cv����g$N��/Zt�I���+&��ф�\�f5��/��.h~�ê��R����(#s>��J�;������#O�R_��'=߼�����P�0Sw:����$cC����s��T.�-gym��
���~���ag� �����+�� �<nz�N|�e<=����q����o�io�c��8�˫�
P���..b���9U-S�B0��~�r��*=�����>|��	5�"�] V�X��s�n�$�2�
b$_��1af�.E���V`�S��z؉ş��"gW��k���%j3�˄vj{�́[�C[͉�9SfsB#�g� �[_,�r2��8҉=��(��&�gЊ���!��/���]�����[-8��~%��Oy�*b�%K
�t�7��#� ,���C8*2_3��Tf��P2 ���Q|x`��
@ŽI�?ٶ��q>��ud0>��_
��
��NE�C�S=�1׽����R�Rk]W
KWΏ�
�a�{��^`��%�;�gs��_T6�^��c��������^-%��8�x��nӚ�늏�I�;�ݩ92��˩�;�Q߬�4�s�"�n��rb�T�!�T�Q�,U)�i�zݘj9�� 5��5���)�>�i-����w��^�v^"��Sd@1�9�HU��U��{�D�Bo%��	`�{�u�u��n�e��S�$��UM��u��]���X��=Ց���u�9%��!LmZ�x���G�V��]H����E�	��{+�f=T{P�'AM��V��&���
_���$��ܿ�7[�2m�Ԕ���v5	DȤ%��j#�D���7�Q{%����zk�W��X���of?�h�;M�gs��XwA��sM^$���hU���#�
�{���ő6��_䍈�nm�v�j ��u��#��v��Kr�dˋ�,l sK���j��Wv����qS��u#�8Ңj������Ԑ��9οl9�4 $���ŋe9���>wu���"�>��k�r34���	.aD`d��!��Ҹ�<:K�/p�C�ژ|����� ���J/��Y�[��8�Ӏǚ���
-P}E�X��bL��×�n
��>���|,�s�@Σ*m�`л��p�7���o�{�f����c��-S�1�a���:���#��9�Q:��:	L��>�,`I���8��9��0��$<�拢�����&K�Ӳ-��l��Ҹ�VFJ8 H*m�K[s�/�D�g[$�甕�|��<���l4�#��|c�!��NtQ�R���H����8��1w��<R�G�S}� ���a�����.?�(v���Vk�:�;pi\�'�^�8�h�?@� F�85�����G�!4�b[{7�['4}|����3�	���.�$uӠ�Sb�9���؊�~j�m��~S�R^ ��|��W��JE���z��5C-��9U߸e�D����rc���F�������9alF!T<�9��ַC���[��r1Yߞ�-l��Nڐ>p��<���=�P��"���_�#�Ob�RAܛ��w�!hr�Q�vq���}pi���Ah�,��Wb�d�����A���6�T�X:����Ϣ�#Z�Gk�3�%�O�)O`'��R/{�-�6F����\��z���̮�;���D��������v�O��`�r~C�!�&j��Fl�8w��7���lsش�]A�hC6�N6c]���J�8+��+O�¾�m�R{����B~Dxl�Y4�=�����C�1ݺȜ;4�E|
G��9	\��-f1?���#�,�����0m�.����P�-8�a���'w�ژ����q�C?;�rP��$�Q��[� w��m�������t�dɉtJT��6s(Y۶�Ȅ'����� ڞ�����-8����6�@4���h-v�r<����EH�j�RԮn]�MF�
Nݣ�+\��\ߟ�U.��+)�>�.w�ɬ����T�S8���Q�q5W�2%����������]Q��$��U9�a��O>+D~�����H�@��E�@�5�zy(/%۰��Do�8:�0K�~�UO�N��β�y߸K�(�{�ra�H�r�ߤL�J!ܫf^��y��g���Q����] ��&]�Lm�N{�����Y��!ww��d������Ռ՝���� ,9�l���&z��-��U��y�H�0gO�D�k�m�[sR�԰0MXq�I�� �Ƶ��;�'�x������ �5L?����g9��#?�U��6�7�$�w�ϼiW����a�#~'���,b�뭌`j⋀d��]>�/�r���i�࿖Y6�����Q;�ԣWb�E�������r:�v\M��/T��o+�z��:��Ie�"*m�g:;rx+���w�n���t�R\'����͓B}�=�P�u�S�
7a+jh��m��G��NE���G������č��1!�U-�����HC�����������=��\*K�Č�Y�ya,�j1�)<^Q>�}�_Ù�W�6�!����Lc~�y���h�Z���Ņt���af��F�J8�)؊\�X �����p��9J�jڍ�&�*w^;�;��,��~Ru����c�������q�;'�(���ޘ.���_ܔ�c
V;b|��E3J�T������K�ջ�!fh޷���Q��1'����e�A?��AI�z�dF����-1��c��rR�z槀����Mfy��fQd� �����[sފ�����#�E��A�.5�$*^�g�ш�v��Ȼ�P*. ��ȿC��F�ưw�O�e^�)�ɴ�P�GF��>���{��H��i�G,Q��^Z�]�o
������揤r+I�d!�}��h6�3m�K�^��ی~�6J�xF�`�3d�ӓ�.�z�舊�u���B�d��`�!�b�p>$K��b T �L_z�	Q��s��[VY��m���g�C�s��j�����R��hW��a���קcU�Pˠ�1)�Todԫ��_LL>n��n����h�{�>&)+���	�i����~�rz�$9�K�M��6nJ���|O�q��o�����0��@��c���ڦ�<�����F5����-_�n�?]vO5>.ӥ߰L\e�g�m�OE�*'�?F�D�f��:����I�<7����>{u��(�U����aB��m����?"t�]?7��d�j!ȓ�8:24�2���ӷ���av��r�?��M�XMPE��/��t��e6�U���(c���J��1b���ߑ$�3�@P�N?�J�$p��}(H{&�fI&K�hv�Ve�Uݟg��@�F��s��YN�T����<��*���eM�l����Ul,�j�9�`��7���
(m۝� 0���5�O�>cM*,>��:D�ۗ#����E��g���B�=����Ⱥ:7�k�ɉ�w|���a�ed�,ů����CW�XZX��~���9A��~RtSݛ��'��w��Q^xf�w���&��<�PwE�\�J�R;5��ɘ����hF:��@�D����Y(ҐL��%��o�;l�#&� ��%��K:��8C�4�[�R#�a5W�4�r-�B�8=� )���&������+��_��>�:21�u�瑶&Q�ՊoR!ԥ�����;��\�I�q�$�� �bC�M�+���϶yui�����4����ǞM���[�(�w�� Q���U�ۻ�;&��e*��A8ǆ��j�tr��j��B��3{%�o������na���`�᤾�-a�ǟ�f����)?��Y�y�`�O�z�Uv�ʦ��cP>KzJ��o� -�|���q�?_��#kE�v��L.E��L[@�O!�Y�&%�>T��!�k��^�T�֢u�Ɩx�s����K@�8|���w/�%������&cǢ����-�нlk�y̳���=�� +�Fb��{�Hp~Pq�w�|�H�o�;9q>��"x�W�$�\$m[�0-ք
�szj�<��J�6ah�߂"�Q71����75��v�����Ƕ�+B~�7�:�.�S�ɾ�pd�G�^��PeŰG3@��چ��缚;�T�4e{Om A��%F�q+��V�;�M�h���5Q��'�G"������g^%�IرJ>%hҍ��Kp�����#�Z�ƍ_�R���1��vPd������O�����6�j�����`M��mfn a<��tDK1z��Ho�tZJp
���n����b'o�g(�0��+>B��lp�e�̉]}
��f�4�|�/º�(V��Pln�Q큫��c񐿽8�?}��2�56���v��v9�֍�f/H���C��������oE�?�Q�b�������v�z_�;0������ja	�u�*�w9�g�D5*&�\o�B�'F�2�(�� �I`G�X�-°��l������3sp'&��MҶO��Ѷ�b�P�ʝ����&"�Qgܳ��<$W�g��)�"c�ZJ���AV
r�xo֘}��kGlW�
&n�啕�|��mS�yn.�C�<�g�{���?���cq@1�(� �i��j����&י62ehM44��)�=`D�2��}YX��e��*_�N�D�o/�2�|�}E=B߆���	�Q��w	r5��b�mP<�q��[Gs�~;�m����G����қ�5Lo,MMVN&�<\�_���;�yb��^8F����\L��!�ɐ��-�T|��<�g$��]v',�̃J�Q��F���zj6~{.�u�4Q<�S�2�&8Rԟ�Jjh�e�m���
a؅���(�'i�J~�����ф,c;�IDĲS�}.�@����#����j ��8�s�,Shcaܜ��ZOt&"+���᷈=�mo!��pb��[t��7:����ј��dC�$IqV�ڥ�v�����vJ���PvL���2���!�&(l_�*s�ȅ L��<5���Z��Q���ͲF�)�צ�bg�7��AA0�AGI�Ip��Pe;R�#6b���S��kqD�����:���x{0��<��0�� S���'�`��zɰA��jmǮ_�h�)����1�$:e*�
�� �}J(I:)�)+u�-��*C��=b�F3�ZS4��Z���E�V��:���U�L��]1?��XD��d��i����xɢ:w�4�����]���[,�O�� �j>�D:�7�S ��'$�R�!'ϓ�s����Ƿ"��\�hU`��~\u�tt���(�v��$�� S^GL@|�(���[���<�>p>4���-G2�-@�[@�0�)�G�Z�d�Ӽ5����T�2��ÉPq�gϝ�4�B�C�蓘�e�od��L�S�s�[�	������ʡ�UH���������9����6D2ٸŠ�2���p�H�A�Z3=�G�݇��}���FQ��D�]�z�x���׌2=.(�������84N�$Z��\P{��H�/��89R$^Y P �Y&ǐ�) s�;Y'H�'�7d�����SS�ه$ү��|Z�5�-6cmE�m�S�)E���.��$��H+DLȲMdD���l:�(5cX00��]c9��m)��m6�q�F7�(r-��r��W�͏Ħ�7h�����B�1ǟ?yٗ��vju�Y�z$A�)Yn��t�L�*���qw"�E��Q�G�!���'� G�E�Q�܁f?�@Oy|��v��e��ޓہ*���O��s8����\���j"-���7�_��Ճ�1�~ͼ�"Hh���s�u��w�M�)C:�9>����.6��S�$�C�{�/EQ M�_�ru�h֣"21�J߻���T�d7y �Jj ֆG��ZOW�ͩ���A�]�?�C�ܭ�sN�!4+<�A,��/_��C�Y��n���p~�skD��GP؞�ƍ�wc�(bx1G,x����C�:���Oϵ��-t!ݶ���2�Aq�n4��˺�ؽ6X'(QO�z-˽�ӄ�N=I�����+X-��/�3W��-9�����4M"��3�Mf��pɄ(r�N���
�wk��-`N@=g��\������D�p��7B$6���h�I���@ri�ֶ.}MG\�^Z��?��2�d�:*�洕>Jɣr�J�1K^�.�¯���{O��
Ms�ʉ���JŨ}��V�i��
C��=���ͻ�I�D�%���jz[y�1a �ՁD�<IgrJ��J:@�>`s�U�8���X���c�*\�DF�g��hA�͍�<c�H!�H�̇��%hL�Zm~!͑^y`~a��rp�X;<	��c0u=�uq�����~���}�|W�G4�������q<���:4�(�w.!�R���KE7
�K�q��=w�j�><i�Vߎ�7���?��4gE���_u��� DY��O&{����u(��XK|`�	�Xvj��Յ#K���v�/�cVob�5�ϙ���E���
���U� ����ێ �yA�ܦ��|�|]\�e�^o��GP҇�Q����y�q��|L���=(�jmE�
�d8��]�WW�}������ݰ��o?�ڰ��fĕ_��'&5�ʚ��=�^�E�b��8��n�N(n*[�R�,�;�V��ػ�1f^�z��>��t�����p8ٗ1)l>����dk���Y܎�w��	�E�*������#F N�]���%Q%-*�ZC֚~\!�Bj��ʵ?����P{N�!�ܸ�#�|�]@c����L0S��:�k�^[W3��̒��j�
�隴>;�D���S��k֘EE?b#HP�fv�MRI��j�a�m1��N�۪h�6tM�%~/�#\b5��s�x10jN��6�|����t��KANa����"}$Y���}	!�����/T��|A!]���ԛ�F���<�hʾ<���[y��h�:��3��9zR�Ag��f2K6,6�+C���h�����<:��a��a� ����/�s��0��^Ԛn+�}9��pI��,):�������}��g'�T�3���H�[6�+>�eĪ
ߡ�&����}S�ԗ�ʍ����P#+.� ] �O��{�u��u����A.�0���̊�ի�������#�Fr��@���j&Mt��c���~yr�%�$�SJ�'X4�����T��\��Ů��P�S��<��+n����;v�E�?U�E��u9�`V�{>�2{���V��l�W����SZ�n`�i�]�к�������r�x��0�.&J|���Q��z���M,�z:���(\�����	.L�E̼U�Ŗ ��ܻ5m����j��8����<�TX"�+�/b��sJiF�')H���˝42��F���MI��F�d Gơj� $�l���S6�"CH����\�ޖ*�K l3J�J�Z�Џro]�hxA�S�����*A�esM7ǚ�'�8#�M�ZF(��� t�R|�Hp�n���V��Ҹtk��|E����K�.�Z���s�J(��@kF;	���C����:c��3� ��Yp��-;6<~W8�_sQ	`;��Б���3�ظ�c�ҙ�a�#�F���;s W�W�U;�gJB�JZv��E�.B����W��3���l��V����Y-	���c��K�T�3���|�tP��J�0�U�n���kV�t�f�s��z�s!$�.-{�c�|�~�*-^J��Gw7#/ @���tް>ט!���Ú RD�B��K����q�eS�=�	��-�rTLZ��Q���8�X2����HP_EwEt�R�>@�O�4vݾ~|�R�7��9,��^1Kbm�o�x��i��6�����������7��j���
P��������ʠq���F}�kV;)N�<k@>d��A5*��90��-1��E�{Ӄ��u�d��TV]��~���X�K��{�x0u>�ЇΪ���Vz6�10t���6��Gp�ak��~g9�HM\�؆O��9u�m���(��À~��'kKK="��"��Ri`,��-J~b��C�DS�$2]��&��Q���^3m�\Z~��r��9��p���'®��������J���Qi�Lõ����H�>�A\Q{���gb�i.ݒ���*��	���%�y �� Z�%��v��!�q{�����?��:���^�����!v[�*����J��yļB��R�X����V�Alt�_W )�Z˨K��gibB@ "�}#3�q�!��+?������i!�0�l��wԊ�߮OZܪ��5��j�'��ЍU�b8�j%��q���w1���T���R��l8Ե�-x��WL9{�D9]g��3�.f	���?|X��hA��fMz��9&����&��ľ�q�r�u�c/�s�X�	/��)��x�/�=�&<�^~5 ��`�졮'�0&�5+��(��쥚ٜ+H�U�_&wPqê�ZُZS|���/����/�x������U6ɪ���ۣ�TՁ�XO�;�/΋|�_���ʞd������� =H�s���b����"M����J�dOgFR�h� �hq�&d2v�v�ڜK��ep2֫üc��e8;�;#�s;e)15J�o0�8ϥ���1�]1%�Z�?@-�޵o��Y�2:8��x"����.�J&�7�����t��M�H���&��M%�Z�?��/�FP�?�N������6�LYF��#��w;5��=M�&V��,��6=d۝�)ER'��i�ՠW,��R�" �EP��Q����U?�C�2�g+��Wu��6y��^����!�Į��݂L�^rJ@�~Ѐ�X9$�4�Tt|�q����H�Hʽ/�����Ll��gN��-%'�����3��!�.H�,���2ٱnI#�eT)������~E�-8��}X�����;s�"���G���zh�=�"����0���>�K��&�%��H4��ع��[؁unU/��U(H���b.���F�rS�-��8L���&��t�d���4�5i���v�i���iHRV]�c2��*~O;l�ze�j��7���rk�<w#�w �����X��_�3��*U����S�̓� e#px.m�ʩnR��H�r-�P�py>u˨E��������l,.c��߷P��0F\1���
�L��"�Wټ�KJ�R{";):��;�E�՝���On�ʳ瞥����5C7ڗo��!�b'�ё���b���lAG�P�-7ͧl�I��qR�.�x��MfD|�r'�ä.=߈x,u⠝��-��_=��G	��bs�f��3b�NSTh�����YOG���o��+
4�a�`fG�˂�Xt!��tCr���u:h]��9&v��;����=�-��!��r+*~�����Y�$G �)��9�~>��ET�L���Ǭ�8��Q~sǆ�r@C>��n��r�z%g��d%k9_*ۗ�$s��?<�lY�|""c�^	l��y��)-��6��M��.������Si²�Т���bd���|p�M�����)�<����a?���T�����ob�2,�������/=�׼��ߑ��h�3>f��o&�Jo���rE���pc��̇��b�C~10���F���[DgNٺ�#���Z������=g���*�)��N�a���K��ߑ�n� �O�,V�Z�a3!���6s���_n� :zu�	����T�9���)�$mIc<��N�,���#�X�Wu*d�q(�.=-خI�y�R��kL�w��@<b�:���juUCy��ş����Tb��w`�A۶$7np�\�8��V��c���
Ft�h�BF�2��w��7����UD��WYe���E���l�A�Y�Q��#��C<t\�9ܰ �_����.:�
A�/	L��ᆓ�z������h�=4؛�<��ew|c�� ��h�8uD�g��Fs�{��i�������\ÙA�0�YE��ji{��
�����;�?7��>iRձ����A�(Z�	z
j�e���2��8Zꀀ7K�����K������m>��w@V$qS�~g���w���в��C$��.':rM��b�D���hK��4�1�f@�����X8����k��#+[4��f�z*��x7|�����I/Q���eki�����筪e��蕜Q�͉����Ұ�p�E�H��EK���M�P�'�H���cv���<�3 ��rM<1S���쒀x�&������@}rl���}�3�]nhH�vVx#02��++a����d"GH�n'̅^(|�)�W�%�Q3;��d���>ʣ&�hb�r�M�/��&X}� u��ˋ\E�P[cw�pb)�|!��v�:��c�3�#U�+
H7ډ����`aJ
����%O��s%��ic) /#�dH�8-<6<k�3��n�:9Sة�(:����m��k5������-hʹ�}6���@W�r�� $�=����S~n>�h��Ŷ����Ť!�kAK����Ǌ�����
8�*�V8�9�	��n�EVq�I-Ӻ3-H����X}��,ʺ}h�=�4�A��oPAbId{gפ���jطZE�'7��Fѱ�Q9�&�Y�'�U�$���%1A��E�����.=:���?0%���-p}+-����39w�2O�����[򛂥g{��|eh�aMR
��+������As槥�/�%�RS�9O��J�γ~mt���,�I���a0���A_SX�!2'�Y�e�Oq�3лo����V��M�v߿96ǟ`��K�
�f {���%4�%�֋��j����a�D����%��-]Q��&m�:?Ts��`*������mL6���q����ȩ�I�;���M�DA"�-��Q{t�b�G�I
"VA��D��7 )O��%�O���$�Ρ�Q�#E#||��>H`��;	B;�N��{�$'K.~�Qg�y���P2��t³'_�~�@�&o5���P�U��`d�Y��][���⸻�WE�契Sj�I�I��)ڮ���{Ƴ'ʙB�=��
�q7�O!��煟ɏ,�O�d�8?v��~��ȅ��I��^���R�:����Q�V�R��"��p����6�~�v�jf������5��m"���-aec~Yg�Ǟ�D���&poo�� ��&:��tl\�����54��#F "*q�Qi�%���=��<4J��8�ו�{����tǠ�'�I+�c~m�v�:�e�ʍ��˘�lo��.��j�-��/�Al��}P��$��?H��,Ƞ�?���`b���t[?�+:Q��u�NV�e��`���0�g9G�Ȕ|�p�5���������ɂ(vF��Z_]���2Ɗ��Hk�j��'�s��_����h�9���)��_I���X�i  }�����;�x�N~,����j4��p��ɒ���`���'?x��D�2���Zq6�/��I1�L����(��5æ���1�ָ�.�
�f��%�j�|�:b�]1�%�n����?jF�KwFE�� d�@�c3,���5^����H�����)��=�A�j��Ʌʷ���;ԋQ:��U'��u
4,��;6 ��$]Csf��޼ͳ2jZ�ά�
x���"(LĸXK��侠{=tV��[:�;��b��k��g$�Yh��P��J`3ƻ�]��yeΊ�(��J8��ݮ�K?ө�u�wdWt�DAo�W��A-�z0�=��G��"r��jE��l�|��/��pn&l���K_8ec^e���w��U��lS5�9e�W���]�
%��۬�Jy����S��PΞ��(l������;�:ƕ
o������� ��jh���8K�Y7�M>e��Fp�_�Y��:m� A�Ĺ;2XM}��)�����J*�q筃(�!'���R� j�(��������������1��9��b��J-.ޓF�8+�@��SБ�Gk��O,�fȪ�ya����Ou��T�����q�:�3)-�Ūc�y�)��0�F�Sj��c2tW�m��z/�N���X�[��R�馓	J;���v|��^�b�ў/K .�>�bxI�ǖʜ���U���h>_e��ݱ����02�i����IE ŧ�6��\����� ��0��b��L�2��#� �VS�|N��9�2L����
y�y[�`[�zab��dc��'�����.N�$<B��I�6�!�i���&
g���q��s!<k��w������u-;囯��H�X`���~0��G$$��@��s1&ɚ�:3�p��?F
�{�l`��BqJ~�� 2ц�\#�ߒ��{�/�SG���q�ҊC4샇�6U�b��V4�:)7�0,��j}�ɽP�*6����nj$h=[�p$D�@��QT�$i&i���쇪.��m�dn1��q9k�.��#�_����Æ �3��7�#S�u#;���BT˪#�5~^�L���G%�M�8nꖈ��3zxg��Q�W�T�k��5Y��É $Bg�aX%��.k�"s�d���k�� ġi�v���7���8Ӝ�&����Bx������*�h�U�R�g�?��|B(�]��E�
�6.��=�1��mg[İ'� ���+4���w`~�[&���tw�TfJ'��#)�"��ߤ�懧-����Z�=�q�O�?}�|D%������R��j���S�����rB_}�3�p��]�.�@Meg{
P ��p2�$H�0}�	�Κ�̨5j���kd��ݘ�c1��9������C��c&���3���:<� ��@U��i��{,oлr7�%-$���j.N�!@q�,�v�WP���K�6,r!J3�|���A(��x�d2>ZT�0�#	���W�	�}�E�l��$��� ��Uޔ�g쩖w���	�i�꽮=�;��R�ۓ	���/��́��4���=�ʻ�)oˀu��]�3��U�ר�Y�ʍ�[�e�r���Ϟ�AI��J��{V�����!�cQ?׸1������HA���]��u&��i�!7�7)Yĳ&�-�!������8G�3ě�0k�����*
�d�{C��@8G�t߳#!�Z�6�F�ML�{�1^�#�*�,�S�� Û��*�� �Y$Ұ�t�"`i'�ׯsH�H �`Űߘ���[�L��S�^�M�`�J^��ad*� �E���&,�X�
�����<���G[��0߅��r�	s�仜mJF��"<�j�����MI�-��O������U�`�%���Ɇ�<�{�y���'r�#��Ho�5��O� ���N��x_��w�X�F��5�mq�Sç���b�"����mG���L9�D"5�LΣ��k��u�ÌT�#���kcO�,��9
<����z��z�^���IM ��8N�tS��C��� Ĩڡ�ʫ�T���ߛ��ya��Ky٧0SY\�,�ߪ�3�m��&rLdKm!;Y����U?S���j<�f7;�V�]k���VU�:��^f�u��U�l�o�/��D�a�w.�ˊ*"���n��ap%gƐ�@���{����O�Y���V�A��Z���C&ZX�'��7��7���8��+\�l��V��!C��艗��u%t�˥~��NB/X��Q��H.�j���5��QVq�|S�&����/�ٸ�|�϶}�Bq9w�����2�����r�<��
�8�<6>pLS��b� ��aƺx���E=��nP)�e�����ުQbr����ғ�7��OCق*T��M'�f �~MQ�
}: �8F�Sh��k��֘�覅���z��
�SF=v����^;v�U�� F\_��b�k'%�UN�}Y���G<>Ĉ����ϧ����qޏ�����|���kͦ����"Y���
�W}�����Ԗ���8s�.�>���jt!q2
�p��RRo(mAv�|�[�QB�V5nne0d��f��8�h��uDeVO|�~|52@���w�I�冩�k���vǽ��#�硑�h*�8�/���Ӑ��R�Z�{� �>�w�,V�'�����Z�m�������%�d��T��z�<�t��Njw�6��`�5�D$Dx����BC�ш�׻N7��N�b;����.�_~Q�J�TC7�8ڑ�k9���i$<����jQs�l�r�S_i<^�o}ݢ2�����L� 3�,4�$�I$3�:?��G����#%�X~����A
��P	Z����6hګp!�ni��Z�tV�#;��!�����|��x\�<WR)HUw��F�)�!ؾC�Ù���3�֍#O���i��Q��Â���I�"���*��Ս�Hsm?\ǭ(�+�Q�!W�<��ӡ$r�YS^Y{��("cD�l�I��M�|�އ��D�\V>|ӡk�u��&xd�|$�UR����ƌ�ϟY�U��:1������:�K�@Xƌն��{�k%���Ʃ�mr��o��+w+~9_%O �r���#�QF����K&�JA��@�$��߆�`w/m9���4�-mX��]k���]��ҙ)�뷗�U%sCrDʜpG$/�=��������%�Ju���7�#v�>2�N��;�$�+�a������c���IS������� {��I�F�ȏB�'<����H8�L���*��=xg
��>�����9΂�� ʰ<��tsX�R����{n?$�WϢ�|3����(�����y����� �GZW��/ߜ���j��۪he�8�W�=���6W/]��8�b��A>|?���-vy<%Փx�d��u �U67"x�XT����Ҷ Js�X��|�v��}XD�B���� e?G]�ե�j��Hn�t����['�)+-T��i�^��:��_����Ob������rT��
����N�<{�U�*��~g�s�f�P4�[�J�`�X��WN�����O�2��`S;f�혹�w,�m�݉��&H�����Nض/�4���_��v�5J�:���Fvh��|%Q������z|+B�h�X����8�	��R`�6a�V':���u�������Ñr}�~OM���d��_>��1�3o��K�}4B,��jH��l�}e������2	�
yP�l@vM���vDj���i�U��T��$�T�����v�q�l ��i�师w���	_�ʋ�)p�@����w��U���T|(��J�w��x���K_簧��
�"�b�R�ց{���Q�C�p1a��ڕu�C�����,VC_<��h8b�3�#!ʁ\���������S�aŬ�טD�u���(�缞m]TP�P-L����,~Cua�GL�S����"1��K����t���/���B"����Ƭ�,����VV&4��ݒ�b `�.���0
���@#L=cWe�S.� �Qi���� ���H3��y��{XE�cr>������׌��� �O'��ݞ�1Ƥ��ei��}W�Rո�^��}�6}�Y������W��xt�Ф��^��t�ۿ��8B�1��(O���3c��rsƹ���,�GcOVU��f� ��^���d��S��4��s�9
�:\���և��\�s'��������ja�T�:��S�� 'Kɵ7M�׽�r�[��R=�5��/U)q�����{��j}IE
𛅺},�p��}�h?P4�fF��Oj�.
�u.x���#�6��P����N��Ru/��a�tϓr/�`�sK��Z��x��Dמ� 址�Mnf������k1��<v�
���[���4����6�T��}`)]χ�*��Ҫż��I�pj�Ie�c��	i6�V$�ƌ���5U�h�i��S8����1�vy�pG<ƣ���!�iZF�Yi�b��s��b=(��=b%�0�Y&ڳ�p���Ӽ��Mj�OU�Z�[6�z��g�k�u�^	��6�_�(e�������>�L{[��z�� �/uQbuN�K�7�u�v �W)+��g��ul|�;aK�ahŉ�6���S�^L�3`�p�'��1G(�$4�4u����ĉYc,��j��M(m�80����t���U9��0_xφ&:�QU�b�nXEC�ZIb`�_�����)���W���X+|��1��l��]N��uh?��ʜ������*��\Y�	��U��S6�M�j�6��MW^C��H���D���od�z�C�%Z8qZx�
p�f��|N722�PX�J�"c�ϺT��j����Ų�m_��?������Vw(�T�+me��t*2��1�滐�v�k��{����m_7?U��omp�}���׼�tN@�)sj�Cf���h������玿��08�Q��";oh��� B8t{ ��l��ٍ�3׎�zU�I2?�$��A��^߇�Ǡ�}�i���0θC
����$?�C`1��Y�m2,J����?ō�X��P[-�v���/�6j<&��r�j�O�8r9��W�@�t�ax��Ug �1�!�T�Q�#m=e��+�6���b�9R^�F?���ˈ�>�b˰�y���a��/��Cۍ[���y�{.��qZ�8r��?����ʫu��w2 ^> �����W[2�A��}xso.��c9<.����7$l���hr�n����ia�������O{t�1u[�-H:"�/=_;Z���K��%�Vd��sxdŜ�1�oπ�|�	b�L$��II��M����ר�'	»*B�m2����t�j�3��H���N���K� ��9��,��g�^�ŁiS��nJ/X!�����$xWO	��͔�A�P+̖�l�)��Ui�Uot�J4b�QM�Q3���*[k���9�� ���@��q���fD
�k�ٵ�^�!��I�Fs�rU~���ɓ��>��kS$�M�����B\�^�������.��}�&/߭����b�\��'-J�-��|w��V��
4�70p���kxdx-�]�cKPW�AC���79�_Ic]�;3r���A��� ����QY�1�@F|�"��]�TLN�OH �i�j,�k��ϸ��Ĵs}�Pm�o�@J�t�#��%���C-�-f������X	������l�E�jP$r4���Ɇ�5mݻ��b^?]:��s��]���irm^��@Z��v��/��&�P1��=>n�<�x2^�[���ut�� <T�sl3�Q�]T��<|N�������O��3k����_����Oj�)��z� L�jj�/M��i=6�0���l'.�3��C.��u���@ف8�w'����5�u�G�8G�Tj�-��ŷʐb��qj��/�t���N��[!h.Q��t7�(�O� �!'M춅��QWg�8r��%?|5�}��Z��"^�'� ��Yݧ�
�M9�'�/h!��c(ﰗ�7�c%n��@����3�	�wK5��4H̰e�BGO�e8��ݜy������a4b��I�Ρ��� ��p2?���cC]��@JFqb�=�V���so\G�x}ᮿ��J1q�`~�@�o�W�ߐ�w�MF\G�<����U��<���\+X8t���>���~�q�*�q����Yz�[U�E�4���1Ҙ�3H��4#�?����k��h���σj����n�䟹��\I��k�oy;��i���Z��0�a
�2>f�yn�O�
|���T�;��'r�"fK�·��������*M�j��ВO,YF��C�9���L��P�>��}=��~�����K��xK�� o� Z/�p�ݻ7����6!ǃ�����2���₤%6BB1�k�Ԟ?�w��$��}��	p�L�II���L��Ϥ�-�1m���*�\�l�hﲚ�NF�=p���|�O��>IF ��(��H���ݩD� "��L�|zi�T�Qe�z�SG���8�hkd���
#MZU�+�E�;�ƿ��}���_��{��P���/�Z(T�W5<�߻���(=�u��^x�Ro&)��8��vȇAÝ�c��K�"#�1Il���ɢ��ٚ!/�ঈ5����K��wa��8�G<MH��?��	�]c��C��<^�X���,���.��]�g�+*GP�
m�K`T&�����ď:��*���zE�}vN���ա�ZD�ʎ]�l��M;L9v؎ɵ����S_��n��L�Z?�f%��f=�_�
ވ���"�ᴠ��ҷ�惮�1�h$J�!B��w'��gqA�����ǽ�7W
$SK�ݙ� H&�o>�uTߺ� �`m��s��sa�� =����׵,%N�3ġS�n��]O!�B�<)}�Ga�G7�F��O&
fh�B�Gc��,@y���?�{�6�7
'�IG�r�{�����:�S��S��j2r�3�6�646���0��lJ6��,�+>��)ؿc�u�x�]��E��>�EԹ�7xA����o�z���վ�;�o����ol�Ã�^#���4��6sRwwae�Aٽ酣	`�)����J�J����P+35h	D��d����qg1����}���3�,b���oR�;*�s/s�!��;��*<�n�{���c���@*�����v��nc@��
�F'U6�2j0Y0`�������O ���T��@KΏ	tփ��*�^k��7�Lu7&�+
��t�-0����Or�N곌0nwa���D��m��1;W�
7�?�3���� ����u�&��g�\��t�T�*(���&���t�#&/P9��`��qK9#e���-��)��L�W?�>Dʸ۶��꾆p���3�u�ru��O�VA��!��<pn��Q쁇.�f,�h�2c�k8�-��RX?��k僫6C"�k�Nts��񷼴��oz�k�g����ֈAQa���2���c]<!���L[�XKa�Y
�8��F�tk��@�ń���JpA�uWN���^!�O5~�i��ٚ�A�)� �{�E�:p��~�a�/�����=�
*�Z�����Sj�N՟�?UGz9�
���n�8�$ڒN�]�ᱡ߇�_䦶9���<Cj���s-�4Kז����͹PU]L5cv]�Z�'����z�ds-�u��Ϛ�ZSu���'�Z�k���/F�8���[C�,G�W;O�D�,��g�HSG�6��M�ϝ	�B��07:6|���18���,�,�XB���@:��Vp[(�U_z�) N�{��C�;!zi��d>|�h�;���HH�[Nu�u���oU5}5�A��0�S-D�l溩�j`g�|^�{6�G��٫й�7��|5H�Fy�Y����c��B>]m�"�C�b2�2S(s�O�>26���e�`���N?�=n���k�I{��%�(~O�������Na�n��Y�|��VPӏ����N�$ZR���k#��Hw}���{	 � ƈ=�2h���k!�@`�y���@�������d0�&�P�i�S�	��.fh��M�Ua����W�w0�H2ة,M�]J�w�1����X;�Thu�Us��:�߯)�V�t�� ]�����HFcQ��wz�.kH�]rR��T�i�䫯=�����-��`�h4�GTJT3�s��h�\�&I�S�O�u	��x�yzV���'�)8�'����t�d7��^0�r�H�^p��u�������P�6p �gB��^�S�����k�k[xvP����o4�� $xT�� �y�Lț(A�����આݵ�r���4��ll蹢���H�m�َa	�wj�e�`�1�� q��G�:�kTFe쬃;~�K�+fٕ�r�ۯX�,��$���Մ	{CG��nl���A����y�a��E8N�X�֟y�KYv`���.x����C���mV�~�5R�"���#��������G�0�͏�2��/T�fn�1>8k,��(���`��1"tV�[��-���%V�+�cޚ8̏Յ��ᖾH���nH��S����Sjl�Dj�!:7D�|��b�9`�������,wm�u!��gJ���|�N<�
r�z��Y�EFW���(��Qi_����V{۾�G�]+c��b���ѷF�>�wfkҀ-�d�n���� �Ë��e`��V��n��S��67U�T4"W��o��Z�[��RWZ~W��7��t�������6�)9�Bn����e��SH/�')>겿�Ɣ���Im��j<x�t2��eo{G����_yΎ3/��h\����[�����Y��ΛY��S���8f�l
!_���!�4&��p1osդˉ��U�B�����P�����꣑���X]_a����Jsu22{)�|��̀s��t R=��8�ǟ?V���-?�=�O��X:�D}'՚�ݳ���sė�E��N�m2AƳ;ó�Y"k�x�X��3�U������fc�4���XU$u#K��@���W��5G��%�^�h��9����u�94 >8q .NE_8>��vg�%��'o9%�ި�Fy�;w~ ��R�j�vX�+�F�A;��%�q��CA>�Ff���bz�z�}���U��dYQ�B�j�[l��?7v��/�'��+^��fZl��2�99��z��Lr�s��^?�`�8/�Վ"��B��PfyO{��ƓR+F^���wی�\�+j����f�L-a������^�ΐ�^��az��m-�v`���N�0�N2��镖-G�p�Q=�E�B�Ͽ�k�/�Qx�Ӵ�a1m��B�V�P΅���H����	��5T֒^�CeJ�:��`�)Y�G�Z��K�,Qi��k���-L�_f��>�4`�����U\y������G����l�\'�Uq�܏ܯ�8G�$�\V��
SP=��T��LƢ���5��w/��B$`��2ϡY�h	�P�I�X�a�̤��ip��ۇ>�i[y�ʳ�1r���X�����F��ȁW�47�^���wp�>#��sz��p��<���e{��F�h��s1�=��~�m7���[��D*gˊ�i���(��*mFseXe?@��O'�<϶"��zh'mNg�1��(�=��O�Լ��^��(�����iob����P@m�o&�P��,&�s��6ua[�_>�<N&\�5���!F8o����R�e���������9����je<��\KM��*_��Ѝ�~{��.�N��l�RT
������pZ�.�NI�OR�Џ�"-P/������!�z�rY�����2c8_�i,��%��2��L�A k�.�A�v�6�n��)8B	� �;�A���V��Z�$�'K^���D{����"�UF��~��W�F��e��^wy%�/�&��f�ɫ,譓 Ԭ=�Z��א@��t孤0�d�����uX��xGIӽ}+Խ�Z����<�=ʵ��$v�֩�� �p�Q��3#T;a�8�L��$ɓ��ZOJ��u�Ɂ�>y���D��P��Jj��!�K:�]{)7!�
�^_ԁ����͎g���k��#� �٢��0Z�����@߀��s?��Ir��p0"4@�A��?��ß�w
l-��q�k��k�4�g��6��<}ٽ��Fh"���[�	��F�כƸ�w��	�Gp� �U�J�jw��Q����4��������Pi�wH�K$�p�.�����RK�{F!����'�3!�{�膟fs.����e#s�����r�G��@�,e%P6:s�s5��p���㊱5:/�z/�{<Ḋ�A�w�䇆I�����K� ���I���v�h��,���T�Bp#����� �������Eڤh�X<���)GlQnѣ�Ɯ��,�*�̌��e�`���߇#�k3΀}� ͱL5��$�T�Y����
�P����CKV���g2>5z'��c|/]*�q�3�-�V���ը�Iz�����<}��Q%����ѵ�qiG��̈́�jJ�N���겘�I�
��7�&�y���ʶ'�Foke L���Oc#�k	{9S(�.��_���n�U����_<��Mh w)�M��ĘW���U����Rl��Ϡ�oA�W��1G�K$��SwSc��[J��P�C�7�aXjcG�Z��F�f}����F�ֻ(��wP6�!�'�1�-��~W��\�lg�5h�c��n0�����`��Լq�\NW��o�W��oڮ�d���'c��z�|�{ e���� ���N�K�P��V�1��e��|�<H�'�Ky����&����뻰�v�R�9����n�m߽����Y���d��Sz�o�5%�t���ˊ�ON� �P#``�flx�k���=��'g���L�_I���W�����2"���QgA��x���r:��
w#Z��KR����C��2�H���A^��k5^T�_�"R0��~9��(.�NEOk��#�WT�M �i�WtHk�t:&C(}w�D�
Ⲻ'�O�д�rĽ~���b�t$X3т����8���>8��˝���%���d���7�O���{�^���R٭�)EKQ��_E�@Y:-�	��:T{�^]��`�#g��[E�� *CV��)U3�!p`6:x�������n���r���j�78�$�~���3�f\�"��1f�� ��C�ٍ���	Y�y1ZM���&j" ���Rk�^-5f��XLH6Bt�(���ɩ-hǞ��oQ"{�z[��[�r�2s�mFiagL2�Ou��ʝ���L ,������Spŕ\�.r8���L�k��W	eomQ���"ˆ]��_��}c��~0������ro�C�,�y�p������d<�A��DW̛�BV�W�L���Z^,�r}$�����=�8R4߹~�W޶�G��S�gɘ h_��u���ǎC"��vO*�k?��{r�{{4p�l~t5�^� ����^fà�	9
���g������l�O��5����9��
��yG
�#�<��RM�ظ<&{ϲ�"�)�U'�O3x����R������'�:��ÿJwJԭ-�_U0�i��2��x���A��\���D2���w�&ٲ/V��E/�W�[�Y����d�'�rm�v��J������ԩ�d���d��]13��7[�x4)��4�ȟ�@����ǖ�v�M[�ҫLJ��6I)�%��L}=���O�ٕ�b7��9B1�����Dͩ�V%2N+�ĉu��~r�)�d7�5bA)6�[��+!�aˠs�(o���g���'��+�G�{7�.[��o^UӚ����t�=
��<�tn5��Q}��h�t�E�~� ���0����%ìgds�@���<+�˭���@�z>��>�9EGs����.f �NzS�!�UrKG"�R����1��(�"1"s���
�2�0d�d��ٜ�ZlHF���� ��e!xB�|�\�5E��j���Q܂@���Ev� �.������s�����I��s��$�.�����&y�ǽ������=~�4Q�S�N2O���N�g���u�v��_ ���o���F<��e�b�+���7@P�\�Z	@�=��K`e�QĺNQ���L����9;5)���ԪClr5�}T�߮�}|:伟jA�q��cȋ�����8�}�_N/�����rv�����*�˨l�2�����0�h[��ꄜ8/��a�=]�apE�^T75/�tƎ[��5I^l�y��S*�F��;�cc>�������ߨ�Q]��v��xaF���i�5��FI�M娙����j���U�+�0ׯg�aFx*�k	Hw +�	�9��q�P�����6���Փ��S�kt?����o�$����r�Q�R���p ��|����R�k]ҼM�����%�@4&�^xt���]-�o�7P�0��"�	�V��덵-D6)�팺��%|G˥	qh	�s3�V{
��h�JX��� ���خ!Ȕ����A�'��9�y��M�,I��BHe�Xz ��B��9�^��N��юcܢWCUwo>��]C����k�����y��Fi�yv]�A��ˏg�؆��iz� 	���ִ��R4�V�H�W�a ���q���-0���7��V�$C�%oYDN����R,|�|��dԾ�h��1�a��,ܳ�k����xH��M�1��|!���
�pP]�����f���mO�%�?�<��XĖ�q���u�p� �D�v&��\�)�b �И+Ѩ{�#%>DK
k.��7<@�U;�'��/�3'_�4J���N_���u�(f/k�u��wB�Te �v���;-���m���<WBrR��_q1�� X���0u�]X�`�v�ꉍ�2A��F��-Z__ED �R]��M���@u�ȇ��<T���%�X��kf��]X�>�55�Q@b��F�G�~[0ĩJ1^�	v�����'?}���A�7�z1c���]b8n75�J>�yM�O&;��\�F�Gu=�\z�J�f���Y�:�ZM(�}�<>V2��'j2�"��$}ւ��a��{����q˱��z~|@4�Xgٓ��3d��)X@'��B�� W����L�z�{�aD!��#Xwr��+�@�����X�	��+������.�<�]�q@&/D��HXe���Z`?2<�j�	��>7�.70��+O����w'�%��غ��`h� �,�ˮD�"�/:�X<EtJ�4XyV� �0�@4�.���3f��[1�%s{7�WCX��gR0مW�6��[ƍyx��\�����	HD�8g�h��l�c�M�2mӞ8�>V�q#�� `5�&���
�N�#2,�(����L3�fc��&�,��l�9F�D��9g�-�x՝W��~ ���OP!�yuG����G������<X��5kݎ��A@5d:A������IN�ˤ19�����P39k�GZW~{�c���n��淭����\�3G�Җ�f�&m,OŭM>
����Q�|�؟ut�R3�51 ,cG�N	���G@P<}���$�6,1
$�}�y��BH�4��wY֋� ַ�+@�v��:��&b�6mk����u%��
o�*=?Rm������P��tLr)JZ�|TW� M��`�Q�	6���ZDq�̶<���Ftjp<C�����xK�qØ�=US!�N��*��y�Ѓ��_���I��^�&d���:��a�;Z�P pף!���@����|&��� ���0�Z����������7������pH'}�l�`��/"��4�������������˩��^?*��(ܨ�q�BM��c�ܥ��7 �8�m��M^#�$ �)�/R�`�\�+Ĺ����^~d.�:�kDQ�Ag/�'�	�����;D�E[V�?���Ķ��u��"�+���8�����O>��������tk� L��,��/�!� ���r*��1���a���]��8KF**E� �U��B^bf1 ��W;d�pߟ�s�\��2�~o)#O���!���m��B(��^��N@L��Bx�jC�ㅵ�XYE�ӈ/B٭E�w�8���C�V��%�#�vR��j_�#.��52��䮠��i����rt�1�����STzs(^�C�J�Ķ����E�t�$ItZ�ǁ��6HW�G��w&�Ʋĵ�!u ��V^��3�?ƙ�׾��[:����EUWS��(�ڇ�k���ԓȋD䲡�S.XICb���j[ܧ{O�-�ď��h6�6�"�T�M��i"V�� ���l�l7V�_`
���h�gi{����p|hɘ���,��U���:��vg�P"��N��E����m�-�4���&q>Z�p���p�4`$�ȷ��P����z�j�!`?�@&-�yz�'q��+&Ym4�L�er-p��qH<�}C�r_���p6/��,2���
y�!��azM��j4%}s"�����띔��u��^W�2��Lݶ���U*�y�?S蘑�O��2�@��'m��,%��䗺g~,�Ԉ�s�_G��Z>Y:R�*����@��?��ȯX`@��b���yh3l����S)0�$PP�5�&���ΩI�2���r���y�P�!�˳�Wy�O�[
�o^�!e'�b���,
���1�HL%�	[uH�ufh��S�|IR}{6�������9�u|(%�������!u=���O҂z�2�32n����Qp��G �	�'�Ξ�* "��-�\���n�T�����h��?���%���I��ڥ�Mm����~FK.a9�I�'��W���EP+�m�ᾖ7 (>%7�f]I��ގ�u�!X���� 1��U}��A��nO��-�g0g�������y� "���򭗛�q��7Mt��M��+\���f��,�?n<��0����;!-!/�6y����:�Z�zb��m��y�P����.������Y&���Q�"s�O����㡙h?xP�o�fC����J���^2��p4;�5
���mX^(����"_A�y�d�#�Łh��IZ���ɐ}/g��v�YS?��m~Rq�ѴX
���w�P��i	�FT���b[l�&0C�%��d�����yhX��������ͤ
��-�d�{�ZZƌl\�w�?4XwȔW�Z{附�Z���3��.��t�П�������xt�>0��V��pχ��ϻQt�On�Oj���r@�e%��!�''�Щ���ƌ����3N��F/�Cȍ�v��dU���� rsD:-W9�=�c7T�*$zG�Jl�+�y�Z��PX���g��{e3�F|c#��0���©�ly�z����e,I��ro�PXש���ұ+j�e�9:�c:��b	��g����-���*�#�����������TW����{���v�pQ[� ��%;㚐��6�D�o#pwt���B\�;(׵�B���VO�f������x��W�ҍ�6�RSm���m)��spHT�]�h�41���`/'���v�������M����'�e��A��5�г��+8��79tp�С�ʅ�*Atm�/�|��^��7�V����x�� @��5�k��5P��x�f��`�@��1
��}|�4�;oMd�Wth��vQ*�Yö�Q[�|nm�t��\�'[g��|h�JRL���ݩ�v9x}4n�^���6�2�_W�i�-��a�#���1O���'�����`v�`�,Q�"\�~	)�]t�R�^%P`��4�La"� T�0�m�v�/q�P�}���i�.��
��d���<=^g�=���<��KPlTh�cn��qF?��I{�by��/��>�d�B����-�p. ��xu[�l��� v���,~L%O���WA��B&4�:�>�("��V�/��׹<X�����1v�	bϟ����XCe���O��~���q�򌇘Ծ��1�W��~����U��k�r�
*K��w��B��2��ud�;7�g��3���z*l��7�i� (A"<���ǔ��^I�V�Kd1��U�SQK☁��(DGqă_�%�W��D���*z����f�s��!�I��y�	d���������]�@	n
�٤�< �d������m��"�\���v�M�.p7+z�wo���C�#�	*e�}0���-�h�Hk���U2���.+��=��"f:�{n����C�iKL[µ�Es�����	�a�:��m.m��C���i\�N�������@O7h&��H�)�v����e��(�2+�@^l�.BA:���R�:�*�C��v�p,�u�)������^Bb�6�va�����j��4GS��ao%�� 7|��$���?c���@Pm_,�r�Z�E�"����i���W��Qx�'u:��z�#���~�󗣕���t�,I��|X�{�e��T�y�(�f��8'欅I�b�h�,�;��V͡����p��]�'c�����3	���RtC�1�^���qO=[�qG. |��}a�c����,D+�׎6J�p�OĞ���q9�sJ�{��z�&k����,#_��*F�w���E�ft�����U��Y��a�~�TN���"F]D;���p�p���Q�=?hw�X�i�Y 셻�p,���:qᎊd�����>�f��J�mc~0��]nIS8/�?�cˈFC�J�V_%�.лa�y��T��D�?��v���4\M��Ѽ��,��tOd&$q�<���[5uș�z*��y��c)d�T'	�D|mً6��'�(}����FѼB4X�Ƥ�n�[�3��ᨊt�y���*���C���=F�@N�PU��9�%J��I�v'I��BبF8�oJ"K8yc�֠N���hH���N�v�^2�$h׍��ZȊw����I�����X���W�/��P��`��o�O�u��&}8l(������M�a�t�򷘓���rx�-����0�Hb�1r4���m�O��{����Vp�xE#v7����	@�ۺ5�Cy�^������2���J�9��z�t��?��!��13j���0���䅢�8&�R�+�a�D�hA�2����|oC�gM�d�/g�i��E-�)5��	T��<��B��>�Э�L�I����zF7�ȷԷp�${(�^�r�h�i�m�@@f�	Q�$A7�R(Ii��Ϋ�b���-IE�cV��ԣz��<a��s=A���qnH��
�!Q�N����ql|�.S�IQ߈U���à�I?0���P� �F[悆]_s�֌��P���.�e�ު6����U�`r�'&��Dt����H�q�zY8r���Z'ؤz���}T��G�
�N���X����I�K���Q>�[>���b��Z����'��f(r���Y����g�@|f�֘k�������Tl�.� �u\���Zx��l�}���%6�\���NV�qG;?H0Lhj(!����Q=�l/�5�}��n�-��yɼC����I����Ub��T������W~��f�l�7�%�l����}�6�� ���,T�Xk��
!���0;����e9��hG-�~*8�BW��?���`����m�A�>R�<�	�EYC79/1O@��ӴRY<� �\�Ϣ�BA�r�c��8s�>��lH5��_�}+���(7�;��M�)rtQ��0X\n���ؠ�\��٬f�R)#�S4;U���o+���1'L�WS��G�aE]���Вd7�P�-W�xn�D`�mmp�S����~U�#��z} #�-w��R��->��,��~�����e��3�Q�<��z@BK�j�QX�&�QY��n*b�d�c�����l���UhY�=x�m���䳣p�HZ����Ҋs��հ�݌W�:"Q���^��$�;tҞ<���@MǕ�iG���}U�ZN����9�3�^^�ʵET�����i��b��O��@؆�]�!���*��S>�$e�=��ǅVR���g�D?��s!<?�6�GEF� R��1*i���N�`�z%�m���H]K�*bEwX���,P;몯v�ϙ\C�Iaٺ��-��w�E�X/h�]�)��<=W�$���Fo�_�]V0E���FP�'V+�OZ��L��ES^�̋�)V��	�4�Ң�Ӻu1���f�q��[b���n;<��I\�:K�	jt!��cJ~ӵ�zF܏��B뭛�#Ec���A�WּI���0;	��n&]T[^��tY�(.���=y�U��,�a�fO,2�g&�M����qc�r6E~`KZ��X��B���g�k/#�0�N,����Q���A+�w�s����	�B/6��G��6���+� ���4[
�sڼg�@u��C|Z��u�}ͽ`��5�J���Kz�>8��1ҏ6-U�b\�ȵK1�,	�~�A�+��L��:W�ro0�G�������M���)'�z���f�۞<����E\Tc׻�;!q���2�+;�~�P�u�HR�s���'[����ܳ�cw,ϰ��j�)f&������s��%��XKc�J�X*���e,�P��K8m���a�@I��X
1l��N�7����߇G��Eq��J�'T���6�i�AO�!��~����8�o`I`���,~�_�u�b7�a��Q˫��r\�/Vo��E�Ө=`Wu�b�B{sfj��+�&ē�X�dq�������^�#l4?F�͞�����tǷ|o	�B`9�iQ���KK�h9e��>��q�O%�4����r�v�.�v3�G���`C��ykj�.�i�MsM�V*�:����I0�6>~$:GhZ��c`�O�X�~�=��h"^i�[��H�D�F�� ��$�<~�X�a��	^}⧝��3w{�����������5	������n�߸]ض�[3� wlH��b�q=���%X8��D�9�5ٷ�)����D9'ci�1¬��-�o�"�k����V��B����L��I�;�.!�h�2�a��S�ԲƱ��F�%z0���~1]���+��Q&��:f��=�d���,}Z�t�#�d{����֖�+Oz��d�ˤN�)l��j�h@��&-�d^��C���Cb�$4����|﹊f�w&�q��Fh����M��r�O}aD��~�𖛁��4�O�o��Z3�:�<�䰘%��[z�D��p��D���뇦U�����3�i��|��T����2�3E,�����ۧG�M�ђ�^'���ɸ��Z(�t���>9��Ȩݍ"��%r/��3�"�����t��Q?{z�f��,�Y!%�Er�w���n'�'6Qe���@��{nyL��@��{3����I�2�z����^rP�䏙�oUR�}*����irU+�ED��.�\��1�Yg�6��G\�(-��
&a e����}䡹&2Ƅ(q��9��6'l�
(Ǆ���d�b jL��8��0�=+iso��H��Q��y����ӜՑ��<t�Ti媖b��?���=��В�_�{c�.oު@H�p?p�ė칩�A�j�J�>�����^�N�U�n��wI�z�9y,���FKIap��2��^���3�]�_uq��<��c8�z��Z!Pbk`4	3��YNQ5�|q�/{ؽ$�3��|u�'^��=��z0�#����5Sזؘ�4-������#!h��#�~��Oa���Ȟ1<�݄�����ă~!*���2$`,h$�Kq��0*�7f��[~�ϙ_/�+=ljJ�"=��+&5��Nʳ`�u
)!��\̴���W�U2�ۡH�[��g��M���+�;�����'S2�+T��I��ׅST&��+U�&�wgh(��㌡�?����ʽ���;h�
�[7�>	XR��[Fc/l�1�b�$P�g�{�,�ԫ����$5��)�����k��>V޸&lPc�Ч��Hb����ة�pE[E�)2���3�?��:w73_�f��kg�m����<)�HsQ���V�+n/}ꂢ�	��}���H�>�;�"�V1o�)�E��Q�v$�J�\a�g�b� ����s�^ �i �g\��D�h��b��|W;�`���(�w+M���%'��5���Q���aj�W6EL�`͛N����7V���	K�o�*P����]2�Wj6'��*\�'�k,��k��~m0���0��np�Kd!�͢+ك۱P�����s��)���Ƹ�5	*y�n�ͅ�0�R�srEe:�x�gr���@M-��͋�zhGdC��@Z{
�T�x�Zw��ff0�؀�̘���Wk��qYÚ��J�F�:7Nf��uU��3���:ɬr?�$Z��X�x�r�xu�F"����q�S8 Ub�ӐO�V�y�f��0��Ȣpa?��\�\���
��OJ�s���d	q��T`��܁����)�B"K�ջd���o����:���h ���V\�L���$���A���nce�&$<��)�_�� ,�ey� �g{��>Bd��C�;�k��G��]��lփ���R��2��gDJ��M0��Sq�"�hg��ĵC>��.ځ�َB�U)1C��`���Z����5�N��z"��hg8A��<(f���+P�-x�Iξt����sP����1�C�J��2%]��e�P�_P��[^K�n_�ppq��+0���tmX�_��O�>�c
g�e�� $���;�`����2$�m�Q4�v�i��ybJ�nN�%=���"��*�ģ�u�@�ĄҎ6T��yA��t������@��8k[y��ܩؠ���?/��I>7�׋Ǹ�VyuL���V�Q��ij@n�C�[��r���;��gA�=B1X|@J��󳦍�T�R̪ 6�U$������ �X��ږy��|�������.�.2�SMet���M�+p�}�Aٍ��xB������N]�W(�-�䒨����j+�� c7}�����o�����m_���9Z�	�bX�P�6��p�H~ߎE��G�3��A�.�s���h+�z�̷6�4ާ��K�,�L��:N1��e��L�`s����\o�l*8z��xÀ���ig����j��Z��Q���݂&�7��XغL��8�6��E��=����ib�q�V�H����<�3X�Yۉ�����<K��;E���:vqF7'���"R�VQ�NA���C�V��Ś}��aK�	p.����т }�w\����}�@02��OJo7t�9���W�,{	 BvoTΌ�����o�H�m�l�A礀O���#6M�� ��!����g�p��C������/�	�b��Hq2YB��0�S�ij0D� �P��[���F�2��`�׾)���EaBM�<PH(P+���7X��,j�tT.�h���i�҅x"ev��v�M���s#�X�q����_W�uX^��*n�&b9���}S�tV��.���w���4߉�q�]��3W|jE���;�OI�^�A�X�0�.KP&i���s5ni/0k�о��,��3�vUo�NT�ȋz�����"�\�i�m�ITm#�+�{�Zd�v,v����	8�>��\[�H��"i/j��bc
/B��Y
Ԣ6�F'N�����b�ӝG��8�L���4�e��ߪ�0m[N��3<���9-��T<5���FR\����I��g}Vsu{q�BnA/H�m�Ú����e����%��ͱ�?֑;�N��l���w_�J�g4�^�� S�]���-��c�v�D��|B����3q6QR��=���ϼb�����`�� 17�n�BkئÉ�@�	���E���A�0�+w�bl�"/m��w�Y��qY�������o�Ψ �.�L���-���`�zȫ����K�Y��8J����FxY��W-ٍI?S�Zbl�'O���H�*!ݫa˥w#8���ͺ�zI>P��q�?��m��v�'�>��݂W����D3���-,\� &a��[,S7��Z�dI�v���qdP��j<��G"$���5�[�Ŵ��PC'˥^q�;���%v��3�y��j�
�/	����51)Q'��((���F#,�!$�q���B�e��+����Z�U�)���,�����cX���*ks�)�%�㟃[=4�v����O�O֦�������2�h�'7�9�}]�ֺ%� [cu�V�'��a!o�S'�Ԯ��Q=zP.A��J��U��N���՝�K}Nz��` ��[cmMv�)�t�ڞG��߿�E�f7$1�IQ�0����ƾh�@%H���]��Wn{"n֗T�!6K;�����G9+^��f�qWaD���5����Գ����
��X�F����� 4ĝ�'M�G����^��\�.����Q�o�r�{ɥ�$�Vj|��&}��=�B��\�	�����b*+�~���fM����]D��ym{���RB���(}��4w�nu*���*�����ܓ�:�U,_MǠ$+�j�� Kkf�x����(���rq`��h��֏��h4��]��84)���|=Z	���h-�J�.�X��ܳ�n�ۢ��?�pY:j��bG�S�e �X�����}����z���'wC�%W��'ʏ6C��p���P�
�-��a� 8� ��`E�JE�:�d��^��A_uw�V0���|�" Y�!<�� �F��\�U� �,�o����O���fC������t� B�F��:�/]���4N��y�q2{�3��q��nG�v8�V���`�^8N�y���I:@��ʆ�Dî ~�	�%���x���� ��Ǐ�hQ�df	�}���D��<F}�b�a���dk��NR�7�m�!�`W!�{K5aD��Q�,��J��]O����Y�Z��:�"i����y6t���L��y�.�RmV��&z�}�G(�? �Z��l�$�`U%T�!����]P�TNެ2���(�F��<)���� �3~g�X�+�zS��Qdת�SSDuBɪ��(ᤗ'���j����&yC�DhP-�.U� ;Bh첃>�b�R��¢�@�q�P��#l����\y7���;#�뿳��躥^V�yu����b7R�C�����r��|�P �D|�˟Z�{��D�6 ͌��������Ʒ5^�p&��Wc����B6�<Br�D���^�8�s��V-j)[s6���,.X\<�O�c��,\�.,~!-����l\B2�}�!T��t�W�Qǃ\b`)�f�ڠ>L�*�ڥ6��[r�xvr��ec��g�C���.�e��>���=����3cJ��2�1-A��[AUE�YwS�6�~��6/�/��\c �E5�� <�;^l���e��ͨ�e��fcv���NGY�
B)BP��.�ӂ<��h��}NCӤ�q
�D����I.R�@�N�
�0�	�����s y&%�*��W�0��K��Ѝ݆ �.~��j�ޠ�V9��YH��Z�6�Ph��-�qCK^�����V���� ��?g��ϊ*y.V2l�[��0���!�@���ܫt�r��.�i��ծ�kAR8��5��jM��nH�p�~� I�э��1�J��ڂG$J���aN�ų��r����~r1[Q~�"̿�<��ِ�eu,$�ɊWې�>���7�q}�S+����\�d�RFIcE���T0f�+9z"�fT�ZX�)�Ĺ��*2W��/�	L�D����"��pNT��7^���?1l��x�."�e~��eMv����ntn�̮���2�?gU_��V �*N�H����tcv������~�>���p��Z��x�n��߽���3���W�^��r���������<LaH���k��$��]����������0(tQZ�@�	�-�P��͎��Ç�ˢ��x��̵:A��~9)��/�J��M�Z�'��ҙ9Qڤ�as�Ä =���8T��=���K���� �V/�����*:2��4"��l�`�z����?�뉩�ԣ�q�&*�WX�����$�v7�����p+[��=.#�RS1���wx����_�6gٓ�
�n�駍]�#pm2,rz�Y�+љVx�dMb���1�A�m��J���ZYN[
�p)�������o�N(-�v5�w!�^7���&�B%�з��"+<���5�p؝�Mp9�V7�E'�����s1|���$m]�$�����9Bl�����
�Y�'��1�d�	�3ToŐx�,���Eh�^J�KsI�e$C��A(�7Z?�é�|����s�w��wpy'a��;bԠJVI�{�����$Z��	a[��m��	+�Z_��g����Z	����Tnp�A7:�7�p���ŗj�µ΍�G�T?��U�������Ǫ�o�������0����%�6:r>8@�/˒U����RH���{�(�y%�� �K#�M27����;*C�rg��̰Hfa�z�T��+H$R���Ae��R�-t��?���Od��s�,�=��ir�܄\���B)ϻ&Q�{�ϵ��u�f�
��/�N�,(�Mލ���,!�2@f���h�08�՟�"����D88�vr�B���SJ��)7==����B����W=�D_��z����>$�'iD��5B��w�����H|@��|0�:��%ObV
ߠF��Y�b4�]��*�PZ���7��2^AyG�%��*�4���R��h>^�;h�k`Tx�Z�A��
q���,Q�����E��`���Y��]v�p���v} R�г����#=�м�vBYM�,W!��kw+����j���=��G���p���ᗕ��	`�(��Aǃw�w�K��cW�����3O���%�%8�������D�E�
u����4i���pH�����#�����-��,.y��g�$���iAh:N`���L�����
�oy�KvKw�9�Ɛml{�a�'v��,`�X^B��U�ln~\�f��"CW�n+�*�1�_��J�{��G�.?W�HH}��a��׉���sF_�0��\�<�cwgS̿�8���U��2���� df)�6EX5d���\F��D�� 	��4���`?kQG����$5�i�NE�	��[�Nl9	��p�e��+0߲����X�!KZ/"��H���*y�2o��Ѭ��C���ۗV@�;°��	]/�A�x�N�ۮ�}���Z��n�p|R ǂҕ/�P�b
ƑaL*e��]�Q��Cg�D�f��i&`/U�N��_"t���x��i���S��{N7��Xz=+��ݶp�B�Ƣ�=��"�t�����pXg^�.x� ��V���6 Jh�.#�-	��ɞG6�*v�H �@�(Lݮ�ؾ��p��j�_�ͳ�#�U&��:�S4A��6�y)]�.��ZƞI}?0��qW3�����4b��MO�xS'"U������$��5h�Z���A �q����[$�q�O�PW9G	I����z��7�)�^Q-���h������%V�跆N)hy�n�tt�%�V�̒������d�~�5�����������d.��f�{�9FC,d]��3T��O*�y'n�~݁���d���a@}�H�=̒�M�����)X��~ҺHr�45
����*��)uFR~�o�P6�q،��_0S4�^���n0ȳ��g�"�h`F6�R�g����د��`P0͛�%x�-����l��W:����?\����M-�a�*(nN�!����<��Lp$]+�&J�(*�Ӛ	�e4�T+h.���3�Hj�?�
1�Yn���� �}�K�E#d+�m��2��oR�g����i�Yo	�?���ȭ�gebfd|6�Sbt�����K���w\�D�aψN X�CNȔ2"> ���~0��8� ��͜n�5���'˦掻��
}��	ޤ�M��gA�0��z�^��;��rb�z�w�i�b����&K3f)�6�'JX���gE��Bc_T��҆GЫ�3.�{�9@o�52���?�/�6bM�1wΒ�
X�g��L�`�����ӣ+��=1)���΁`ZK�]ɨ��UuoZ����!�6��t��bV�o�40���CjC���;\ ��� �ɇy����Xo�֮'�����1{�s�	�=�
�:��1Sd�m�cӤ86��Q�^�齁sB�d�M�G�W����P�&��ޗ�� ��m�)��Ӫc�x?!9v�
��Q�U㙖c=�B��;�^��#))X��u�,�c�k1� ��qD���o!���/�n�oQ��?<���h�'�R�̵6���F-%���z���wo�MztC,BYBEce���ۄ1*�5��u�b$��6BdIn	�t�Q�ѷC���h��rm0W��F�sW��P&��3E��~`Եe:-~2�ن���xk��{Q�S�F�g�k<�	���t$�ج0uVX�����<�$��ܤP*����0��S�B P Q\��H��z�N��5�DtK_@�28��#e� /��`�L�;��6�U����I�S㥚��T�~ۚ�iu,Pp�P��#�S<\.�hH�������e@�؄:�t�O�I���H�m�q����z���k���TtAтW�ea���x���5L�U�q��2�������\,���K,y�vv�.������ΌvY���|N��.HE�p��}	�,=�oѸ�?G�n躤&cV��?ݪ4���!O��	?%��J�Q_��Z���9ܢ��d��
bd�3�^=m�fev~T �Pn���g����%������*�����W�je[�>�~<���(^�k�{�>O�1���Љ�*b}�Kb��\��IVvOt��S7B�Ͱ�d=}2j�G�?��i��(�3#��OVDd�b\���<t��\���E�9 J���
3v��ۣPW�g���	��R��%���0�2A�>���P-ӎ�u:o��\�PK�]�ֿ��I�RM�
�����r��2�ˈ3nC�W�UY�Ш;*�����4�o G%ߵѠkװ?�(0}����I�w-�r{�?	m�A���ǀ�Q�,5��e�]�S:�`c����E�ж��L��!��SN�jH�����L��Wn��]V�ZW�RF��)��ӟ���8�i�ؖ"����anG��J��x�����r��o�/94�a�nx��`��dJ	�e��>�1ƣ�a����/��� U�i�hH-_����(�Ƣ�y^��=}L��>I��'���ǌ�x\�"�U�4�A_D#A���9���6z�����	99E| [=��6�]�pp�=e'�(���;)o�D�8/
DY��>�f�{����j����k��vW�b���͍<�/c�]�k��e!�u��e�´j�P Iwa�2�󫳚�s�ȝ���Q��>�/h���<��s��|R�Vϡ�V��ǉ�WU�u��&�'oG��#�_�i+L��wn����W��1p���?�E����!���nM��9�A�S��i��E�����]I7R�bݥZ7@0$a�f���%I`ҫ]7�%]�+��v�~n�N�)V���,�������>����A"��^6�7�ĿBՕ<fel���͇*���f��0�[�8rN8BKO���9瘇������3qc�F�FH&��i��W�I�gI;���9��z���w±	},(�g	�E�wQYšj�3�{�V(�òǒ4��k��fKϊS���i���W��e.R�PC&����Y��xrH)�\��DZ��2]�H�fє�9�@�D����,�֙!}ѩh��1��²D�����O��4Q=�)ƻ�q~W��V�_-RƯ�v�ҳm���2�W��<���0[�
n�bYS��5q>��pkJ�'�{O��ޘ@��رI�82񉞖���Y��OI��!熐J��x[���n8����63�	]L���������z����P���,"�]�`}��� �r��P\����2���;V��;F�:ޞϾ"��q�f䟵��@! yә�MO���3�+�u��y�����Q�{i{��~�Z� }��!�� �&�eX������[�y��;㓤�E�g(��}��Y-�34��\����w�w5��x����5�)w��I�0�I�j�%�@w" Ѳ0�BDp��%�h:W{[�h�o�3:�c��L��Pp�%~������b"�\��$��aC̓;G�.(�#�R�?��#Y�u�d>�-"��"VD����cعJ��0ԍ*���%?%{��3�x�1�Al�h"d�a/D"W��Z{R�$��!�w��'���wZ;Pɧ�N�Xـ�����y�}��N�C�!�t�H;����K��%�Ӥ�as}s��/1��r2s�R����R��{�Vہc$��*#@O����T��Z�7��p�+� �V<t��>��M�?�3p@�c�4�-8S �9�r�x��=Z�<�]����i=��7���㠬�à�۽%W�>��|���q��bP7�v�A�풉G�@F�x����by��p	cj����!Եy�����3�[o�)!��K�9u�3yҍ�N�f�H�$;��D�F#fY�:�� *K�'�h������W��5����6�W<C�z`�e�>��bȔ�g�w�rc�I��Z�iz�޹�(���ƪ�y�����Do��jq�W>ǖ��{9@�g��\ۦ8�3P��2h�7}����i�A�@��03��|��`3%?Td��	�dmF��@Otp�P�qc����g�Q"w e��L��.h��tO!�����u��d��s���L%��Z�"��E�D��}ҷ�X�l{�뻹�1�6�R����ZKG7c@>B�[z�
z)�`;��s�%�S.��B�%ď?�ש�r	�����g:��w�#�,a�;R��4�i���v�=c=���>��{�h|�vг~c��ǑZ�]�ME'�XuW������B�i�a�!	�G�Y�ȝ#6.@��底H	�!��wl��8�Exd�o|��]H :�:�s7��P��R�"�-bɷ{�E#sW��|���z�2���l��#�7ch�=@�3h�1[����ǁ�-X��.77i�z f3��ٓF�A)U_�DM����d.y��Do:׵�K����1V|�x�/��⪃�7�$z��PeI�T������,�V�.$�+�`�cg-&�[��1L���U�e ���k��:eH�+�v\qD�e�h�QD�uH��y��._���5��'�����z�6�1��C��������N#�E�]>q���J�vq��m���p���T�.A��6q-g�W'�=�̗��x���S4fsB�P���X���n� ����T�n�ܣ��?�;�q�-��=�P�f*˴D8�Bj�KQ�0�:~�`U��ɼ�)ά0ϥM��U�>�A�es,�#˿A%�|�6%] O�0�Ą�i�l�R�(^|g� �iXzPOUtjD�Ӟ�}%��V��"��.���Y���2pE)�z�V�k�h;�W�Y2�����SG7�Kv���_�F�F�����p�/�/����/����ҟ1�5�-�K����1o/��1��\�z���d
[�Jn�ʋ������"���z�(j�zsZ�Q�:2�}F�YN�c��v�ῴ��ı�_m���tLy�QlE�̒(��hb��|wv���ӆ��v�8�6�F�<޸��K�4.�v{��$�t����E�Xꜩ�%�se�L�p�H�.�g7�f{9���]��tpc��&�LӨ�,8�Y�6u�B�k�� � ��R&�l�6����Cz�Bv�u�3pu\ĵ F��� �S�X�K�$}�f��.�8���B���%��m�S��'���ۃ�a�F�������"à��gc�2'�r~+�����q"�0VJ��8#��~(ИT]TW�yK�k�+T��x�*3 
nO�}R����Skd��視�IP��1����|����/�������d�`Xd��[Q3���܂V������@0��N�sP	�On'��8��>\�G�8���4;$��JS`�w���c�҆ğ�F��{�.K�	�[T�$^'�ҝC�N�w �����gp�u��3���-3�^�K��ۖ���u�����7Ǫ��1X���>G�,X�x�m{�Gp��
q��qK��_0+���a

�r�+����tG�U}�(��;cً�g��TX��W����6���EE����d���]Li�q���Il���Vm�Yފ�S9P9d���Da����i/�q���d����q�R�4o?����\��6aY�����;峫T�}4�,�^�C)�ͨD�U��y�Yh��bٗ��ҟ��z!�O��G��<�R���OF仦����6ed���d� Z�(/
���ؖo�}��������Zh*ףe��/�'�v��5�Ѓ��6�⧲K�ʋ�xT����X�p����>�y�d-7&�o36h} �ʔ��D��S �/�ǈ���8Щ������(��^���NUG��}4� R�N6�f��{؍�vLA��Y���2;�@��ߠ�K�p��� �p̚7��!�W�a��	�ѹZ\��m�]84��/��>�/�p��2s��1SǕ�!��6��>w��9mCI�V�~��g�<���j�[r�)���'��co�{��u������b����I���9��~u[��y�'�A/��������[�;3�N�(���bEQ]�y����mp��P(?&͎�3͜��?�]>�q俥�*�����sj�=�b��0�����tg���"[n�n�f :�W"ҹr�vԛ]����`��Kv�f���U�A��<�p,�XE;���j�N�oAcF�@�/�'�����@�:k�Ƃ���\=!0\�:�J�l���>RrJ��uFe;E�8r�q�����)��w��"�	3��@Q�ņ �'�x�8�����8������#�.H ����Z�1ȸN�0��`J�v/�{ꮴ��e��V��JQ�Q4�)S��N�]��}�7�V}B��XԾ}��Y�c��(�1����8�,����6���U>���e��5VCQ��<��݃�S�e��PGS�3��C}B�����8���+&�)�F�`������Ud<z���Ѕ��cT�qG������;��K#�#W��Uy!�� �3��n��)� I���JV�4S쳏q�~v!���#-μ�)��ezh�8���v��\�(���c��[i�)�L>�r�/]<��T��tV"l��Z��_u�G [�R�%B�.�'<x?^��CD�?9�n�d]Q�`۫�UՓ��r ������<}������G�s�N2��0;�p���nL�^Bs�[���9��йt8Fz����c�`�������s�!�{D�J��7�]�� ^�sA`1off~n��]R��9Al�f ��bg�3��/��7ԈR'�:�(#F������KژÂо��t�Q�	A^��~=t��C;�|0���Y���z_#�Suu5��A���/Rn�����{u"Q7kr?ۀ6*:��.3�:�����Q�ң8*bs��ra��"ʸ��|>?�q���a�i�����{6��i�s�ks����&�V>�Q�A<����M��G���
ѺfS&U���}�	 ��}�����
2({�����f>oyV��ɨU%!��v ������'��\<�i�Xo/���I���F �0���=)��|��&�Ɨ|�i
��IM���|6�k)�o"V��aG���S�ӣM����W�Y}V����8X��`�=B����W����%%�Uu��?�� ����V�`�9���!+3Oy��~���t��h���Vᗇ��̠ݍ%я�NeM��+-=�t�����["@F5U4��&�V56�U�l�C�"ǆ�
�A6t���T�ѳh��v����SW��`Z��}f��a�lL�����ƶ,�$�G�m$tm���[?�E6�rP�Q7�U�BjF�9��{Ҵ�3c@�a��F�!��Ų�P�c���:�_<��4Mk���S3�z����z�����Cƕ���G�P�-�3���|�)Ǣ�!.��I^0�i���w�5�0\z~.��=4��+Pq��� �e}_a�A�xWx����37����RJ�lu�1i|��hPs�@����Cn0<���ۄ��3-\�gU���P��J�t���l����n ��m�O�����+�a���Ć�^f3�BO�g�{ȩ!gE������T(�c��_(5�P�ywJ2�Q�X�t��T�b���՘��6��/:'=�z3<�#�=�nb�Kp����r�7~���K<%y>�.�Xl7����a�/äx{
����J��6t���4��t�j[�����kW�����O�����@�f�C麚��ԎU��H��=���g`^��J�����[^��/ 	���4B��LG�������	��姗�={*�50{+�6��/�@��S�d���	mp5IT3�f�<
��`�!��]����] ���^�dv��6�q���a'�^�c�	�͠4^����y�_S�t�'��A��&������ds�*E,�W�����Gک��2)�Q�Kр�)ꋁƃ����6/u��f��m8�|te��3�ڔ�qK����y�<s����m�>B;!��w`�!��,������1�(��qKw��i��n�c�A����6H9���+�W�%�af[3�(ߺy\gU������4p<���0�z`m����4����T��Q��V�#�'��u�[��t�c�r�"����E��;�:C-5�86�0�����F3C��|�{���4��.%���M�|�s�j"G�{<X�c�����՘��G����Z�5��*U|��m�8�f�:���؛�!�J�4��t ����1�dr$�-Z8��j�}cJ�`Ih��b�]��H��?�oXrG�݄ڥ����͈�fV"���ALre�$j��\��tn��B���p%�O�T^�	����L�Ę5�F��
!Xr_�2���$�g��#$�.�Z/22�\	�Fla�J���q����o3+��^�	��xf�X�"�H�xJ�N�]�����C�������k֌Мs:0l�a���&�A||ԓ)6wD�}c7~z%�����,�9����� �b9+­+�1n�R$d�8����#�c���
�Ds���6��R[NĿ�$�����a��l��;����?��V���X�F�Z݈
>GU�>�xP��*�*�A*��=���bA.<��^����9�Y &��@+�w��y4��N�Sˬf�燹C]�k
����\��;[��ۢծ��BG0�L�#
�,R<.sG����*���I��#�w���}VTIXI���x�����B[ʢ�D��8סU�y.�1�4_N����������<���_��w�
�� ������Uk~���+{`���c5(dd�"���b`ZJ��ܧ���`iI=�m�ڵ����c�MΜ=��VI$Ad�����Q%�W9�/T��0��s�=�N5�\Y-%�}w��ח����[�H�G7(|�{����Ghf:�=q	�O���� -���sg���$��:-�}������:�	0�kU���"%6�A^�:t�S�K�vM��E|c6M��
,�R>]?�*Ce71��QY��z�~���J������-��,6��Ҟ���v���	��|;P��1�I�����A��v�Rg�#
���2�(�T\�&���p�ԙ�d���Z]�c��	���L���kS^"e�CSJy��)���cT����+'���/n�B����[f�]N��h�0[�{|�IGT�p��c����o~����@���eu:R������Ash"wC�	Wݦ:;��w����R��uu���گ�0ɇ0��0��r�m���O�E_�.�:c����&(�qn��c��O"�@9�#rP�z^����1�f8�\��F9e� }y`F�)u5��j�g�"�9K���&T�6�Y��K��@�߲�[�ϊT�lKq�)A�T�H���[x˽8��]���������k#+G.�d;& s� ��y���n��PH9<��a��T��t������H58�w�4������� �(�:|���0$��ש�[�4@f�El��L?�`�l��M� u�.������
P�[�&��&x1ȁ�`	&ϨQ<�R�@�z[��}��*v�8vl��?�mk�����NՂ��@��;�pQ�"ζ� �,c�T~q|�i�F%�_xǦ�bk�����ӕ;P�觷�t",��5#���D��*L7�J�������pm%d�R�&��j6�4I�0��s�bT����d��f�\�7���
,YLgWH���v���rbR�]��^����p�q!	�#za�}�F�pZ.�Y�X���䷑��N�~`y��	(ÿ�աT��]���)[���"l+t����/ʙ?� �@��qal�K�DG��ē��&?)��I�U
%��⚋��;/T���0:���㉴��M�{���B�Q�� f��P�MF�ͥ(Msa�2�׬>����d�g+e6J&eF`��zU��	�Q<������P]z��!��ݸ��~= ;wp4����^/�K3��z��=	Z�\����% �J�����R�������J��`ߋ�>���\n��(Y�V��ik�C<;��(eX������%צꙈ'+�u���{����k�aC��dǘW\_3Ǌ�)x�f����<�~�#{u&�j�L%G�)(g���Nc�3�)���u��G���s�8D�T���l��ߺ�I�Jb���5B�����XȔr�&]^+���q���>fW���#����4E2y�h�H��߬�9�"̺�쇶i�*���8=���DR3ZCխ�'�0��G��_�H��"�o�>D^��lu�)`
?���-^2� ЛB�1�8h�E��,��8P�?}.[U�CM��=�r�`cSU�'Ɏ;��h���7�������x]F�U2m�g������˭�c1���2���P�;I2��Q��qhQ���5�Q*Ap)�$���D�����;E&�L7?PSj�1�X��{�tA�	�4�2�D��D�O�ڕ�fԬ>�#*i��I$�%?�33��%o�.-���uf�Q����I\�#����Jc=��gОn}ƺC�c���i
��#���S����p|\ ��\�E�7�t�u�����8����lH�#�!
����"�E�ө��$�D؝�}���"��`z,�����ΜW���xcg5V�M3��i7.�\�,-.c͉�矟����XΆ���^��)t�A���͔�~v4�Q�W�z�[6�R��Ͱ'�n�}NMß����妃�|��b2�/É��O`�O*z��f�X3����f>�!�bS��t2q�O�a��a̌z��]K���ω��M6�X2`�1�G������Q��M�<�P��dY�-t=8T��YK<H�[�ٷ^]/�'����r���r�{#��2|$�5�4�1!bm�]}�	��բ�8�7> \?��1E�[J����Jѭ���@׫�"-�|L�O}o�"��{��刲��3ZB\,���~-������nD���j��@Ċ�A�$a�s����'y3h߯{2f��� <	1C�E7��O�%гe/�dj��?x"�����k^�_�\�φ	kz��Yc�DU�P�v���4 k[2��}?/"Q^	�(��,B"0�a\v�������qcHN�Vٕz�yXߡ���#�+Q�J���Wp�p,O:�����4����iq�#C|W�P���5;�5ԶF����;o6�&�Sї?پ=9>��I)[�H��b�:|Ra%#�p� �EҔ�� ��C�2,}������?�z���u���6�z���;�/p����6�d��"�����8��-��_*��V��e�K3�ǽas�_n�\�����o�+�m4����%Ӓ�圄Q*:ⷌ����'��� t|�����F
h��n��;�MA���ȾH�i�ݜ�D��Kl��|� ���G��x��x��3�ey`��h����	C��ճ�m>�Lw~�	r��������� ?o�a�ț�$�-� ���
�=��(�@l|+�zɁ9Dؒ��HIS�l}b'X�؟�#�LP������{'����
�i�}���<SQ��6��� R7z�hq���e o��mT���Gi8s2k�^Bk��AV��Np�h�u�'mX��a��ٙ�����7��ţ�8��:�̤��Z[���V����A�{6Ƙ������=��>���H�^U��q�쫥(�c�1�X�~��$E`��[�H�K({��/Ou���z�3r�_��]�7/|�X���*��-Q�E݊��/����DPK��bd�6FS�%+5�#����n���{�<��M�U�����G����O��ʍK�c�>x ���C�gm
�����z�`��⿚�Q����i���Y�piśЛJ���r�,W4�u_$
9h?}&��z�,����~�t�{�&��\|�9SC�yS��ѲG�{6�����Z���8P�.���'����s�8���*�BSR{ ��m���i�-���w��OQ-Z+����6y�)���
��G���q�Ԋ�N��g��]Ohؤ֢��ywق�K_ݠ��/�[�m6��"|����=kAl�^�Ȇ�8�}��"R�MS8����A���W�4���&�:��a�0�F�8��'v:�����1�ƣ7�1�07&q51��#��]M�5u��(�~$jd�x;���lX�j�'i�����e�Q�*6�B����~`�W!J'�����/�n#Xů9,�1Q�H#"���@M� 
-7��0�դ��c}�!�I�oOn#�U/�*䷤��CJ��q�oq�&������wC<����}}���F���[<��ľRK�N�B�����u��m��h&G�X{�c���m�݈)?�8�*����gF�5��FdZ�f ~D4��	����R��<�A���P��^�s�@E��~���'�Q�:U"<�`�#�(G_.�C	(����7�o����:���3٩G��
��kDo_U���K{�y0�+*��_ ~�O��3�a��@���Oi���j�X��&3�|�Hn���n4�U�V�>��KJ���a-D�6�������?YjҬ*��M�|�������LV�i�!{��	|`:���S��LB��C������l��W�N6��Ǽ%R�#V,n�׷(}@�������V�#�U�󰨂j��B��XR�2'�OEJ�@n���+>�ӵ�q}�D��@8�2��a�Q^�s׻ .�-,�X�AK+�>G!w�C���Tp|�@��Y,W@�:�,�*��.� h`����%�(�sh�sp'���3��r8F���i�8��#��ak��sF�$�x���7�������m�Wݯ��#M�����P��!�>_�l���!\��,�p��	��$��@Gx����)���r�z2��S�e���/���ķn�䝇&����*N�^v�γ9k���a���"0�9z:�k��E�?��5�Y�U1�G�������FXt22���s�Hџ�3��o�^�Jb=&�6���,L&�þ���cy�[��E�,��]��[)!1�$E�9�����^v�|m�(H��0@�V8�;�=�8��r�(�@�pK`,���Ȗ�e{�-05ֈ�]b�B�S�Yҏ_D!����X��@����rK�3	M�~�i���8�Ǝ�:���r�z&y15�1�j��7dS��4���I�N*��Q¶U���ʵ�
���,�?[RyY'""�j:��"őaȊ%�\��h��z��$e��8��.��_
���A�U'T�^�F����R�"��GD�����:��fI�>�vGN���`�6�l>{ܽ3f:�ANQ%0�b��h��~1EE����F�a��Q��P�ς�c?��v��	Yw�8u�_83���xE%f��PH�f�ޱ��_&dP��������\���C|�i~��1����T��M�;��rIv}�on!;��I�>�`�3�c���4��5��*!|�.O��d�:
���=}�� �N���N����A�g?%9FmĒ���RjFiCS5(i�M-W��.c+�MH�"Ь(�M���n��;�QF����:���?} 09Lcu6���V����5�|Rfm��'���A�`BD�"<u��p����h��$~�OI����=x�ʹT����R������F/�<e�-���I�Ŧ�~�iق�,�n�T��ڌN�#8�g��M7�z�=(҆ȓ��>�1�\!U��4]ŐC�g�:WD������[_��z��]�es�aaJ�=A��ԍ���͇f�n'�xr<]G$3�1�.�d�2?ҳ%,>�%[>�&�jN'�FF]�=D6AD�J�C��$=��+>`�{T���&;�~����^�']�10��qVc\ՠ�ݤ�=�l�J2��I���WA� HĞ��l:/����X8�wtr1�����c�}Ӛ2�F�P�
<#�-�\QW�8�菭�(�߀��aŦ�F�gSW�K�럧���q/[���X��}��GE��Xذ��k;�妸K���ߪ:�GB�R��)}/s\]1�q�l�;���%0��?pzX<��xɔJj�?��R�$7�fg.��lr��خ���Z@�CzaKi�VC�`]勹koO�ٵиy2dQ������u�Xj�]��Zv�4c$��*����!���C���i|j����9%|�ٞ���q���]֚mau}��Q��a�>�� �T���tH�h� �֯1Mz$������O�ssI�?%�/6v�;���W�Q��u�j��}ƹd���:r�(@]�����6�W���\|gxZ�q�o,w��������B�tlsvO�pڼ.Ҫ۴>��l��Eږ<�W���a�.6<��玑ľ �)n\�;���%ӭN��Am�y�A����W�q����HQ7��1�+�?fm�\H������(��:���V���{��rQŵ�S��x�R�>����?�U6�e�:�ˆ*�8�o�=Q��R�k��r� �y�������QL� �^v���[Ѯ�}�\�;M�Vl�qƄ�~��2G�C�U�1�^�D��{���`�D�d~�C�8���Z;����ݞ{	��~J�zE�@�y�G P����9����O��3I�}�z��]?nԛu���y	���Kv�&��ӦT��zi���v����*�n�0�e�Dw��$��h����9xԞ�jзnt���{�BBR��v,i"&�mO짝x���EH7J i7���)���E��[EVnL�X�YDT=�DE3T�j�S� �ga��Mܽw�3m�����+̺�x4�`-�Lk�/�$�XH�>� y�"�:��L���G�1����y��r���H�0K�fIP���n/����d��+;�n9����|��e}޿�#���L_�A:4&J|�ݯ�=dg0)�����ߓŵB��f�k/�7ER��S�����?�~f�1��&>!0�ѓg �W�)(���� �R}Y����Pa����O�Qdi"N{`��/�!�l�_��~,�ϣ��J����ٞ>�댾�ZI~	R��7z�1Lg���u��N�$�W7q��}���
�X��M�!5������7�������9�6:	�D*�sd���� ��Go��5�W�K����_�����nf#?�U��5I#L�u��h���>��@��{�$Qݨ���f0$�YۆN�-��4���׽�����r���;T�{ɛ���vq�T�VՑ|B֛�l���<�"�5���[��L_0�,�V.f��h��b�i^	�Џ��e�7c�ޚ��٭R�َ�x��Q!�`Pj�� �GL�y,���aSK���;�Dbu/~	�4�޳������|��~�+cA���B��N�dA���Av��4e�ĬM%����+���8)A����q���o�Ym����v�J�y�߯<�g>R��^3"�)¹V�BR7pJ��Wⷥ,�l�y�����k��0��q�̂��g�1�J �����aٰ�7�6y���s�VaT�#w�P��(��]]���� ��gR�緒�F5�&"O��^�8���\�1Bv��:���N|���/�F<���H���7Fy�4}�Ne	�x@}���P�3�?�y7Xb1��l�|�C�ۏ���-���l=9�iC�)��P���($]zԫ�w5�_�].��h�":�it)M�t3�ĝhF�I��T�9�P7����
�V��ʗ��*���Ĉ��?YM����@ԛ?�O:���6�W��0��B4	]�<guY��T��ʔ~l��m����]!�*M�M���=�1B9-��� �E�/�����	��N�P�ݠ�D6���p�F0s\8��i���\�q�.�����J�J�������&~M+����� C�=�5}�l�)-��I%q��N}�M�R���F)�y��n
BW��Zr��m�J9n�{��q̩�"��x��/����6Ǚ�����]g�9@��4�� ���:���|Q�W����ϭ`X��%�`�h��*�*��2(�qª$�C��68:\�t�)��Մ(�~�6�J�/9B��� ��J������I�E���.Ȩ5���_��=�&d�%!Q=>�d9Y����#�(\O?;�񵰩!��@#P�׳8S29��a�V�1�����e�l��X2��^/<���m�a���R�D���t��}ʌ��\��>�;WJ�����eFR���H���e#ӫ����(�HRh�ڕ�<@W���蛃X�hN� p�ѓ������w��c�(�QOFB���4b4Я�!��O'��
�V��voc���R���Q\'��,b��݋_��e
��K�˅?�����,j.�a��9Բh�ڊk=I��2�@��ei�,�W���̭yv=��W�V�ڦ޻�Ƥ����ْï�%_PV��sK��\Wx���H��k���%�:e$�n�{�YW�%�s�8vëP���
�':*	ޣ��qΆ�/?.5#��?���T��9Dc��[�V-Ɇ�&�\���!�`�Ё��^W��U�(���̂y��0$3	�DhwO�+x6/�H�[\(�yc'�w"��3ɚA��|'����R����v>ہ��DLQ�ݱ��A^��B��Zx��@����j#�`�j�3������~���wAy*��r�Ҝ����ڞ<�6�y���N��})�;�v��A��e8�Zϴ��S��!�yb�a��&����(F{Y�c�Y�p�y��U���-�ܺ�O!H����<4R8�9�(�bV4�?N+H��VX�Qz��x\�(X�����y}X�4��,�Ⱦ���.Z�6�ܼ��(	?��[7a�Wi�icRͯ�©��{�^����e����pyyTC��kėI-À��dz�.K�ܚ'��m��ai0,ޅ
��Do.����	�&)+��(.i�3x�r�l��3������,cD s�U��,��4�e��qT3Y��8M��t�Te������L#�A��F'����앇����6��$e�d��v���_J9��6.��)��#�/\�.8��b�;�Ʒ��%e�6�Î�L�롁��Y���.�J�_�㤘��r�/=7G�k1��8)O˔�8��9�n;��h����>[h����l1�ZZ�"����B��Ȇ��艡�GǸ��A�*7*���L�I�<������eɚh:!�	�/�f�;=�^�u�rR��7�J��`�d&�Fu�Y���՜�ɧ���j��@����� <�s�����!��ay�>���_8���<%Z���PP,8V2��s���kQ�8�h��Ts��ΩA(�]�
��|^�,��چSS0L�9WїY}Z���ն��o��[� ��A�>I�RaЉ*���W�_�"p��,�]��ᶜ��k��,�+��O6��@�|������s1�X�	dl&o~?�ժ�^5�}�=��"zF~l�Bv{��K���{)��lY~#��x-'B��.�l#��[뉍�м�S/�����K�w���^� �G�qP�ʁ�̀�zC�¬����K�=���D��D���K�7�.]�$(�.1�
���{����w�AJ6�Y���f�=�zE&Z��i��1�0�������|~�Y@5KX���O�Z�E�ؽ	�6e_��FP�i<?���od�;^ƴ�E���}��Ca&�	���;�]�(�9V
.)7������s��%;��VlǂI�$U�r[$�	N2�G3�°!LX��v������3#2ū���*42Eֆ��1=me���.V
��X�EO��%F_��v�F7`�͡�=e¼Ai��z)]�c&jBUim��e+X$��k~^h��� �W�s����2���Ҧ��p�C��N�B�ZN9~�q,�i��Y�P��2ө�s��^����$����L���9����`�͡��|������B�֬��bϨ ��y�ayn�p�e��dn.O6�k}��d�����+'�� hJ� �Ó~�0�#�y��5Y%Ь�g�G�׍h	8�H��].���_TcT��K�0V�|2�j�����ম�d���$��|����΋���:k!:�!3�����	�s�VK����w��3���8�	
@��T�4���"G�ZՒZ��?^/�|�͆ytW]�{-�����0TT��������e��d1^��Zt���:9O�C1x��Y�aoYxq�'�����]�g�7Y��W�u����r��:�w���jk�ٛ�-�`Tۈ���1(l����
��/����~T<M��Te< ׬-T�5j�h�)ݡ^��ڌ[6��G�h�|ի��v����ck�E��=�2u��N��5td�������5�>�Y��N��vH�E�h��L���72�7s�d.��b��l�J4���џ8�+��Hb�9�;ي}3�g�G�W���9�|��}�$�8�$o�z��Î2�[�,޼�t����s��W$��n9�T>����v>[�!�.�E%u7���ޤ�{<�򍤌�����t�p�@Vq��S.�b;��%ʲ9�G������j�' �6	0����@}+Z����#sw�0��.p�KZ'v��х�F�艒f�j�ry�{Ar��K��?+F���J���u)o�G��C��+����ZPn�· �3@�`��E�����z�48����\%�c�NΩ.�����}���s���LBv��TsWpJ������t<��+��d��l��l�y2����ݎ#���Q.4K8BU�q�z��Dih�%�t, |϶�=W�
���@��~�!I!�v�=,�}��-��$.�m�����bGk��CB0�D�=�?�0j�K��v9̼�� Z<α�8�o8>h�|��Z���"��x
�	�V�(�v���y.���"M���Ա0�U�-��>*]�v�S`�L��~�Q{�+D��h��DB���B�	[�Sɸ�&F�&H'�G��j��[��@Z�7[�/�_��s.�a%�����_L8��h=�H�ٸ��)���J(L4{&lǓ��V2O���ٔ�^8k�a�$]Z>�GUSd���a�^�F�#Y��d,�$8��x|��n��@k�B��`��=��1��!�K���(����"ga�P=��Q"	~�f����:Y
Jl���E��q�+I��B��k�HEj�I�+�c]4�9��b�ٗ�ȝ���!0*��w���oq���x`'/�{
6���VCX�n�ӕ@��_��q圑�
	2c�1��b��/�3��/�@��D�:��iatd�Ϩ�O:����߹�����d�&���5�!�1�YK�U]�\"�m���\{Lcv=��E�����)ua1Hs ��4��O�� �����j�JJW!CN� :`�x"�@-��%ˬ@�+
~s�/4܋��QzDJgy��������~���F�$�JiQ�8��i�h�2�)b�Ȩ�����Lǧh�)+Vga�J��ye����ij����mL���sh���#*TT���9~ﳦUtV�.(j��'��)���8�	�.��E'sO&l�����:��΂~�1@� �PS��t�܁�I;ͳq��0���C���:d�lX��K-�6e̱���Ec�B"��V��[�����r� �@����/[+f�_4�3(^6߁lŊR���-�=�����Qb���[fHpF ���Ȣ�m>�����t����4�vJ�Z�J 3��ČAl��W/~����ٝ.rW���:	4z��J�@{�ԛ�#�O�j���R�N
��@:Z3򵑨O�ll]��h�	=�F\}2x�P^�Er�5�F�G~�Q
:,1�HB��6{�*� 1�%P�v��<5�bc>՗�p\���^��Te���n�ф��C1��g& N��3 f�/B�M����Trә�t�a���=���to1hWrq�\W��I�{O�ƶ;I�Q�:�v�����W7�yV>�Eʟ����7��+�ƁOi��|�٫Y#ny�i���,!)�󻒸��Ds_X�h��S΅}�}W�!�Y���j�+���=C�.U�Z7�7�c\F�_G�tK>��:��:�7�k���zs��|��8W�V�7Hs��I�OC�K�,!��{4�� �V�㣩�n�v<��'���]b�pX�@P��d#�N��KkA������	�;2��\۷(Ңm~�c�"�� ���%���׵_�sF�.��V@��'�D�x/�h�[�FHѯT�	��F����<-��VN7UH��b	�M�A����y�&8�ؗ�:C7SQJ�!��_�0,
B�g��Ss���}I����������'#S�^��]b��QIͬ�_�Y���Dw����֏b��JawȢ �Q�O۩�iȅOc{�W8۽�G�2�= 	͏�H���ְ���@�C~
���m�������\{}o���0��ݧZ��x���/\ۡ�,�2���j��
�[��}]�}SC�^�l;@/���Q������bB2�7,�f�%����XMokNYApx������X؍v=%��Q]�n��@�m�)oW��V4_6���$*�⓺�0������&Y2�����7-�A�S!׏j�6��0F`��\�0��,�H}x�Yi�Mx�M�kU�����&k�h�b26�jذ��X*��
1���0ZLE��'f�K���6p��0�X�M ����=>�{�vIqK��X�OrFb��S`���jR{S�.WC���K���I��f��j��|f���0'0p�Z��UW�@�W�O�f��mN:�9&�zz�.N��)��(x�J%^~/b`�0��k��ON��L0,�T�I�e�0����1���y�9/~6��/�d���d����XsԿ�_3��^���,	��nwO� �6:��oQ4����!éG�J��Ġ��NB�6#�+�8�sJ4����E�=��B$�V�>��d��bSݟ�}�X�;t���To]b��gjx
��Ɯ��6��t��w���K�'~����"*�R ��'��L.8ٛ Zq����J��Q�϶���d����P��K|*P��~Lz`J�A�O�jt+�;��w�&��P��OKB����ú��\5�I�=x��(��Ս ~�A}{�22�Y#�Q���	�yX#.��ei��a�&�sR��xe�s5��	efͦ��½������coY���~-�gahp�f\#Ī.~��]^�A�v�q'��RJ��DL�wlۖ˾�(�׎������8+yEM0ݐ�����0���9�ݸ��=��(�#�0��Ά�JF�7[+���Ҧ�tA�*`�;2�����Qhݾ{2QN�(�r-NT!�'�&I�'$�s~�2fk�Oi/�9�GvX>�4|��G$.���P
G|�a'?e׷������B-�t$�B�{s�3����9���l�/�a�:X=��.��DI�za?.���ȧS��C9{r[�)#�v�[�G�ct&�
_�d�u���6�e����tEym~$�=�!B�P �`�C;�I�����yL�����8�&9����@+ڂ��k��$�2`��ӽ�O�v9V����j�	��~�x�te�?���ce�q���X��C�Ζy��,��SdV]cKE��Cȼ����?��錨���HU������j���-7�C��p&���B똍|�+h=!����=8Ҝ��Z�t��+�����j��E�#�`�|�៝���I�[�U�Xs`z(���(-���-#���j:��K��_��FuP�:��N�)X 9�Fn��,�)�n&�І�[}����a�5���Km�����f����B�-m|��c�9Q�KF�P�N�1���*/�]U��Ѹߙљ�� ��,qq���Iq%3$l��.<����6�!�,`h�(���0�BMSq�ө3��{�Fx&�yU����y��$�W��0�zt���p��T����Dk��ef��O)��m��PoQ?�Uۦ����+*G�;�C��hM�<C/�8�oΐqva���Z(z�L���⟭&'9�%zr(>��y~q�Cʥ���&�վ9c�2җ ����p~��5��A�X�grb��Ej$=���F�W��~�$w��F����D��{uP�.���7��2!�Jg}���M<���䟥a����4��t�a�m�N�ȼ�=�ˁ��8�ǜ�s�'� K�^L��m�3&�������̱�r�W���vlE����}2dL�I��yMÕ�#Ff�,v>+��]3�̩��Y �,vʃ;�}|����h?2��b�B=l6�d��
�K_�{��J�!�y�-�ۆ!��i'�-Ux5H�|��8����wG�q{��t����?�_���9,��6	b��i?��ΐ�ʉe=�"��Xꭓ�E<�8�EB�@���G�`�#-�O��RV�'�~�3	�݅�h^��	�%}��I��F��v�oF��>7�"7�5����N'�Y��j"��;1�����%�y���Z��E��kY���u����
��s�+�~�癘�77�gJ��i\���c�m���.�/��bAL���o�_�vI��y��U�w<p,ԤЉ�a� R�5M/�i]l���=F�c��[a5 �-)���C���I˱�P�c�#�
W�K���wlh�Y�4��t&p��0C�m�6���� !~���z�B�\��J��VI�eq�i����K#4���֕Z���x06@���g��>����s��MqJ�"4������e�}b($!?��h�\[pq6&5\��N��s��m���	 h�>k9��F8�x׉��*���6����\pQ'���,x1?���S�읋�F��a9����dا��bV�4�lp��������]�n0�,��ۉ8����'�b�k����a	�d�y�} ��k*���q�L](�7*T���]kp���-`ƹ�o�e����G���^��;Pe!�'�����h���6I�g���� ���c6ƣq��~d�1�&�t��44��x��?���a�};k9�ښ/;�Ii[&���*s������M�1�$�FQ�5�X[���Q������y1�-��$�!,��XQ"`{*eO\E�?Tj��>�789���{��<��xNb�N�&�[�}����|G�qk��Y�n#� �"�ƴ����2������"��.����ScK
	@B]$�����$U��kF�o����M0�FRߛ'bۓ��ٙý�Xb����;��=$K|iL�4����$����Tc#��r<#�X�5v�����?����ͽ"�M-6ü����rFݢ�"]DMe'�V6�V7�{P�۸������؀�C'�nC� �wD�%�t�x���*E`	q� j�	���솯yx�m�r��y�C]TS�e��g�Yo�dl9R��8�^����hM�9+�� ?�-b����ҽ�_=��ARW��\(��aY�V������3͕��z�����;�S]�M oܨ�8�@��M���0�F�Iw�r�n_z!�:,��7?gSf�؈�=i*�+6Qzo-�����T��L��d��,�-�J��w_7�ޔ	�*������P�Z��)������:�M�"u��G
!��6dg�j�~)Nb��8�孭E�!�L�+��(`ꏧX"���񎤽V���G
�(&�>���%`.䦕��}~;�����U���uy:|�̨�ĵ��Dv����f���r��ch���E����sY�F)�5T ��-������#�r=!��$RJ%��>��U%���Y��@��Sl�Ҋ��o�)5URW���7	3+�!b�J3��p��{�blCY��I�<�������,����4mӣ��yZ�>5��AsC|H����Tj*O%��T��r�`�
���qp�җ�tU/�Ծ$w�3Ƴ7�����-��N�������n����[~���1���`�(E}-nb�\Ӎ��oMd���0� ���nd���Ê� 爈���寠�� l���ruק��D�Z:^MY��V��E�)@j�0ج���ă`j���R�vҐl��[l�`��-��`O��<.�e�3�7�4Ā���	zp�����}��A�44���3�'>9�	�3����R�ػ9on
�zv.�A�U<��[�C�[ʧT:wo��RyvS�4����To8�S����I-'L���!49�AAU�Nce(V<˳#hA	f��������,�C3���Ŏ���p)W��g��y(�H�~��Q-�B^�}/��\�s�,�o4�ڶD���,h���ڥ��Z�PW��[{�R
��g�O&F��i9�CVsN|C̒%�?�����ij��F�o���WU�×��OZ3eq���0k���J��ޚ���H�Fn��qv�$0�=����Y�gHe�d/b��q��W/���"%s���^� �Т�Y:�W4�_��d�a�8���	g���U�"��]u ���d����"�p2�@������.�$��VyWj�����E^G�@®�*9I$�Ls������H����t�5�� t�9��׵9�g��!�[ӽ&-cg�f_�tZ�C�����!01:�T�چbD:`S�ʛ}qk������AIb5�ζ��Д�����Iz��?P�h��4(۬�m��,/[���/ʱnW�wр%�]�B�|�]��/��/x"Lj8*]��K�&Cn�I��ŗ2�;s%�s ����1��>�SgĎ�����r^��?`�����0t�ѫ)%`YQ6���J״1���J�/a�+1)Ij8,2*<0��5���{UT�:6��P����r�VA��PJ�@=Ox�y�5�i(�MB;�oT��1��}�~>Y[W���]�:L��"��:�oYWqC%p�w�AR�ⷅcX^�7* R��񸕻>q�=���T�:`���c�c��~�$�]��]�)=�'o����?횼-9�iʫ=K��(U�U:+U�6�)�3Z�"R
��S߮�Hh��]	�a��ōyjLB\D��a}����!�}\�㔖(9�Q:����*��_96ڹ�O��/&%�m7��qb�s���Rzx��q�n{ʯ��L�!�	R��f7h�$30%0����>'���I�whl.-�(-�] ��#(򩧼>'�ǉ��'�6�P���X��D�������D�k`/o��i���V	]5���udg��oz�E�r�~`,浫��_xJ8��G�Q�;��"��vqO�Y�_��^,�$-躉zG7hö�0�k5&�Y�wP%�1�V�y��! �����?�H"���f���Q� /��qZ����T�P&+��ߔ��)���ᐴ
�h�"L1;��7P���2:�ۗ\���˃I|07�#U����#g�Z(�6���)�##�F�;LٷD�Ѯ8k-����㨷� �K��^Z�s�y�f��������6�*K����,��v�k�e��4F\��:\�<��4p8���=��E2d�z���j�,WFǤԈ�+[q&0ݚ:i��*�j�&��ZSDӫP���	��nX���Hw��`�y�5��Ll'ϕv09N�f,�L���W��P�#��zCS����ӂ��!3�hT��݆c��K��"С�j5���5Xu)~D�8,*~�_f�&&,�<T��x��֌l����D �
cN��/����堛�\������ 
&d�=���e>/�f�*��6�u�O�oad������o9�#%2���0��y�c����g� G��g
س�u��ʇ"�U�Pŷ��#�8*\�+�wD�} �<"]�"��w%6?In�J�"i�вLU�'r%x~�NY0�m!�`W��\4b�0e���3��z�og��c��'-ď��GB�vl$����O)�f,��Ku��^�L��zVl�CjP&N o�#��j�pw.ŵAK&�Q�ݲ��T
���!?Wʪ�b��L+X��]d͝��#����m�� &j��c��� �jL���" �2�|xKD���d�^o> �hv�ѯ���|���"ߊ�v�#������n4Q���}�*��g#br���2L��x>Y7�&c��zi��i�zS��*���5^��!�Q��NV���e�jm-����1%�a��vQ-s���WXϤbS�?���}�=U�@��Gٚ���ߡS��H�81}ʃ��u�M�'�;�E��J�]@!o�6�SK�x묾��X��pD�ƐuJf!����	<�#DT��.YF2"/�5�����J�N��p�|�%u{���1N�֝]x�I(9|H���M�4���_s��~Ʌ�V-��&��<�?�':m2z+�i���\�˹R�rG����]*+J����"�a�rqSd����6�I���.�d|Rx�7���8�&�|���Dl���� �Ƒ����?��}:��9�?�Ŕ��]_q����OCF�Z���g��r~I��k��i��,�=�ha�z�ֹ���p�݈�@��B�2��K���	\U�g����K({��\���`]�\�|TO���K�9}��F͞�0�z�s~r��l����+/�O��}ߥ�ʇ8�e-�� ��k�+�EM"BNe��;'R[�Vv��<�Ӄ�ա'꼉��|,^���k��O�1`.T�S��!���P�V�Ho�Hڬ2&IY=��1w�^�7��_d�7���M���s�#Ўʎ\|���ʄ!�
�_�>������$��.�b��ӳ�O'¾c���+T����%��NC��_�֟��IӪ}�U��>s������H4���Htr
evHf�>�r�F>O���~��ES=��]�fo���7G�VEu�?"�˓oyc�|sjk��^>@s��H.�����i�����R�@\��x&�~��X�gya7��J�[���x���Aq��]�ԷU;�%�S�)|�U��/n�,�FK�if"���$zI��[7H��k>_�'�K��f~�Ν\(2.����F��i�4�G{����=<�����$�k(�ʊ�"S�΄X3���r�:�X�ʳ~�d+)��H�
�#���쑓m݌>������bi��'�7ǁz+пν�%�"S\��ơ5��#�U_b��/ۗ�0�:%�l�O�=)ܛ$M�`��<���{�@-)]⏚5�|b>���\�Cx�o�V����2xy���ϋ�k"��|�����ۀ�HH�F6�������Jn�Ĥ��I����js�*��;�lY�;����<�g��,���:o��g��M�u�?�ӟ��3X�+�^z�b[f�+�W�vO�_4W��9$�)�}_��%���F4I�\4�/����A:�'M��R��KT@G�9d����}s!�օ��)�N�j}ӽ���`����D����Y�8_��x�*��T׆F�(���]�1���o�t����VagN��2��v�.����t��s���.��'��y����\��ʎ��I��^-�H��	�Q�e�f��b�:��ۤL��ȟ��T^��T�3�������NQZ�`�p|2'�k�D/sa�$(}�&0$��t���D�`�������,Iӈ���v���h*X��{��p�dcSy�|�<���rIS���gr�5�ګ�Iʠ�3H����nˆ}c`W�żk=K'p��X��I��.�41��fH
���	d�rXZt:�3�_!� �)��������p]���RZTD��+�A>���2�������V��8��]��lm�w9k�a
2)$��}oT�
��t`υ���u�m�Ew&7@(��+vd�4''ra-���&+ی�'�ܴ
ik?�:"���/F��_�1�dH8ň��v
��%� f����r�$�������+xd(�u�	Y���r�E�Xp��d#M=ϧ��0��a_³t��;�ur��`��9޳8vr�8�ll,�׭#�rw��v�+��CK����Fn�A�twDo���6R"������]�V4�ݷ �ɋL��ʣՐ$��WY�T2���`�[�m~MIH�A�خ��e��y��� �B{�刳ն��+�r����%�{k@[5�RS��o�T� �B�Ƴ>��+���T6� ��mfD[�4�=�Вt�q��2����%9��%�����xӤy�l-]�,�V[e9�ׇM�@�D(���SK=@Zk���	��������E�T�x�%i���j�����e�ь��|2�a�6��H��/�2���F���m>#�-����[�xỮw��0s,Í%�3H��/�L4�Q+�ZA,�b��!_:�<Rf��\�U�,�jCQCu����X�Z�9�f$tZ��P�Ѝ�RUN(��(%��9�G�p�9=���;`�f��8Y
7E|�s�5��O�Й��1�	L�]���p5?Ȇe��7����1���kB�bL>�U�M��-�����G�yl�p;��ZnHM��k�Ǫ�S�\K����,�Q�i���G��p'�j�@��=��4w�R�f��jIZ�)���s�A%:K;��ߡ���3�/=h�<�c�|�I5�jj���Jr���D��Q�P+�� ���{��x�ʔ_K���g��,Hs#���8s��=�]�F��#8�BLbc��
��:7�v�rP��N�Y�^�Pp���N?��!P��Q`I�������]H8��,�C�J�J̽a��˩P.��"S���ZчWy�������lm�pq�����JKнS��?��M�1"�����ϑ L�E����ȨP�#ϝ�1 ��h�VJ9)HIY��LI�����z�@~�=v���@�y�Wg*7���k^�����Z.����6��%LA̗]ه"K�{ �@g���~'���\<�ꓯ���)f�<�r� �s�S��v�%��[��/�9TU�o�U�j9�|��?��c��t�2��r2��������q;�Q�~^�����he�=7����������΂iI��7||���}�貪3�G`Q0�{�c܅���["���5���������(+����~8�3D�UƧ_����'@+��{�tk��ff}:��B
�%�}/��ܺ��t'V��U�	|�ŉ^�6>�\���v�-�㞽fodHM�:�`w:�ͽ�ot�ݮ��aC�x�rj���`l&�E�а3_%�lH�E5(�~����o9Y�������Q/�vB��%�E�lPD]�Q\a>wh�2^�:dHq"~�	y�,�$|��u+vS�o��,RF�#��')0B����-T�\E_�\��U�w�79d�&.D�3x�`�QjY�Úp{��[��hz��/q�R`���m5K���&~(��2���j.V8��!���(Crkf��ˋ"�*����ۢU���e�?0����p!�v̊Ƀ�Lv����8Q�n��%�PS�{��Y�I`�S���U�7�>�n�˽�W��kN9�#��@�-����Nj
n 
���12n	�|  ׫D�C�7�Z��������	��5F�k��G�u��{��zr%��j됡�V���H��`F�ue�>J2x{��ƣ_�I�E@��8�6�*k�	�y��Ƌ ���2D���Dh�a{6kx�z�!ʆ���:�&��ռ��x�X=�H�oQ4��U�i	.V� 1QMc�����h�S�<V4=^�C�!\�i\I5b͍���R{ ��-PE������
i���u�B�Zam<@�	_�n������vt�������J���Q�&J��Y�K��B�}���3���[�������nvӲ��Ky��q���O_ɄU!��|𻠎�Cm�j�+����wu�����{���i ���
_S�}�S^C�!n_v�{�i���!�r�y���T"�����uJ/t ��py=�̴�wz����ʽ�dD?~�N�w���+?�&��6x���71f��j".KW�KBXى���}tP:�p��h��F���,�\��A0g�� {�C~�ߚ�>�wc��t&4)D��ո�H��E��+['j�D#LGio
hq6q�Kx��S�I��d�\�t�}.��p�`���� ��/9��9ž��l��?o��}4�T���d��-�����;��hq�_�&�)�	 ���3��tu�)ު��{��vV�7� 4�68�'������oz�ZA����T/�c���Q����F�A�Ao�٤�D�\�Ġ�{\����&	�'��-�5O�p1���!<�x��x�^��F"  ,~rB��\�s!@�x�W��56��Z�w�tA�q���7_A��dLY��
����0n!K��̔8�fY��5<�#&uY�	F_qV,	��'`DR�[vJ�N&"P����EC�@���Q���w/r	��?�_���tioI�mܹF���2J�����uy'�ǣ�3Rn41Y�o/��ۢ���n�:�6�"��qݴ�S���9�Px�mb���,Z��R�X(!X^9�Q��j��Ъ[��I�zf*|����,w3*~�嶢]��gQ��qk��rqy�O��q��������-��.&,fܢ �e@&�Q(�B�WE�`ZyJ��~c;�G�7�/
�<�`4���y�rr�49c�p�f
:G�p;Z�Y�S�� �y�i��� <t�	Icf���o14�����K��Y���tG*Lv����ev��?�����lQ���6�	�L���D�Ő#,"t���mn��ƌ������G�.=�7~�E�0�02��yk�EW��T�� ����@�uu	�Zx/�꺈(LGj���T����:�h�c�l٪�b��o(�c2���o�
>�~܁<����\3��-]��cRwv��q�q^��o��\����2o�e�7��ɐ/�:[�x��=V{�0���nC\�pC8d8x��h�-��T��&y�����d�\[�Zq���g�@N���w����Z�`��F��g�Xy��E!>\wg���S�E�/o��	c��A)�5�y�~���Hk�b�l�t�1�����c��V��0,�e6w.j�ϻ2"Σ}w��]}8�1.��2M����6��j�9�S����,���?�vwM�� pd��q���s���ޭ�$||󟌅#� l�={�L���[
%	M���M�иS�j����C��^�xM�/;�2���灼2�/8N��h�x�xO2�DUK�svDUZ�������r���z(�T����kH|��tI�ѕ�?x{"���c1V�`��#�;� ��oS����f2�m�!�!"cbw�.D�V��(v0�%wB����mݡ�6���(k	�wuREwm�M�h 9���UJ�<��f2�>4) �(��~"����k_�`��"�'7	�d���o��:'�3 Q�c��e�+ �~3�/�B�E:zFW4�H��d��򞢮�)��b���g^&@�8��M�+Y��#d*m���z���Đ�ΐ/�oY�.N�e�=�m��L�L�3��Q�=���?(���8G�7^F�q��4�ֵ��"�W
�@��s�}�9g��%�ˎ���k���4������/^���2?�Q 9\j6[�v�с��\`v�6Vw���j:З#oxw�iU���O5��vS���GibSy��Hj,�BŜhE��FH���D��2PW;�Ӟψ��j��eY�#|Js&Bm0�� \��c�('T첏b� \�@.���B��[��!dV)mt�V�\�v��<v������}"� 6�ҹl𷧕$c)�[�t�@_�j/"�}).������V��}E�So�F�������=���������0�_���P����5R��Z[�o�O+�����[;��Y��ОIM��j_�$���
<SZ�ݭ�@���N{\�D�MЧ��m�̺1�������v��1pgI��Ld��z1O�������F��� �W"���؄��%g�������3�-����J�XL��2�*CYk�Y9��$��F�'����d�!7t�/Z����N�M����A y;yy���$ⵘv�p�;L�,�s��ը�ӂ�9��X�e�7�a������P"� ��p�5q�J�z�h�����@a���J��eF��C)�xUVh.<t�y�LԘ�(#�����COY�b�a@�;�� ��.�]����D��h3>И��t}�Atz��29kf�#��|7�>����r��~;7«��>���\x?�㫦�*�53�V��r M�s�]K��6/xIH�l�W+M��p�27��=>޼�H
�Tߛ��B.�(�{�|�P��*�]�%q��VY��h`6�$&㰾��Hg�'�S\z9	r��Ja����c2^C%��Q���m�
�w�r��� �g݉�6������W�4+[�^ ��;#&q�5��3��g!.I����1&O_���g1,R�W��¿��&f�H��$�Fe���o�x�/:X{��5������x|L&kj(#{�pK��%�e�L�g=��b΅�?���� u�������5�2��6w#@?�	�����[{<hg�'��χ�0�i}�l�A�ߦ��7ryj��mS���6��||���s�niy�Q�N1��Edc����3-�G�7o�0��O׭�缠�Q X����)�-��|]e&��\<����5^2�1Y�tk�.��?���N���k�؋|�5����$�g�e[w�h�Z�cM�e�Cl#��k�noCZ�¯�d����R��:��;:VrCΗU���Q �ڋ�1��\�lf.9�t>�����.�����$�g(��k��� �O���$e���څ����S0���ɓoxtuu���L�{�UK�P�yjy{���%z�8,��n��՘[��
P�%?Q�7�o%(,�/��޸��غ����<�쁛;S������ؼ��zA���Cҽe�A��a<_7٢�P齂(�	�=?�7�eX*��i�eV�e����h��<���eQ�Z%V�0��&!�+k�ri	�¡9�xB]�L��%*�L��w/W_A��F���]�y�F3;���힯�s��(���gGY�W��g{���+�;S�wY	&C��63��,��Mϑ{�\�^�GC���4�懌��%��NQ�b35R�`�� �lb eX'9��?34��ಐ�C��d�:��2�Z���l�+�`UR��Q���p��\!|;V�	�9��N"��`�tQ3�R��fKL{�<���3� ��$ٰ�?���l	���c��u;T}zxg���k�{:|��f�����+���V��n��r=+�T���h*XV��� ���RF����E2鏫������}��>Ǥ��ȅܩ!v�����\ɠ���I��Z>��{��T���>���LE[������d��H�����ɘh�K/Cb�R�c��(?�L��"-�n�L"��.T<>W/���'h���zU�\F�~���m:=�H�[R%n��VB"P��������5ۤib	��OI�ڽ���0��� <��6p��:���CF*��9�8�eh�2Kr��D��/��V̇��鏟����Q��u*��%J��}��Z�BݷV��H:���%�(�2�8殸9�Q���XV���2M���-��t��ր�Q�O�u�K�*�0§�`�\8����v��5?@��#��|��0�y'�W�Y
�����OR�B0�.�"�U����v�����M��;��
�K��6?5�'5ZT�k�|�1Q�7�*%̝�H� ]g�̺�pIU�}�lF�b`Q�ҫ�:6~GC�nw:���4�|�'��+�P<��J$(뷤f~5�9�2��hm���T� `�ކ�|�g��gg;�c�a7^a[�n'*�(�b}�(,��A����N��8��/�kA�G� ^�iˆ/iD�Р�[�����K�� �Om!�9�Tb�N�
դsS���Y��ik	P�x�&/
�
FP�B�����ӤF�#�����ӄVH~��̻]�ƫ4V>�gO׽��Q-1B?�S@��T�/L�0���ؘ�4�E�>�p�݅Ǐ�7[!m��6"�O�7��Ą,�k���K��R����q��y�Y��ߊ�9kf�1_�ETFK$��J������ M~|Ad[R�W(ԑcf�yW�/>���r�2T�3�R��"��Wז��zN�_Hq����Rh����?�g8�.�B��cА�e0'���"T��d���np>ݶx��Zq�¤p���%�U����?��l�Vo�ޙC2?e-�k%C�o�0���g���9�`Sҡ�I�H�@�.���IC.�\3L�R��t�2��>�����l��K�\��u�zrN�>��g"�*to5J/;s5�^�l���!$򑅔���`��=&���ظ8HW�
̯8�t�$��A�Oz_q$�QK/�4��F�]K������rQY�/K��ަ�t�R:TH��$ 1���@��&-�"d_oJi�D�ufW`������{�}�*_";�
�=�;,�(�ʅb~qcR�T?��ݓ���!{��ޝ��}܉�RXx�ևAؾ��	7Z*Q�#3R0gf2� [Vز���A�?+O)�*�K&U�6H�u�7R�[��/��!�ۅ��]���֑�r~P
��yT9F���mY*<'��\�i��}�9p��];��AF���?S�_����$G���=�꽊3��:|����l���&����,h)��C*5��h*Ǒ���	����u�	�P8�	��-��B~�L�D�B0���	��ۑp�L������9�;.&�����W�r(]Ac�����4��L���ך��廈O�/�s����.l5Q���4�̺�>�]��� 4���V�Em�C�����+�Lk_�k05�ݚ{�X'xop�,?B��ձL�\9����f���}��1����i*x��e���y���/�7X��.Ӳ5�|Ͷx<b!�y3@��Et`�x��p�����$��r�a� ��<������|G1�3�Q`&'��Q���>2>xV�[�z$L�3�e�+�x�wї�qHxFN-��[�U���s��o�.��Jıc&�?VlK=5�����ф�;�$Ki{�4��Ǐ��V|Ta"��G�a�<9������2�ʿ�܂��i�ފ�f^�K�T�[5��0�D��W��`@���j+ N��|��q�ƭ� �Qb{O��v������������b�6�ul���i\��,�ej��l7\}d��TDʥ =�
۞k/�ʳ�Fe�^H��q��)}lۉt��h,�1��%vj��N����`��i�+E�6w�=ڿ�x9
��Q4T��܆Uχ�"ϻ�n�(m9ɮ����J6P���AJ��_-�n@�KԬbL�B�tj��5*o�jjF�?�	��j� "�pC! �� A:�Ү�<��FH��b��&���S��R���Ւ�y�K��5�{�/���{h�����l�+yT��$��u���Y(QRt!��Gϴ��$��M��p��,�6nc.^.!���ݮD���~���)A�k|P����v[�
eh�!
چtD����*z��|
�,T7/dX��:�a��먉L���hH�Or��5�{PT����At�3���x�b&�W!=-C�"������U���U}X҈c�K�H|o��s$��ڇ�m[X��B�b�I��_A�����9)�<R��6��׮p,�Q��n��2+	�x�E��ERXfgwŀ��j�M�5�V}���TFq4@������a�EO�g:Y�tG�V%s�]e�H-<~ȵ#�y��1�KQby��l!ɾ9������I4����QÁ����1��'k�͂�d�%d�\�,�7R/��O�z��.];a�/��3�>oz��K���5�삦�[��*��ݘW�S`b����͜����v/n�U ߘ!��5H���[&���v'�#_m(�R_�5]�w+��P��d>��ʹ"c`z�7��3��;�vsP$~"ӾIv )갑2 0��=lM>��Mj"_J���|O�w�'�QI���M�K�Ċt�O�\r	^�[�LƊ���I+K8�����J?F�Tk�r���9���i�Oi��E6V"���N��� ���bW�B)�OD�<�v7h笇YQ{g2�]�QK����oX>	���1ĺD��ћ[�5Y?�0fwd�v�	���H-�/�@�GQqUm�ϰ,0�g����xM��U��wrD�ql�
/%�������I�A��jv[I~�f��I78°Q�e�
�h�B�jԗ0�99�����_�v���Zʟ�	Z�m'��V ��h.�ɧԽ��M����Uǟ�IRڤ<��N�娎�99��hC	�
�TR{�[Gʒ�ӟ݄p�7�A&�D|A�=�Z�[����6S�E���5���k�g�bv@؋/��ٲ�8�D˂J�R+̐gv�傺̮5+c���V��AR�4{�
A 9MF�Ff���J�pN����	�5:�oГ9j�jo���v8����\Z@�L��ι̋��M��}�'Tap���l��$��nȈ"M����_~wzϺ��@=�p[N��d�yg�c0(�[���q�GK�=�&��qc��U�xK�wܱ�^���!��0��Qԭ��C������b��4��}�=�^:�*�����i�/�������EA�ɯ=���j�*�!�`4I�S"y:H���g�qb�2�*e=�<������7P-�p�nx�	���+	��8�kmQDA���X�ݍ���d����ا���4Gp�NI9la��zS��>�L0��qZ��7�&���4�d��)���K~�W
��]�\fh-~�M��.7��mm��o���`4��iM�5(/S�%���seU��0ঠ�2Nu�f5S�!CS��.{���q���>a��)���C�&	V/���ȁ!�����|�+A8I�m$r~�P�_��g���a�'��L���mL����/�����U>%��O��ZE��G�<h/�s@o���,z�7�_<��Tg��&��O���'l'n��e_��#�#�MR���l�K��b�R��9ӭ2�D.`��Im|]ssvP�C��'���M%���:"U
%�����M_сf0�E*j2�AE|m*d�G��k���)����45KGV߮+��ʫ�2����-{dD�v�:����Y�������c$G�?eig��kJxZ���)�mz��@5'c�ʦ��bx��ĭ̎$�� (b�(���ad��D�:=Y�����k��ǃ����+�����hڥUP�Y�6G�����6?�#�l/���~&�2Ur����2$��o�y�(�@a{������&�\>`�Q :B��?�M�2T�l�}�=���L�#��Am� ��������I<���Q�֔H`�!��e[����R�@��(�X���[eGI0Va|��z��*Mq��74Ȏ��]�p���)v/5��/K;A�)��}h�@i���)�w�VF�� �0�L���y��l��c��0+��	���LN"5��4���|iR���O\�~�������U�M{?��E\m	7���)��ek�Tߢ�j)����8a����+��`��@4��2$!�=L�`h�=E�'E�wE��H�_D�T����ҹA����������'��B�"��J��:��D�n9����%��:�o_�v��������w�H������`�@^t[���s�/�`�x,���E]�yL��}��^�O��r��:�?&:O)�^x5��� ��4�ڇO4�k��6���T�:DMگ�<����� ���D�F�o�+�V&Z!�S��Y�t��FL���3�2�Mx�u?��~���Z땁~y���wPEŶ`V�RF"Ji���n�G޿�r�Ln�Nl�$�h~\%�6�=Z������� 6�{�v;N�*�g�8!��<���E2��x�-�t��<�?=��])�U����(���=�U���@:�vˬ(Z����\�ݐ���A���E�����2������b9�$\��xщ���)���W�:�$eЭ:4QE�HG�5�Ъ��~���Bi�ܒ�sj���n<c N#�i�B�#P��2v�~?�K�}e�m�	�]t�u��mDQ�̶�
��(��%���n�}�q�
�ϕ��~��/ Vb�3��q��	m=؆��[x���@�1R\��L������p{\��8��bFv���Y��s)M���&Puh���;U*|�fU��.�ڀ���m��W`�;��Y���q?����S&�=x9Ė�~��� ��_�wSG(X6]��
}@�u�I+lט���O*� 
����|P
��+�+��Yb����������k~��{���.�nV���9.�ñK����%7<�_��1NGK��g�Xk�f�gھڐ�������+�$���l7��d�R�f1@[lDA�`H�i	*3�����g����Y;��/�"�{�����I���1>��m���-�`�V�"Zr^퐽�͋��nB�u=��cĤv�\|SѰ�UA�OW.��V�!��@����+�������/U��~4�S����vW	"�S���	jy����6����Ī{W��H�3G���]�����s����NAH�U7csuK�_6���1������.^5��啫�#L���~˧�v�~ؗ9���$t��9�Q���?�{i��<� 
W��*L��|����ʳ�U:�&�u�B~�8��)ͥ��@��[���H�(�Z"TU�=O,C���V�l�L&M*#@�L9�e��z��s)`ɗo`����1�2̣�YzٝC]�H��ͦ�7a�r����۲�"O��>u��]qm��'�7�u�1�YS����@X�����s����R>�5���Q�ePS��<����!�ҭ�
�ڶ������VV�D<T3a�R�j�Bo���ڞ�T��m|H����OС)Pn�M�e9pn����+���ů��h��(!�u�e��Z��T.8(���>x��F� wZ{v�rE���#]Rnz�v���lGu�|I}`�B	u�r���M�����D���B��z0!�c�y�J�O���HO󿬨@�M�ރ%F���
�'1+��a�旇-�A�Ճ��e=�=�C�6�;$LhR4�~�&�J
�c� ������rJ��%}X�|U;�U��]����vҧbT��B$� �ǆ�Ř?�|��[o�p��PV�p3�@�K���"/�db�;FUz�[���$eJlS�VB�8^��@)t,���>�7��b�}�&N���J�"�����{�chU�樋<�ui���&7�	Y�n��v���V<?�8OlOHGdO�~����gc,3�Z\���p��y�����k8�T����ލ�\	��$)�Ԟ�9K%��ϕ�=�����@ci��!ac�)n�]>G��?��^-5WXj�'(N)g#��k�ҧf�o�I|fl3� (|�7���J[p3@��ZC̵����i��<�-�C����U	���Ou�[Âz�hi�l��:{�$��GEʝ�[�n���������F�Wk����V��d�J����~�~03�lV���֘�g���)���\�9/�������I`�<�l�2=Q�';W�zp�[6I���#|�+�Ŵ)��2MOS�%��<��Q��j:e����y�^0�%��daL���gFc���.4�4�f��	��I4��rH�P��
��]��{++�k��<��:�&�� �?�}~T�����3�
���n?y`G�nRUٜF�e�_�S�Ȫ$�*�5������.��z���TS��oD[��̣�����Ծ d�dE{.v�����f���f�h�\�����v�-Ra�?�X��U�ڎP�h���w���6)����|u2ԫx�=ukT�|"�mXܕd��Nv�`��p�Ѩt�W�{���$mia�c�jP[h��8��>���}�-�V�ȼ�ٲ7��M��Lφ�Sκ�%!PV�>�S��P>��W��ƎΊW��og��v((_�Y�;Oo��������<�Y��c}H�:w�,� wc#�� �4Vk�O��[�|�k:PcG!0�Y����P�S�d޽T[ >�'���B�a�����T��߇k.����9��JXcZ�O��0/��kawߪȨ��u�Xԥ��m&��%v(Ǚ)0�"A�+��v
rH���i#=�ɂ�@��aI=�#6�w�t9���?'�W`m˺L�{��cr�͋ej���9!-%@MH��=SpSz���l,,���e�b|����`s�"�C�X�5s��0�,^��{��ۗ?���׃����1i�>��C��8"�-��S�p� c8��]�
�9�	�K����e���
y�xr��w�A��>���P+n�&�!���|3����0�m�s~Qb�����'���v$lO�{��(P-��&�����c����LtN`�t��&�=��һ���T/A��q��ݪ��z�������jPwݸyb#P�<�uk�i0^I8.o[k(p������v����s��!���(^4�_�E����B�O���L: WcӁy��7ѱ�?�I��¾�5R7a�D��濥�Y���!1�S���23i�l&�k�XL1ak����m���$Ti�����P��ē!A]D��4(�9A���]9�t�7�V$��Z��֏J<{��H;����˩,f�~}��uXDli��*�/?ˀr�b��(��`�"U
{��������͓�������@o)d�i�u���>Ja,C���"B^Q@}��"���-�0^sU}�c��-ߚ���SG��ET;��Tp�#��xY��\H���њ`+��2���63��HYg��:bE��#T�&@#̝9V�s��ĨӃ-q<�d��x!��������C�%��K�����Γ��]�|B��ȌC��R��?棄X������ߓ�o���U�6I7�<p�&Jp]A#�<�`��4��Z#�_�x�ݹ�<zpL ;n�)@d����y����h؄�4�3ݴq�zD�Wd-(r5��9�}y�9n�`�ֻM��z���lT���������V��mN��&�����$����{7�/W��s����-��ψ9.����O�u0\"��XMwz1��B�=��������*�囨Rvt�;C_E�����tQ_D�{g�=���y��νb�(����nR%"'��w���\%I�h5����JAt�2Ǭ��5*���<z#o����cV6��W�o ;���k��_���R��7}+�i��?e�2@ԙ�WށC�C2mY�̸l,[AT�<�L�<g�l__s���Yj� �ݪ?r�(N�`�`S�� 2�vք��ˏO�pV�;���	��E��6lW���E~<�sqa�A�%���p��p�T�^��[&��t;/���:ftR�y�z[l#�fhX1v��Xݲ18U��BYLҰb$���R��"���^C)J�A�E7�{/4|؀�[GTJw+��"H���.*&�q77P��gi�gƦ�)�e�w�[��l���A�*��rу*���~]�B����\""�0s��U�u`!�T��mB ���dm&�A��ޢ�J/�T7>I'Jt�/��m� Y��`�;A����I�r^�}�=�0MD����o��"�.�l�RB/>'�����^���\���se�Ɯ��
�8G�������19�]�Dhپr�+n��r����me�dU�פ�r f�$��8�N�J��
D�G�i����q=D�Q��c���K9��r�vV��mo�f��H�����e�[g�MԌ�#A�'������P��8Ş-�6oQ�'����v{�AԆb�N<Ӱ�7�H��s�N���,�J�8����w�K}b8�G��(���sO�Π!�����Ϧ�ez�����!�R�x�SK�2�p�'�ݞ��q2E��)7�3e0��V�O$��m?���.�ժcKۜdy�����ܫ\ri�D�\��X�p��O�==�~�`5�CP���~}�7������s�I��X���ꕶ��F�?����8��;��w�j���b�� �@E�z�*��rMdU�=*t-^�[��v��ZSA5X	�T Y'�f�)�{du��M�@[��3ʑ�M��&��j�����IU�!8}z�#�� =ʈ�N�{Ew8
�
�<N�ߖ5W$Da���s\��У��x����.�H�,>��S&�\!�A�V}�=0b2����:(I"�������O'���Y��i���>ƮS���d����|�GՍ��bԗZ,��"~Ϯ��)�/4�*t"�i���r�LU��y��P�Ϊ�W]����ƣښ��?E�Z	�����;��0��^��I�+Mި�%�`ĊO�w���W�J3S�@����6�[����A�L�6X���3����[K-�מcY���c����&܆p�VEF�7*�(t�:N7}��z��΋�����3��f����N�\�tk׻�/9�Z��ZDq~K?p�L+�|���hXf&(8į��gm����t�ʠ1��6@���t�R�[����I�}Ib	µ܆�:D4@,�P"��Ԣo�Il���ݝm��D����je�K{�ڤa�)���^A�[,v	v>���(B�U|@5 ���6���|t��۷#\˶�i���2�G=n^�D���ۓ��ډ�g`�@�X�vV<��SÅq�>T����i�����"�^+�xL���[��Q�X#���a������G����~#�
P�=�yh��D`�
�Z{�t�Ny�޶�u���{�v�٘����*�SI���DԼƇ	����i���CA6�����&���=��-q�y�ߖZMݐ�/=�o�l՛'�*/���4���nl:���ڱ���v�k9�֗!���1��47˲^�s�(@V�څ�9Ba�c4�/�|!��I��������QhjZ�u��)'i8ރna�TQf��(*z^�A��M�6~T���0���7�iu����QT;�8�d׺s��t����퉟��{gjdv,|�퇒l����'~�.�BK.MUN���2��)� Q9��8�PB٥�`�
��:��7�q���Gy��jO�=_Fzq� o�g�Ã��FHk�|� Fs�]�-�O���y,����7�tg���m��H��/���vO}�TҦ�����V���|�7��p�V*��\ �sizy�S{J�\��2��K��<D�\��;S)��B�rp�n����u~㈦�82Jɻ����h W?�ZD���L���W����\�+@1Y?�����Z�|� o4+Y1ra|px�2$����ugLn�:�q8d}'��\�R�(����oԽF�Z7ةKb����r9�ii#@:>��y2J_r5UT�8²�~���l�/��?zx]���w������N�*�S@�E����
��H���ӆ���]�Y-)���E+*��>�؝��)��g҆�ʒ��z��jt����i ���o9��&���� ���/	���	k��eJ3r�LvO&D��PN�eD�b�o����~��u�s�M�,֍��!1~�De4?�١�V�MGW�ns��jlx�A���(�HJ��D�B�����;�-�����@�&����>R�e�����LO�H�����7�l�Z
O�����w��iH��gB
t�/ ]��|k���7Bv��:�^�p�YO?�%L� �E9�9���8�괲�b�A���,~m�xԶҠ����Eރ�{�F�4VpP��G�G$e���A!9I���G� :竱�@��z�8Sg��5S�m��-��ɚ�j���"�����7���/�=�$�q<��M+o��t�!���+��I_�3e��D��H�7�~�iwALN�
6�`�JYE�4�y�'�����bT�f����!:i�%�e2�Hs�t����8c�s9y���d��,�ՠ�ˈC���<�xG#ə��ͫiR�u����<^�!e"c@7'^d���4}��¿U&N��8�y�{�q�Ws ���N8�Rx�	G�ෞ�mY$=+���?s:�����|�a��Ј9����t�S;��0��'�E�6�"�Y@��� c&�NT�����7�(�~�x����:�]�����Sa-j�~�YX8����H
:3���mj���������h���SL,�$��5�E4o�{[9̢ެ�`pV���X� �����\{�/�h��ʂ�;?��>�+eH:a"v����M6ڙ2>/@��?�\���$'���A�mۃ؅:����$�l�6��|IV̀ B�cU����]�	c��9g�ڙC�'}'k�P~Nj.5����*=+[,d��&.[�{�}��PT@E��.��֙r����kz[���aa��݉�W�RmQ� ��A�ݏW�t��H���T��"��?#����̾�۷F�/�ȋ���X���T���;�<$��k�ɫ�|�� ��6��q�����������ZM-[�e��"|N��x��������sBvfD���^t:���'�4`��"Zq@$�c2�J5hHrr��@ Yh)-^�۩��d3QUX{��FuI.�*�Y�|*`�G����DK�s+2�9�;�轑$�w�Տmg�	�A׽�9�-�
9���з�Z�U�ϜB�@�����\��Bh)埍�Ո+�� ��ϻ��	�7��G�8�ےZ�HF��O��x�N��]�莨�?�?��Փ���������q�r�q���xa��yY+��L�&��@�^�E&�]�2�u:h˰E�RJ*i�ۦF]�"���C�4���j��@:t�FP���?_�m.O��/w�^�D�cnb2�xap5Y>��5<���i�t�E�����
�C5K�rcF5�"��S	��e��TS�ў�Y��П��ձ���g����X,%��=��L���'� �\��})�����ڡ�6o�i1��̾�d��ն5�3#Һ����[Di��Z~�"��٥SS��d�|U����g�����sV�$V�7��{H��# ���X7��f^)���f6�"�n�D�S���\3��w&�����>NͲ�����X�%�ws��8I1��~���s�.�8M��ȥD5�I
��/c7�D��HlzXy��+�Ҩ<��%�;�V���1�����X��@�m�����"<����G�6�G�-�ɘI|�EcHB�4x�'�*�ݘ�	�"1_(Ue3N�L�KE��Y��55� 9����g;M >�̢�^�I%9�g�pT^p�g�+�B�����:v��P������;A�A��U��$ψq��}���E�P��C�i6R�.%�O��������'׆�ˎ�w[��i{K���e���d2��5�bv�REe��*����o/�U�Y�ϞR�@���?Rܹ�&Ʒ������,�{ъ�����*p��J7R��>HOy?�Y�S�ɔS���Wl��
���Xž7+�z�>2��-<	c��ҟ�69J��s��ٛC�bx����ո|5׍�A���/{P9����=}re�C���i�<�Ԇ��f$��0j�ː38#��8���,Lv�,��: D�/Ş�#-뵾*�x8d݊��2��'L�W�L$��s�f�N��C^������?���l]�I�لZDUߝ��4���F3%nɄI���(��<lf��<���-�[��
�E�I|H��a�Ҟ���X����pC��9@@7�6�C���9L:�C�r�H����!��xf8����N`BI��i��� ș�Z�,?JVY��H�p��gVc��$ i���Ԏ�!�,�"M}f�2S|<D�h�D��̼�����%�����|���ĸ�>8��;�-f�Ս��CV�YSo|/�0�+ʐ�&y����VO�~��2��fl��,�<H� � 	s[+������+1��z�`=�Vu�|�rmg���=P�5|ܸ�L̸T��<~�A/��r��1h�
�k��[I�:(JV=!��3[�͔��f͇�L���\��`�4�F��-(%�L�j�B��K'��"�M��Z����ZV\R�|=�����F���=;H
�����R��1�^��E��3s�j!G���4�n��jć��;�\�M?+ql ������\�.��N�ت�?GBV���ܿX�������maJ�-�
U�N�A��[��C��]�4��`���6�`A��)���LG�rF�$���y�V	3![����{t4 	��X�ԩ�ƽCS��k����.Nj�S���Q4�I�1:i�'~
hׅW�C�RAd�G����2�~����Z�Zd��4���*#`X��Q}ѵ��Z|�@��ٹe��A��-�?"�GP�}��iZ� c�#��L�<,yEU��x2�ahp��G��:�G�.�`�D��y@����3��A�0f��O海��3J"w,���4jwJ-�N��A�^��R<`Or�]R�V��W=�"o)���}�AӨ��}.)H�� ���l �D����>�#PI��ܬ�K�5�k�(�ˑB_�k	��m;�X$���>�	�FM $i�ۨ� ~������*��p疡�-U��l��a�z:�ۇ��N��JQ�A�u�]�^MFHۉ�2��a��������6Q����l�Iٷ��;��$zTe0�=�<f*�����'E�`��AK^E��W�ɥ�����N�z;�/�z�8�o��g3Z�U�h����,�J���gV�Q~�~�1H1YI�w5|�4pm�K�u�ٕ|eIz�+��x��TU*h9ĬlUI�t~�֖"dTc��'� k��#Iׯ&࡙*C���0���V�@���[{��s ��'�I����BN��T�H>��OL$Oe
[�?^��葍�����[����������L�R�N�	oA˼�L�?3H*:Rj���He	OB�Z����������2��v(�@eJ�5άw!�bl�!U��T���6�Q��J5G�#�]ښr�lT`�m�:���}� ;,+�~^��������W��P�t�V���Q�/��N�(�T���[o#Xl+\Lـ�nj�M��		�w׬�W�M��5���b�ftQ���Yu/F��/S�3�%O��J\I��\Jf�I	�u2#���o0�Y�]��:{X��Ծ�H�0�z���b:*ϗT;:��,���wE�ېߖ.:�����O �C��������s�S� [3vA%���N�?�V�/l����3����������r������9�\�]@���L� ou'���\jз��n^�*a�[��f<2K)g��*'e�c�-�c�>�AՒ�6-WR���$;gVI #J\��kU�o�\��� +$*�wô@�K�0��W�ʕ�o�E�*N�%������d����ȃ�&����Z4��]������jhZ�q��=[��3�Fi�'�����[��{�$T��w'�p�Lx�%�:�b��3v�A��'lɞ�=�V�'#܈����) �n e��N�<Җ��%�<Z�\(�SM;!˓T������ ��Hu�O��և���!�y� �lYƽ��*�������9h^DG�,��O1㑯q���{p��sW?�(*j%Di��<>��7w^���OƜ/��b0�NK��8w��!���]��q���G��������3P��ݓ����ik��JY��ʄ��7(���z{?�u��v8F�O�0�������f����U]^�E���d���QG:��A���󼺮�]U�zh9a�����\�K�2U�:��0�����4qS�M;�=ѥnp�+X�F(MP!Xug�t81Z-L�Ż{�<�\N����tP��#�߃�G����NrpQ��uHȽ��)�(�Ʊ��豿A�%}V}����n��/^�?���/�/���J�ԏ���n�ŀ��*�|��9`�">���]�(�j��!f4�&��Y���	�n�f���̆U�����̢����[�U�%'(/��Mf.D���J
v���̎��E��I[d�L�i�9�3�{��.C� C1��:?����A*�
̈튶�&`Юu4�y-`krAXS�Iy�D�3�u�-��SR�w�7xR�gcg���S���@�K0>���4�a"��+w�/θ7|�C��������ʓjE�t�rx�J9��M�}0���<);4�܊@+�9���rծns꺀p,���9&tPsf-Y�^�:��> @R��β-g.��	ShMA�� �Z��&od�i���q��,�:$dk��Vw�z|��o��/���l�rq�xzͬ��c�a~ � �efX0�Ͼ�GY��R
t�	������pO�$Hi�/k&)9��.B:�qsrK[�h��v��dU���97��AW�4����lRGb����y�s�d���]/i��]��gn� ���������K]z�xR�� X�5�:�҈	mS����z?u�>��h>�7yn�;W���M�	~��nS�V��x�����=+ӱ{�j�K�EA��c��.km��V��S����Rd��C�4�Y��H��*F��ZIpO�}�GM���Qb״2�^#|U[җ�"���[�� 9;"E���r��mQ"��h^�?�\ٙ�'r�s���W�A�N(V)'��:�奶�/�}�ow[ӵ�B���$���%��P2�	$�z���T���'���`�CO��'���U�b'��r�6f�3���ub�������<�w�ģB�s*I�O�7�E��.��]���0�Ư�2�����(Ny�q�hc��0��vӎa|�
g�������R5�.!�2\�v>���y|�Ɠ��ِ�:�~TAf��$sRȬ��$'<
����d��\����ə���T�ovg�׆4�s��] Z�c��רs��*9+���+F�g�5J �V
��'m��T	�$Ԇٹ���哘�0.9�<a#Kۨ7��8��|W�dm�=̏T�w˴��6����6%�c���KIC+�r��0��v�ݽG���$���p�M��n�kȒq��{�Mޓ-��@Y�<E���/��>D����]Ȣ�Y��')�~* h��%L��O]�:����`H;(�����a�ޙhr��:y��7�S��˭+an+��_�؟��M�1�pI@��t$mm��C3A5"��M3�$���ѩ�ω�^��pѹ��t�����ͫ�Lcd!	�H+�q�Q�O*�t����l~ph�c��_�+��c��3�2z�$+�MA1oy��S�(�b]![��v�Z2d���a�s�=���ȵ�p���w�M'�n������M����Xm߂5:���ea��]P
�����D��j�]�1T��ok��VI�m$dƌ�';bJ�eb����>���'���.�'����;X@���)���9has�:�.�Rd�<������;��?7��Oc���B�p�.8 �9�Fy��f���]5=�L��Rn��]�O1J	��@�>��<����i�e����!>B��)Y6}�K_%�XA�Wu�ń�&�~e/�q���}�����i�^B�Dh�^����ct��/�rVg��v){�t8���@�3��W��̟�����W��f��)_"XՁKN����gY
OA�^���3b�]�ϴ�Bd�I��HC���ynbW?[J[���G빝j�Q~ 8��l���I�/��v�)ٵr�˲Qh�SGș˯	���*)X�T@�5��1�9^�QR�1Y�7_/���G��A��cj��h���Tz��_����X�M�h�����;�ඖ�пP��8�RWCZ�)��xM�	2Ct�����A^2))�_����;�ۨNS������z�n�a���� U��ww:%��R�s,���4t�� ���Z����u��J-�����_n�l����/=4P-�6�N:�k�	�X��)���ઉ��T9�c7�Q܂�z-�����m��{C3u�u��MK��N����J�k|��`{���^����G�-F���m!�8Je���2d��M(�b��n�{8�DUϺr�˧*�@��$w�HM�v��3�u�
��⧷`�_�&�S��e.Is��Y!��&�y7S�e�������s�y��s�+W�*{@�Wx���"d_�:�@�;YR����G�V�1��yg.]�֑�j�L�_J�]mў��}��?�<Gc\'����(�e��^NL2۾��E��m`�m�t�U���+h~��?��<�g� �k�OS��o<O��6e�l�ο[t^�x�ӈ�9����k۬�M��kX��RX7G�S޺i�^_�[��{awh���������+�o&g��ʥ��#��Ĝ��d�bj�`Y*���s��^uz��1�h�~/Y�K�
�������J�a0�$U:	�Y������L&�t|g�Q���$<D�Q�?��O۫��2N�Ot�Z��R/��v�5���^�vGq;�Y����Ox*0ճQ�&����N˲^ߢ�RFqd�J�)�����'%���yX/�e�~8"�s$��>Z��mhPF������6�����	�Y���!�q?]?�A�W;�]m�r��K?T������p��z��.h/ta���8�1��׫〩cu�����<���	$����������k#�g��{,����q������xe�MN��۾0-JT|�����87/�7���:S�G�Gʘ=����Ul��lv _�Oe@.m��d>�V�@���׫�B�M���[�yB|9s�`��u���#vvfq�i�Z�S~34�$�A�fYt�¨�S]!������� D[Z�r��'�C�C#�It��̫@�ǲ�^7��=ܫ�1��J ��~��k�o���F-ii�9����@\�D�a��V9��.o�j�m\8��"b���X��j���Pay�K�n��A;0f�ӳH�Y߁+�ʨ�F�A+D]A�M��^�������Wk�)�����gdn�S���)jzU0K�*{l;��?>�oPV���H��X�����瘏�v��3��9V$�j����!���p��=
�,᾽��8�l��}�$�$p��A��|xů�?,��}�����.HF�����%�:���S�R(f#+�(X&E��v��m���,R��7��b�'�v(��᩽�:Dd��������@L۞��qإ�O���7�D�J!��`��&�6C$�c�9�6Ǯ���N1�]�V�[q��nĿ�<�>8 �����շ��Mʈ����h�+!��tC?�Va���އ�_
,�+	�r�H�i9�E��85d~6�+�q��s'��՗I���"'vōu��N�m�h�G����DA���*h\��i���LA�4&lT��O��,��/�z����Z\cMp'�|ЍT7J��N�	������#��P=-�Q�7~1*�j{趁�l�?K����܏��YuJ,�ל���J�
aK�No(z��!��x���d�а�K�~�ak�8�W��3L�'�Y=������vV��ˮ4
����(� �躒XlA��j��uK�w)������f�F��$�������Dy��C�|{>��Q)��K�H(]-^v�� �����ݦ���y�ߧ<;ݩ9S�7EWl;a6`|͒�+Țl���
C��N�E�f��VՔB��^b'OUkX��b� (�/��EB|�R�X1z:��!Z�w��b4��߾Q�����n[κ�Y��~��|���k,���C���."��b���0����y�ߖէ��� ̍[�\Ev0�b,��7X�;��N�O���5Ԉ��uf2�$�T�FI�O���(v"�7��U��ocK�Ov�;ı���.���sVF��B:��(�&��@���O����Q$~G��ȍY���?���$������)�����DV1k��O/�TZ�|�.��~7�;�v�=�S��!@�dI�� ��ҀpKW�sR��eb \��M�����99�G�_�l�;Ϛ�d^�V�YQ�7������v>��_�'�?��D���`�q\Āf��ӗyJ֫��B���:�E���)֙+�V�� 6Sځ	K8�Lf������&�=t��D�O<�����~�/9ֱ}T��[X�2�J+m��ɤkWM�� 
���B�2^E���<��5�s>P��Nu���Ӝ<ft��/�,x�ݡ��Fl�W��8!ۧ��j�\#'hd�;��y*:��K��Չ�����ǀƄ��>)G�~>5�ȯ[͝%�������>Be�צ�yS���5�g��P�7nYV��^�x�r�r�Ԋ)����.�?Ʋ���_O��÷� ����1.�l'9�+��'�h�+���W�ѕ��0Y��G���L��ÅYęti�p���a ��V�>ۻjəo�8���Er�I,*q+pM��̰�C�ڇP��v�.��U	�Fhr+=Y1UG[�y�������9�/�X�1�`Z���ܳP�բ������ݛ�_�Z��ԝ@�{Ы�X�@"[����X��c�r�+S�+���ԢڔDp	��}�H�1ch�������"b�
��;��y��,�t�1V�����(�f�fCcڭ��=��w~������h���L�+�Q��^?J�ygb͝;` 8rN�z}���0�^@e�p(��MsD|��`Г��e��@��&�G	⭲���f��Rl�Ⓐ��AV�7;lȺaf0��gz
�|�d�
d,!��cJ&!	��9�O�U�
eq�9����S�������dE�6U�:��㵡;�	��ŭ��^�:MX�?�SF�7�ޥ������t��吵��y���J�6��$1;�y�b'g��j��e��tE~ֈ�`|r��ݘ�N!�\BK'o���"�4`�.찄����{y�L�.�n��|(���f����s?d����X�c�3���"ϓ��/[N�e]x��B@ ��W�;�o)D2p<�Av
��XIm;I��Ua'5��@��kX�T������y>�FLz�*QV�]��glP��A�J��E
�,g@�x�v������X�eQPA
��Ȭ�J�7�f���AHN�P��vrG��0�R|6=�}�a3�޲_t�����"v�X�fGa��XǸ.f�)�ߗV 3��y�^x���YiW x;3�F��w ���VZ���+/`�>~�ʂ�R!3���SgyU���e�2,ap�k�Tʋ2����*��C]8K��!Eۗ/�ʶ-c$�'/��LqUW�S
�/"Kb��U�:�*�3�,�(�>W6�'2�H]��&д��5 v��?��X�5F��H��.��7B?�W��01��j�h]�,���:�"'���q<�;@%�$�@P-��	o���aX*T�s5��Or������!'@N������V���x�PI�Ͷ���=��;����0���M] �]��,�k1I�N�������۰.f�d��g�|B��*��퇽B��D�E79Y��������h�n���k�v$cmX������+��K��O��S�ؽ������y��.����'6����mM��<��+��_�������9�
{ź)�!��2�<5�:l�����{M�	�p�l��!l�<ml�u�QrG��"�{��@$W�Ze�晆 q���uRAOvw����P�\@@�Nԗ&�]��2� �=1J����Qc/��|}{ɐ�//^Or$W m����C���&����dX��)v�M�?鿺���ޙf,T���X1f���1Ǹ�)H��X�quX"E�������2����3���'}��a\A-�V4����\�+I�YƢn� �^꓁d]�0w��n�j��Usҷ�K�I6��.;8%i���{��|���p�$Ks�7/��!��p4����uLV�ȅr�b��Q�gX-x-��W'g��,�!�"^�q���p��|���EC{�db��o�`y��H�U��^iB��ì5�6�$
��?xB.�K����t�܏H`8�V9ѧ/WVv�39����W�h�E��+y๟�O�@q$��l/���H��d7��ĭ��M����(��� �{i��,U(|7��8���O|W�d��\�#�l�m�P�Պo�V��dW2��g�9�hLrڸu�|y���L��d�'�S�Y�R��.~��&Sul#Z��@[pa`%Z2�'H�\p��b�_�T	ZG�U"��MO�Zs�n�K�»�_����G�M�4� �Ê=�ā�c��g�"zu���n
?1(w�p6��O�+�2�R�d=�.�Sp`�t�Z�����\~ĩ2�� �9.���wYPxA�E� p7uE�&w?���]~��-��c�pc�_қ��`�����-���y6>ٽ��L9���x3�w�J�Ϻ�!o*��GHϏA��|A��tSG���=i�=��^Is�'�s��^#.-�Y��+F<�)��_5�Ѓz���'ٛ)�t�+�K{��e��t�����^_��̀�Ę�H�\�v@7�s��ڌAЈ-T��3zi����7�y�B��E���4D^��x��Bv���@]%��'X�x��*ʇլfG���{��{<�v�Acbj�� Z"7���U��@�EO9�0m~��s'�iG�?��WX@��0'ξ�i:�$ń6j�o����f�m��8���|�΅����*5."򡾭�p�-5bl��mi��g��RG$���z��ym�35$4��_%���<`C%jU�Oy8�ށ�V��*�@�j�ˇGn�/)����o�^��u21}1��s-t���wd�3�>���^|e>GR�3�ޱY.��j����{��Zn��b
�N���!��
*�x'�/X����q[����G�w��SZ\�Fϛ �-��&g�`�Hh:���}{ ������	7���w�O:`��X?�84�Fߙc�{��b��f�����L���p�1�������i��h������g�������zN�՗�|t�����c?/O������RP�?Nǖ��!��|��zx����d�*~ZE#�������
O�e[�_��o����@H�5i �CKG�M�O;���oB��b�:����}�nC�O$�G�/?�+v��ϱ�:c~mVBF�8X>fp�2.-s�v�54���(�۱���
�i��~
1/�B��g�G��B\r�[�j�����=v��������^�~����'̱\|�P��c+��*����~D����ვ�}a=�C�3�b
��2��z
�P1Bd�\���ُouQâ��;�����"=��m"�,$M��9R����}'�ϋݶ��{cO]���1�QT�7��+�7�����R'F7~h��;�F���ULu�S�Or�a#����*.�9R�Vx��o���n?���`�$"��s�m�U�hn��&�ɖ�/�>E�׵��h�Ь6����\���� F��e�~��[���g�](�~�����Z;c�`��������*|9+w��<W���,*��є�+���<���������±��բ'�ӳ\+r�u5�?a� �p?m��m;�g��T���-]:�?~���T�3�WB��Bh�N�w��ˋ������2,+���=v%nݱ�������x�s��57����$Y\Qa>G�&����[��v���r��.şK�0mCku��Y9��L�#8��]$$͘p� F�6�QN��1<
n?+�k���;xhO�PUs�Uxb�"HT���g1!a�o��".'0��}\�@��f_h����o��Y�<���j����#:�}��ɱ���G4_˙>\��8��v�>6��6�T}n0�c ;KOa�ےnRćX	�C.A+�3��M��=�]�A�iL��Ԃ"��%)�z�^4f�!\sNH<��m����G�yF8D綽5ǽֆ#8������ �qG�㵥�f����ܒ�-oʖ�	��`��|��1����7��������%+䎩��G;u"��i^�{�ɁZmU� ��a1F�tG���E�@|�&.���RI"�{j�����o����j���Έ��N d�7�3������]�ju���B�.����P�D�	���揥ST)�\ɨ/��Yv?�#O:�=<�EǞl:'�Ρyݥ8N����j�+�v�]Vw����2����)p����sP��Y2���{�{�3;�8�>��a���v��-��������' ���f~��'e�ͪj��������]G�G��Î�����s�5�����ʚN�][邙������7�O�lv�ŋ���35�5�J�	��.�C̣�53~aT�k�v�"5z:�h5i�����)�*���_�1F}�U�eӍA�8r�a�7��j������K����%H=N�2N�abP_���zM����ʮ��UJk�[�&Q��&[ލa���[cx��c�+`����/��"�����72���t�XR����k^��A�"*������]d�J�����R�x�9`��x�f[T|�W�B�b��ɭ\1WC�N�����������GE��tCq�ϸ7���q���;�f5�.E�	��:o�}�� -�,{���l9���n�M��@�F9$DTzt��:}��]+j��A �+<���I�I�������#��v
,��jD5;�i,q}DE�y?�S.2�sf�e�h�?Ѓ^{�4a�d��떗p�]�������V���M$~l�߸��UQp�����b���fc駑���Գw f��Hu;@���Ls��i��㛽X�X�rZ�\�̖�ݓ�O��/�El�{+�\A#㩡�T}��qLe=��5ҔwR�����^��q��e֌lL �Q1lyK��~����l%`jP��J5MZ���m���:�!��&��ZtHQXL�7��.�e�T,a5�*�$jlu����.p�O�&Nwn��C���c���\:�Wo�`hrʚ7?�A��0�M�ADѣ�bW?f(P������]\�����V�sf��>N`�z��1���+�<l�56���r^�`���+�ȬTA�%�P�tq3k���眦�vu	��dg
���B���m�{d�,"���1�"�H�P��������^Ts�f���1�XIp�;�#�e�t�r#V�oM2y^��ɜ[7���,�ٖr���/�쓥7�w��3�S��_�}�сmE���l@�<��� ���8��"�� �cR\W8bua�z��-��]�psbĿPm#}�2�,�d
�W�_�ڽ?�ۋ�W��)s�H��+�,��W�1Z�"kSg$���:��
E��b���}����v]����q	xd7�����{���<g)���*��`*:J�D�\���9����V6��]����/����"{^�����k}�Ko�|�����^+\��G�@�)L�F�J��^�o�r��Y����V"C�{��w4mˉ��[�ח������^�A�׌
�.?^�����H>|�J-�@���o�P���)ⳍ�x��l�{��=ᗬ���z�K@Bm@�+�����$"�sVjx$��'14�[�1@A3Z�ω�8�Rn�pz��[��5�����ݠ4ƙa!����c�I�>�1�&~/S����@\�ӝ=h��+�	E��M?���xp̡E!c�~ 2XI�"�,�Tl��q�Ne�NVR9-A�D����$!�Bj�6$��̈́��W(��Ո�J�)�^"��W�o�-�6��kR��>!:Z���0+=b��4�$1�F��]���Rg@����E�'���؆����P�4�&�K�c�JK�o6�}Oӗ�	�u�B�	��兰�a���6�=��.���ӯ���p�����i؀
}�?l>	���Z<^�h.x��h-�M�+i*��7�M�.ܒ/"�͌�w�D&�p��)w�-�$3���8�f���^��� ZXt�\�#P�$��OEfi�I5K	ܙz����u��5�g�b��a��>�Nc�15�W�(��Q��\H�T
Y��@Y�s0�*mKw���U���k5�.����`��QT���|1[ҍ��S��A�u��|���G��a�NS�8E�H&�R�`ó�B ,P f^��v%]SU�9}c0#"�#-����}��P���2`�"$~
Ht�P�D�R㡛)��L�����y}�Ŀ�9$�/XRv�˂?=��96�#��g���D/(�x�n/$缵4�B"g�kM{��>��FZ��:�g��s#o)�K���zϣ:ڲka�zw��>Y�뀍hlAЅf��l'm�>�����	��Z���N��->�@�QO��`܃� ���ߠ��?�A;k��F���@zJcNap�.��S/S��ӼK�!��p�h %͕r�)R���0st�j<��V:3�g�M,��%e�ZJs��7@"*��N���c7�ͤVZ�w|I�Q�+�Ԯ�*	�[�O�篥p ��������������d�H͚��T  ��A����? �P*�"+�,^NA=���hM})m[iWAs��D"��U	�2��B%� �@�����@+6��0QPCr����\��Va闯X]�:�}��r�^�۝��h�bY~�v� q~�2���o�d-�ʯt*;��ǰ�.*U��'%�p+�/}�Zv�u�
5�S��5ߜ2��⢽�S��_s��UJW�^~�E�v[}�+8V���	��*	�߀08E��W�d_޺^F�,�
Q���X�j Jޛb��wj���<��.�=
���b(����~��1Jx�q\{��k^���qn����O���m�e��r-�Hx��T�Q�NM2��������%mh��`ߟ2H� Je��(
�T� #4��á�7���'��#�^�nN�̂�3jE{p?a�֦H���/���������m?��ܱ�qG��Y^do@��Ҋt��K͊��D�`r�� &�sUzȎ��ӣ.SM}|��u�#^��?(e��	�=9(=ٕd��ۼ�IŝKO�^���Rh��O&hX�~4$v��K�Q��8��k�go5��1�S�5�6��+���������>_�-���M!s���N�������A��xtg))%BB�؇�rUN8�E9��\� �֪��7�ٵy��u�W_����O�05�O��+�l-A$�g�2���k�2���E��31\��a���	c�o���a�RX��`�A��m�!�g۱V0�s����ܟ���y�4]�an�5�;��xMxّ�h~����Dعh�e��#�;`����������e��(����7��ly�m�B�lŗJ��=Y9��{u�>���Yg��q�M���c����la[�L�;��L�
�`'[�vC2.���O���)��Iǆ�\#�A��^:�c�� sݾg��΍�M�.e�~X�0��-��k�u�_�,^Rw���8�a��q���A(��Q�Y��������1�g��Z�%�n�:�0����������sB!����0�[���&�:��u�j[3�x<��ۆ�ق�G([S�b�, `��M���C$>x2�pv���}�͸����Œ>	մ��W������M�+���.���I*�9�Ĵ"�Dh�h�Wa};4�|����U�^�7�΀4��opx�E�T���o�Q)D���y�1�Sc���:.��5��>���:;(�*u���[~�e��wt�^��%W�`�)�4� W���iM��7'%:��LЬ��ݟ˻1���2�~�fR����a���e��<6�n�:hp���$���K�#��Zӄ2�fv�Ȃ�Ӱ�B�ǵ�H���s	b�)�����`�șKx�:��e>=�l�s�F����ڱ�QBo�ڍ���׳�,��O����+�֓��;AK����x@�B*�G�C?���[�'���_��,7Qj�,��}>�?�:��ۮ,��P?B�q7���l;���?@N�z*@_G	�M6`ɯ(�^1�&�k��0��Ë���s�Ox�3���!+��ʖ�T*mo�ۥX�ϴ��W�
����9���LO~<�}{�\��Ȣ�����rE
��h�[׸	N�&��+�zv��B��tZ� F�����҆te�M���7.q�hǲ�7�>�M\?w"�W��徳����YN�K��;�}�S�E�����&��9���Z��K{�ID�� f ԹSWXc��56ٕ(?�qb�O�q9 �!�*��J^��>'Z���u��Ưt�X| ���,�?�c���R,�&�J��9���]4-�����0|�b�	�~��%P5��A�,�ɿ������d����AYP�*�(0n"���[��$�W,�p�q�9_U���̻�>�*f<�����t���nIW�ι��K�}�h�O�!���h��w�s{C�Ak �}0S8]V��u�������5���3��cx���
��e��k>���2K���ϔ�T�� .���hZ���@av�4Ɓ�:�Hy�NBˉG7��e����;�C���:��1]D��*�uP���(P|6.����l�)��/!sc�1n������Դ��k!�Af��)��n�X{,�He� �WE�0�mw(��I���Y�Wd'\tUdhi8��� �riGu?�|4K"8��x��\������S�irA������ �_��1�L�UAa��
>��l��U�
���U�E��k9,�>ښw���A�0�h��#����(�k<������Lg.u��s��n��҆�T%�T٣)"�U>'9���V�uF� ����4�����;#��
�-u3
��ޜ�U���G��>Kb���?3�J�Oe4^�d7}�ZE�g��j[�����-�ܭ̻g(�l	r	�A���ʐ%�_}�#�?�;Up�9{��LJ@����&��C��^�:A�Z��	?1e��<){Aۢ���6�e��t��$��^Oz�YZ8x�#T\5A�y�K;?���p����4G�{�քxPR�]66��P6*��k��ت(EA�.��"D;v�h}���Q���dgQ������Ao�C�G�D,����~�m�ce�R�&��zGq#��3|�q��d�fL��i~|�,�s���|��u��Շ+m3A`�r��=o�׵�6�3/��69{�;u	kg� l?igמ�/��u��A@���s��`�[��Y�Om�ٍz�ͳJ�������ek-Q��҈�ӏ����0�����Q�����W��\ѲnA��R��m�|��a�˟c�^?��QV*��M_�ˏS���%��.��`&���zny�����vHpY���{ne�k�y2�L�*������ǋZ�ſ�/9csK� D�5'z��d�{��l���q95������+�mA���(�镵F÷D�k8�왿;L��3㤜qO���y ��D�Q3W�ǣ�{~J-0��������t�QM�SU�q�*ոS^�����{gX�VTsb��eA�RUf��!9g!\~m���}�RF��IYŰǘ�ēf��dѽ���j�)���y�6}�m=��F�l�Mf����}�)ݹ}l��؋���a\(]*J��C��?x���_�/��g�Ab@T��������nC�V�aX�F��@@����@T����T�Zv"��'k��\Q� ^�G (rͦ�MlXMş�Nd�2�&���d�éL����Yu���c����kf&(M'cM���`}B�1�
�D*�n�D���Con�c1�������%v�e�ᤪQ(,�(p���u��Bۚ7�5S?B���s��g�)�^���#mh�4mo3� $3�2��I(ոՖ�b�`نL@����w��	@�XO��B���:���ʊ&��'�.{!�	��u8r�)�Lk	'�p���ǳ�Qp���7+F/������s˶31�U7�����♆VAK	Ce�Z1������e�Zϲ�ځݟ��[7��WXV U�iJ�ۖ͝�I2{60=��+�Vs�\e˰�dcgk�c��bE���	�,�3�jU ��0�ށ�g缒p<���ĝH�Izo%Čnx��f��ɇ�ћުp���l�2S�wl	,-E(`^�eT�>]5�x|¨��&uA!\�C���p��50o|wh.�����yn�W=rq�|0�!N�����SVw��?��%@������!/��.��ߋ>���EHt�?nd��IF���_N7�H@�/J�K�E�v����>����K�;�yڼ���
�9��>�z�ˣc�c�;Y,�8'rl����1�"��+����u:{�r�i� M|v����%��7�r�R@��X/�Hg�Հ�&A�ޘ۱#
ƀ����]�C�.��)����ȸ�����1�c��d�\a�~�#D�o1��GPփ������^��S[��O�GAWج����>`?f��vC
OLO�=kM�>>̽ޮ��I�+�H1Bt՜G�����Lm^�MD���=�kp���� lъ��C���w��+�Aܼ�-I��Μ��VDᗙ����"��
�k3�ςjF�F��֍54�,��{���i�BO���̱���u;χH�ׅEh�kh ��}�/�8!Y��/r &�p����\R�l�:!Ő�ý��6W*� �A}�'aA�[�n��=>/ف���㝍%1zPM?�5Fy����~�.���9����`cu�Gy�4);����E8�j�4���!Y�E?��c�����z��(�U �f#u�ȩ�dۄ����e�_0��h�c����!A�8VU��T���"�ccY!7�?"�?��=p>H��.j��{���=�j�/���hl���`�C\�&��W}:C�%���oV��2�I[�3�ܛO��Ai�P{ŊCo�NF��ZzZ�$�wE�����v@ ��-�!�n�eH&Q N��H9^j��C�:�-�e�R !�/֗��.S�;d3�A����Ԁ�}6���@CJsڏ%]3�SL,��?H��0-��~�(w,T���PW2c%��%��8����E�id�$�V��T�,?F�H���@�嗥���7�)��t���#�ph�Æ�j�j߉|�b)����T����J$3�u�w�ΰ(8�5��<�7�Q�����ED=v�&����K�[�}�h�Qg��r�K��%6��)lob&��0�
q2���'�OA�OKQo:�(��ST̅��� �C~�Ş	���zdX��b��$�4L�U��Aψ ��c��;e.�/OY�̿e��ˉ#P��ޥ>���g)r���_�� �[%'ʫ޿�/u]0Hثk4n5^р;�!�]��6|R���F����H9���{���K�6 �8!�?^�N|<��d(6�A	���T��$D=��B�q�@������{N`�"qKj߂B�P��������~q	Շk+��QB�2nd�\��O���SJ����"��P+�kv+��Ig@D�>�HU�Z�ݒ��E�tt�w�*�� �O��zs/�Ӷ�ɨ�К�Wyܳ�d���T�E��z�+�<$�-�&��(.{7���veJ�Of��5(G�CU�R��F^o2M��K�-�şs}��+�cD2��G��wr���:#���N��nќ���`(LK����r�Qg�	ɣ�C��|����3)U�yl���Sm^���`0Q�B�O�p�Ŧ?T�]�v�2,�?^�񟽬,4��{�QZE�&2Q���mK'q�I,�����9�N����ŷ8C
�c<�C*��V�����;��܁h��p�s��M���T������k���t����腇:�v�51���}��h��N��j)�Ao�1�hU�)k�kDK%5���mu^Ǝ����M�Ն�ŕ"���Ў+CQ�d~�Rg�������-f`�$
��� �Ƿ�.)c�Ԉj�D��Θ,e���ZR�?���*7��D�CQW��)-�	ȥ��g+�r�S�l�Pl��ul��4?Wk����S�^��4�N�5�	w�����R�c�p�s� *b+8IB[�Ф���K���^p7�z���&�?������9�߽(T.{tM�;�
:���R�#Dxa�f\�^�g�z�Vj�D��7y�ۭy��E}��p7{����6��	�*Z������8ם#�XtV��CV�ɗ������:���'�b.D,��pRc�G���y�F�!���2qx�� 4ӥbE��~O�vK�4<i�Hp��o�n�!ɎN)�O��D"�G3"�'�0��VS���1=���>�N�u�_?6�p��nb�vm��]e�x�nz�I[͟P��½dQ��[o�U�9u(�{�e��qt�j��lm7GS�8lRC�{����B�Ff�4�.����jQ�i.qcרx�{��J(�9���l�#�g�����B�5lj{��j�Ѓ�aw��Y���@�1�)�EĪ��<�c����ZEv}&��u�Jg��c���nިz�_�65��:
v�sB�d���H��B�I];9���4���@��y�u��T�����N�G��.	��H0� :��]-�e��/h�$�"�%B�r���Q�� �E<{�z��TQ��`�ty�cM/�u���ώlq?r��S3���.a7��i�fU�dA["@�~`�f���U!�c���\!`�&=\�{�O�%G�(L;ܐ���Ș:E+��A��ofn�a�4�����*l�m2j�p�kh�
z�Лnp��g��� `��R)�0��\�QZA?����F��OSv��ò({��}����ӵq�#r�;�^�@c�����FY��J�P�8GTM��D�����s��]�l���BGtA>��f
 $���W�_�p �L���nY*�@ G�v���+'M��{	;���: gk�0QX���J�t���"��2���M��I|G��Z��]Ha-׋�6�8A�s�|�G&PD�(���og�fh�-9'���8|�E T��w����LQ$�L�sca찜�	Q��ԍ'-G�|G&	���ْ�ë��؁����X���oS�^���|&��)�ҋ	��Dw��URlH.�%��]�[D<��kn���Ɗ���!a�97]�.������wRc��P/:�8�	�����,�Й1g��6G��G�����>���B�J�V�~��Ļk@ce�9B*����ab��2�@!
N*^۷�K��/�;�h:��5���ϼMߊ�6��=?(���PI�?�*6��n�u�����
i���N!�0��[�Z��r�W+���2O���}�����秵|��dK-#%�9���k�*+i�#�[i���t�*�0n[��YG&Џ���萏n9/�j��o�w���l3�'u6b�wmQ*8�$�s�.j�l��L���<��o7F<������}�e��
�W��l2��`ߚ�7^QF�����Ւ,�w:��6�f�נ,���� é��4�Ǉ���}��~|��u�F<+�t����غlh��.) $rѶ�LnO���ј{�/Y��� �i�� U|�6�>��&G���@`����d�l�B��֮^N�㲰T�k���)����]v�G����G��"��3G��9�o{X�� Y�?��E婂�wQJ���©�'�C�L�{��݁"+�?�^�F�hb�5�>�`=�1O合�����7��)���׆�����W�3��~�g��`FD綦�I�ߧ�B�n#��z,|�^r�"� 1��eri������Q��k������ڳ ��L��7�8u�+���c��V��� �x���
�ܦA�������#(m���Hi� ���)��<hq�/0�Qo��~�$y��0([�!�r���W����\G] (|/�5�5DR�65�k0+�N�[�B�)��R������i�V ᅕo�R}�µ������Ҹ&�E�6T�I�'��E�Ab���\(r*��^fj�#�J�<�_���?�y�;J�I-c�bi32/ +TWD��w�T.^��ɔ2��ӂB���˫������p�Ľ�rO� :=!�[���.r^����J�s�h�1t�6t�|,Y��ezТ����/��{0"ܙu���B��Ɨ�GF|��1��&ʇ�EnN�Xf�GR�m\�Řw�PX�)2���{�JЫȺk��m���
���C'�o�s��D�f��n����*��3E���]��:�?�:�WZpmQ�V�w��!'�ڼҿ�Of�8�c'Y�1�)�RP��lz���˪�w��TWϙS��R�ek�O!���mw�޷Iҳ��_�
Y������\�u4�|�x�[{{si��8�à}�c�U�B����� �dVSk{�K���9�Q
�9�KV|+1$/���� kLҨ[�D��I�u�bQU��� �c]�*d�-�NܸFڟ��������D��:p��R;���@�X�*Z#�fe��m�#5��P�|F^3��j�5[=�mE���� 2�6X��4�7Ɨ�t��o����B�Er�����-Z�|y�x>Z��'>�uڝ��-�lJ��qn��͢W����k�|����a$]lmAHA�����b�k����B�ð���\K��}R$[�>�,�E��{P߹C`p�v��_d�����D�a/#<�� и��1 ����|A\�CD�럙�!'�&�X��˥O�����~6>����[�.�,��;��ڐ�>p�zR��?��Ӣ_���A�b�$�l\?��� �#�n�p�B��'#l
DAȺA��H�C���3?j��˅��n�N�s��Y���q�Kx:ALE�YP[�0Z.�	��F⧿*��n)/2����z ��Ki�׳�Jr��6�(B5� 8��rY%1���Kj�bTrc��������$���at:�F���Sy����5%��+ȘR�_��
��|:�2�XĦʺ__Ͳ�tK��D�����Q�chˁ���j%oh��萗B�[�K��Y[�����{��E�!,-{��U���+�/l0;F�b�&kC.T\D�$X[AVU��W���%l~�Hb��$��ٚg^w���p�<��$�is���a`�r�y�+>g��j�'zE�����E�?F�KCa@���n\�a��1��m�����b3	���G\$hIL�q���hn���DkO�煎}�+b;�d�K�$�������Y��U�G��i��Oo|5j�77(P�*$�/W��cx_����r	_8���#��c�\�)���@�mX��`��0V�����ڢ%������P^ա�$��n����i��7z{y��|�H�V��������h%�!2�_�[d>����y��FGg.�`ͳm��[�[Z
˦A:e����!Z���"p��죯��z��Vx�<�z%E;���ɫ+�(bwSHau�j8����b���>�&|����!Je�@2k%h��+:�ß-�V���Ř_m j1�x��վ����S|���i׌����^�NJ���O 2�>���Qu���b�΁���@�@S�! ��I�}��@�$,k�_O�Kg����k+���,�D�خ����U&5�M�|~:�P;���Q���������j��V��W`���X��6A�HU.���c3�5]��
>��p�0�9)e��` ��p4y����x��_t����G��^��خ�^6_��dz}.��/�yx������� f�%���'��5�B�5���,]�"=]W,��G`���6%���wt����JWl��gm1��{ۏ`�U�A]�{�'����k��M�e j��R�R��o̧�ܝ������Ζk O���+�z���Y/..p�g�4��NYa����0���nu�m���sR(�J�]�U]#�g�K�Z���I|��ݡ� D#�Z����r�**�n�$�,�x�!�r�d*䴆��hU庙����w�g
 ʙF��|<��>Ί'���xt%7Pnxў�'i��������R��<]�?�X��l����]^���yh$3>�̹R���}���7hڃ��]$B�x>�,�vZ�!<*�:dr�n՝�	*H}�ً3B��+��b"�MT���&8_������7]��QSC:٣�)��]pf4`�Wfb��4�KYnSU�pp ���
W���L6�Z����b��[n��6$���[n��l,vJe=Ez؝����jj�j��I�x�o���#Q�����B�#f�`��b�f�P�V,�6��6�e<�=�� ����q��|�����^@&��y����X���	=6dx�����[�	n�U#I�}� �`lz&^��Ɵ��`Ֆ���g�L��_c9ƍ���$����}~�H&�+�.��I��o��D�{���Q��9.Pڢ���אr�����-9�O2}>�/�3�,�ښb3Y�u��@���^�j�v[/-���d�(K���a� cX$�eA��Ŏ�
/��hb���p��v��k�|����8�X�ys�
��6�\�6Ts0��@y����ViP��g�}]����P�3R�r|GKVrr��<�JZ��9�F.���E	sL���a�<f��f�n"?ܿɿ��ۯ���K�D��X�:��vV&�
��d�M���Y����7��Y��Phb����Ъ����{�r�%�4�?Z���w�����σi�p�����M����`j�K ��+,љ
.���bi�o�e<Y;����o����G�Z;�\�(ߝ�V)V�\��������m�#��?d�;uΧ.�� "w�'��m��6�σ�f�<ȝ���Y?���[���)i|~b��4�ؓ'�;��~��}w�.��i�@�.�Sǈ�B�_;\C`��]�K�J7Q��hq@ɖhxc�~7KJ����J���ȿY�S����?]Ǽ���k��w2�d��z�� �J�e7_7 �L�j�Q���.⽩߽v�.<��4����Ք�*�A4]�A/�ד�������X�r��m_@�;���~�R��	Z��<^^
v4�(p�@0SU�.��U���Q@�	@7cQܞ����¬x��"sU��Gb���Cw#�U{����6��&AK��s����z�}���&ϋkU����a�Hl��{ԥ�QR���K����u��K�x ��Hw��������Uz�������u��.y���~V��~5J�7+�v�$�/v�3����mv�00T`�}��m(f)
�9
ap�S�X�aV`o��a�"��$�p-�޲�ļÍ�����x�QC������Ӵ���X�.C8W%)�c�V;�Eap迕Ď�.�񕜴��@�t=��<�@l]��W�do��s6�%�W a�w[�ml[��� r������{�V�8�6�����iBE�NJ���k�B�u�~{�Ѐ��'�a���I��*E��/kt+��0���ZHE�+WM�,�b(��a��Q�� ^Ei��{1�c�:\���N�cA��+ ?D��:v �r�հ�\j6����P�-C��z�(o��;�#�فb[�UJ˻�_�c�,�|��r��b:�SS�29o1�/��[�m�v���=��!�҅�-�&<ݪц�8�Yj�k>$�h;0%�L���D��:����޺B;���
�X��TfB��R�R�*�jn׆��\ߥn�!+�eM|���G���B���X��~�R��.F�3�ߎs��2���n��~����(�
w��Y�O��)t����Ͱ��N(��p1nH~����I�,T��$&�4�_��c�尌:��߾hPf-����hR�+�j�Y?��s�V=����,!�;�X�_	"=eA��C�����Y7�&��~P"jaa@N\���Z�N��<֓��d��L�k�Ի�v =�g�����0�W<,�˽����G���F$̇*��"2]��@xeς�	Y�*=-U}$V?%���smɔ2{�;�A>�A�:����J��|F��ߏ��D��HXo����=����1��H^����+aZ��/�EG�`�l-&��S\�<n[�Kĭ���[D�v	~�D�1!�zVk��gs�h��%���J����j�����F�������P^�����;:1�h�f5eݞ��q�t�����V^6�R}N�h
#I���-,�Y��Zm���\_�ALj�R���716�9A��Km��䬆�on/r�lÕX���r�V|c*�1H���O��%iW��[�,�P�Q���Ǟ	Vպ�C�&�S���cH�C���?��֖�5�(��$M`��M\q��z��
��)eۇc�0�:���t����EZ��@��<xi��ù�g����KR9oY&U�{ˣ=a6z?�|�^#��m�t���^ҟlv4OW̬��i6�.~YL���vqntF�c�e�};�����3n�J�laVi��Fm�=��&�h��y�e��^.�#S�gK*��Ii��jN�vy���������R&���R�XAe1�4q���1j�;���
r�݊���;	��c�8-�8����_Vk3�v__���GeI��:���90���}HLs��(�(�>�FK�M� ҐH�P:��z1;QŘwTtb�$����tf.�5��@��͐��i���/�c���s켝�k1��_
�iE1Brې�s�+�nR2����i��/��m�u��������	D!���*d�.��f��䷳��v�&�ړ\��qF�Bi����oe�=/�S3?��f�^���x ��j���'�Q�m>q�Oj�H�h��%�4\x�Z/�.%���06g�Z��.c�r�޽@���(ޥ.$�J��Wďܹ�w�v�p5�Fe�rR���mG˞����jW�E�{�2�O��~|�������|:6�@b�#7greB9@�"WZ�&���x@xS�P�9Y�/5���@���ć�>�Ev�e(����<u�S�$������˦��_��I-@w��ɂ��
�Ĉ�C���@��ca��H}*��lzAb�@���YQ�L���a%��>�׫��$ò�[jW/K-�<��cA��'*�����#.�\ǀ3	��'�z���-x�j]I���]Ǡi��~��Md��<0]�;���g ���D�sm�2�I�ˉZ"$�k�"�4�]��h��8c"���2����Kd�'t#L�r ��U��a�hv�
�?�A�����qzP��w5�*��Xl�WH�;O��U��	k~Ln;�^:{�Dr(���S�Y�v娭�R�f�QW$���v�"�]�j�Z��!BMY -V�(Spt�7�g:�j�V�	�M��=�){l�@��Y���y5A�d�� ��h\�Z
�e��w��@D��hPD�oj�o3���2B��!D�����-(���jב�k�m\�֎= �7J~ �H�������P��TZ��m!A���#7�f�N�p�s���i���ŧ�3��h;]H�ފz��Ҝ/%?�M?��������+.uw���>���E�ͣ4J�����,Z+���H#�i�4�^-I)\�r�I�
��qTc1	���d�i�ۅH8&e�	�mϡ2<����A��,Ke=u7�{MX��P�\�?�U�H���O�4u�f@-�LF�;�MB��
rz$�����v��2juoK���c�D�	´f�S������w|���t3h�0^��t	5�$�(X�	Σ]�S8�{�A�&�z��aA�:�x���,`6K����_;Q7
��L*].�2���(�n6��b��W>	�FM��F��H
}���0J�oL��u��x>�����uF�D���X����N��J�`-�6ኄ�
����Dh���W(9kW�ZЇfgT%&I�����V� ��|Kkb�F'�5'�̐��7�lk�f�MF4�t��&�ż�{���+K�=rn)�~����Y/���+Y�(�%Zy��#��kn�=� ���<�2�w�4f��Ew�̈́��^�x�uf�%��V�H}�I7]�� �ޞ�3�%FA�Oɦ��H����8��fg�����)IFi��/=��C�h��:k}��!�\}"�V�K�`�Ȣ�����AQr�_����.���h��m7�2��}�}��9ѿ}aj<.I\��;^!��C�1��8����K��l�f�-q$|�dpmbsB�w���x�;"j�m���7�&lz��<��>ދZ8Uc�n
�~X3v& �;X�@�b��$���r<[�2�8���i�����ǃ�D�P"��N�UY�y�fp�tڊ�������h>&وeS}�^��/o*:���+[��h8l��ד�"��:As;����8��/B�)��✹�K�i�r�wX�o��t4m�	������K3r ˊ�A�4s��5zf
}<}"1P6OѠ�D`?s��	;0�]�$�i¾{��0@��X�
�=��)03����x��ڸ���RQd7�wo�P~��vpPj�Tn�'3���S�w���]�C�9I0��n}�ˊ�i<�m-i?�סf�aAʁ�B����)w�U���I�K��!>f��j[��X-��I�ɯ�a�(˚^,m35x�I�{�"��o���x��wdf��K6�u���<�i(j�·+���l[��ɘv�S=����P�� +Z$f��F�FB�=q �[̸��I�����lk-z������DBCZ�`cMb���M4Bﲔ����ŝг���]�R'�eGp�A)u�8�O�db;]�4��C����U4:Q2�Ai��4���z�z�v-�5H�)�~��By5��w��v��Ʈ\�X�Έ���(�,��}1{ώ_�x�����})������|�fd⒳��[�O�L�Z�nHm��H�}N�hG �l������x��/� ��H\�'��B����Wݸɐ�=E�}��F�F�8 (�#/ڣ�1e��#u_W�$�,JS���r��[x ��(��G�.�_%���T��#+ �d7t�_B��;s���e�l��7���.Ʀ͐���L�bD=1+��#��Z���Rs�_w,�H����N�t����-��Z����{ dJU�Xd�q��9ߠ���ًw��@��F�i�n�s�y}����t�*��YtH#�
L�w��B��y�V~��G��$�0�Qfx-�PωQ2��Ϲğ�G}�<�IV�|�v,$�}�؂�$R1��N)�XC��&y������?�
�4���N[����7�g�sj�]��$�}��Ͳ歷�P�>�����.��v�]��E~�in/�a�=��R��Ŵ($�O��&Za�<�g����T��K�����\A�� ^ �SF�p�&.?�ad⒢8g�̃���e��$O��u�<	�ǫq��j��@�d$�t�jv$���Q��a8��1Xv��!"U �Qh>��
�j0Z%ۡ�L>ѳ�!C��K���i�����%ۣ�b�V7O
{�Iw���E���Z��f�������Nf��z����l:| Q�WJ���lr���R��yѺ+����W�q���P�H�Qm�]�(�2湮�)���2��!d۲�@�%�����y�XmfEC���l���`�(3N>�<��+BQ}|��Y�ӣ�>�Ӗt~�_E]eh�/���kx�e� $��"	S67�L����dUں�~���/F��dwǅ7��+�<�Q�5a�JD=�������'�¯/��&�-WEou�2V}����xMc�?�2T�M�*%�\�˾0�G�a��6Z��ox�J��]��j�C+�ؽ�NC޾)_�6* ���%LnA�e����z���(
JEiXi�2\�}"�6di�:Tw�&����\����8�Lm�M�!)�ӊ�@�WD��W��_w�d_�?-��O"�x�:��O�Ḵi�lN���x\:�l�^�C�0�ku	b�\ƅ֔8���Cp��h8�Dhu�s�(���zp��X]Fm���;˛�r|#s��*��M*w���"�FW��0%�v`�]x�k�cv�n��4�8`55#�rj|�&R����}�I�į�ߠ�u��]7�J�Z@뽵��Y4Y.2d��<�-3|�b`��&^�3�v����Z߳�+p�V�.�����E-�� ���.���H��X�@8��*����S(�[�Zo��'���I*ŧ$U�V#�/�7&n+�j��5�K4�K,ī�mud���d�ǝkq�^ɕ��H)��U��Zqi@ژ��30c,Xp������[P�(݂�To�yD�������0P� �weÂ���f�qFmy9�\A�|&�c�Q�I�I�I[�bp�T�5Q�ۣ��PX�K$��h�Qm~�u٢�%]�*@0H�K��{�)82=�{G��0ס�~/#-�-kn�L�~T_����J��@����A��,q�?����k�S�}�>�����Ѭ��������(uK8�.}���|C
0q)[~t�hB�Ҹ��)!���9ɤ;��dT�L�}d�#�@"/����_k�?)�\��
z!�N��h]�.F���"�WM
�����]�&5Nc �3k�lM�oIԥpԼ�D��:�&�l9O?H��oH:�/ސ�8���v���^ۊ�E��z��1��Rwil��:ԕ2��H�_���D�y�D��-;�6���:;��t���/i�v�\���"-���O�MN���`R��X�`���
����:�I���~3��
�f� ��e#��lQ����1$H *�@�A���(߹�Bu�:~�LOjŲ5U���.nަ�w3�*~�7�Bo�7@;��2ĭ�V�oGJ\)�_sX+r�Ѳm����>�\D��+X�hJ~hc��-#����o5d��[���
��k�p�J^���?�IzG�OPB�m��e8�ō�S��?�*qwp�Ȕ��|Pw���tS�;\+�qT: �*P�8��a��\�.�ɺ���S�]���K`�� ~k��Z�.:.\�A��R��	K����k����h���Ћ5T{���C��w�*�'��P�f��+G�^�z���厔W�� 4�Y:k`;���\/�T3:u�э������q5����0��A���(��5
J��=d��^����C#p�E0P�W�Aq��k�ߎ0��+P[�;������-Ӂ1����>�7n��8i��'g�5�7�P똱�L�s�M�~����;*ZT��,���Wc�\����l�%��=�I��q�*>�֦�Y�5����5r̄�f�eɅ�b.vѝ\�8ӌ�՝��~�j-�Ok��=�JC�����!RR����CDa��(�oޝZ/]��l��m O0�QWo|L�ψi����nM��8��8*����()�750�����=�1O����ywrf�����H�|`O]���I�+e���@�4�5���a*<>DJ?�u�u��g �$>c~c��C�G�
Њ�0��D�cc=P�[�wN�3If�}ey�By6�J�g�)�@vB�N������\�΍��4�?x"�S����7{��X�!���`8>Z���sn�L�
頟��"�=����ͯF($���B�_ֲQӬ��&oө""u�\vբ�6w_�s�uo�ۄ��.9��ehtpM���<�=�zn<� ��ZA�B��Q6��^fvv�#�����^/"uD��(|�=[}�������&���s<�'{�p���$�.P?!�׳} �5�cYO]y!/�J�y�[O��pH��Z��d����/���D�����Ku��w/:�n�dDl�po�i������曜8d�r��~*�i�ra4����-Wb3�=k,��ԛ�2"p�BI�y������ �򞵉�mH��2X���a�p-��<�2�2_�x_�|:o_	W~� �����)E���z>n`�ބ�����$� �28}d9�t�|ju��"�����9�s��cD�Y><`&c�nl	��y2��<���8�;�z��~�;�[~�m�|�"���Qi�>��G,|W���e���	�N �_��-q�J��ȶ|0ܰm^�kg���������#���f���X�B�z��o5�a��:�QX9�f�������%hZ�	92Bj���_�޷"�����ɢL$��Dh��j񸺒�w�#·�CK��`�e?q�T9Su�C�&tAD-<ܺ��{Z\,�=GZGXX�E�,r5�'���ΰ�y;c/�sT �����аHA�$)݁Ϗ����qNB�) ���B��㧮bnX{m���p��e�iξ����#Rn�^C~�dmU��i9��,�&wϛ3iB	RC�9)}�.B �G�*���M�~7YΫ@Ge3l��Y<{�D��}�����q��@�/��0��#H����
ޅcyG�xn/��%��*i;j ��ua���D�W�g`��2�O|��9��i��z�4����V�:��"b��HmrKr+��o}�f(IE:b��;O<�k=��5
�i[y���
�����վ�F9Fs��+/�����;X���ͥ�8�8{�̄F������6��,�=���eή�ByHp��Q^<�%�Zfi%��=�,�O��rJ�g�K/^����9L���l�Zj�#_�[7US�3��P���,�L�w�{����;���9!B��/y�Z��̬y��#������d�������t�E����j0a)7�T~h>��ZC���"K;�5s;7�O�Ԅ�\	�n�����ڐ�1� 
+¦�|���̆i/��e���L���)��B�j+�[C�M����h�����+��P����U[��R�8�j	��;<�����1r��e(�E,dZ�c�	o`8J�ӯg?O�ȓ��F�4׳��M�Ku���щ�R�b��F����fl���7�X_߄��5�<�%6�=�̐���mCG��4[��^և�q-Y�_~���>�2Qp�V���(-ƣ2ms�ճkF�<�vks�S���(/j(ȁ�ۃD�{ŋ�Ń��q�ǚ�~���{��0�>��<� �t���+������D�>`��6Pc�KUY�5)l����%E�,�+ҰQ2�d��}9��}U�*��w��!���Ixh����7�̀�y�*|�:�`�e�Ī�
��̪V�7��!���Ba���l�/7;�&^9<�HDMV* P��'�>V�M��Tpx���pB����?2G�>�R�6�X~�84�Ƿ���� ��3�m(ZI�|�/�_�����3�"����}0|��}��z��?=<�ͻ�)E$�M��}4w�9���ĝE����H�t-[���Xqto�%?hV�s�V��S�|��W�£��.�Z�S)� ��#�5�P,���2C����r���y."'�¿���?]^�y���I�%��Z��Y3�������>4��u�o�eiê�F�t���e<��v6����%�dch'�+Ę����ۘH�2L�Zpl.QX��Og��!�I �R#��'@N��6T�Gď�A����`\��(LW&�!�����r���ߧ�����ܺ����q3?T��� 9�믫��=2�"O�ң����%��������e�V��U�:a5��Aˡ�sts|����5�ӜQ��7?巌{�F���^o 8���1�Q� ��^�h2|��W�3���6yf�x�	�9���9�-3e���c��}02̾�yI�&���oG�_}@�k�qO�Y���C"��v�#���ܧ��_����U�w/��܅�G��o2���׏�dF��!QR������sRJ�ӂD��.���H��D��ݵ�P���d`�ܵMVL�qFm��wL�O�0�Q�G�ʕPT&�ਦMiP�C�͑�lz��V��p�.5v�je��<I���? ]B���� �2�Щ)�u�v�l��p���ZB��6�הT�R{�{���|�{OX[����V�����̅�]8�����|�85ŝk!e���~�Sf����7�p�_eq0y�]ȿ 1��%C �U�ՠ"%�=��w�}�oZz]ܭ |���lԯT>�.ou�R�o^�-�k�Nt�s�k�R�7α��#�B��
�\� )�_{��&0���0��@Q4�Sb\�i_��[���������i8T�}���j|(~��o�G���k<'��Lh��"�^� �`SJ'MΉS2nK��S�Cw���*չ=u?��Z3�HO�A4��BDe�����Od�3S��	3�ٓ��)���0�=�f"%}�|C���V%��$?�(���A���`���y�aZ8T۩8@�^��r�kҧ�e�|�8�A�P�@6R^E��,@r�2�C��`�B]+Q���-�i�H�$�	[PW� LT��pިʈ�q�q��a]q�ՙ�kkZ�Gz�_��2P�v��u�6%��i9X1\�S 8��!E���״\j@?���u��%H��^s��~��-PCU�<ӝ���cR*�m�젲H@i������@�X�5�K��y�	0��<d_��m`���ۨ���D���B�q"8��E��G�n28U$�F#���_��p]w����6���)�V=!�J��vE:�0(5E��ԲP��v�.$ij�c"͢�I�'( Ɖ!*�?`���t�߻���g/6��8qU!	痤լ�I�,��rк�it���/�G�Ƭ���� 4��5���f��w�@��x�,������9�&��|o}j
l��+J5����+ָ_���듛L9��R�@2�_i�4b35Kv�!p�\y\Tg�<��w5�6�Ȁ�2ù�r| �3�U὾x�����pg�A,,���C��cb���lCɽ����봾{��R������\~B�h=���`�Z�A/���L�|-w�3�B��3B��#�Rҵaz��]B;��Pq���
v��h����#�
z���
Q�B��aCV$g�R�Zq��^�~o���X*r���l�ڲ�]��~	�'=�"+����#ua6����H�\	�^�oh��\L-W��]iK�o�>�:2��aP\��yڑ����Be�!��-E$h�q
�N6���Ko����oO*t�&φ����>~�l��Ut�6�5E^�k�3��q��ٞ��ٱDʢ�q7����cLZm"���@��l`k<��Z�-(�����Yd-�@$Ѽ�+஁��Z��`S*r�^�[82�-J�a� �:]G�ؓۙ��Z+a>\��9����Ef?7��H�\�����k"�r8(j��� -uj�L�'(�-���̠��,r��8aSb�Ӕ$tx@�p���:�����f;�ɓ	.H��ك��-%�o��ʬ���Hg��Ք@8ƺx[���i�dv�H)���۬�rq�87��F9���촾@S��h��-V��4oy)�䥝�k	9�v�k�`�a$�y]�1\ �S��&��+�F������Ϙ�E2{�py�5Λ����[h�sE*�|soK��a�RXcRp����.�G_:|��&C��0�����l�i{ǅ��R�_�Sݹ'?PM��S�p~7��ƕ��k��b���H��>��Q�v�+F
�9Vp�U��>{�5(&紨��w�PY�aģ�ȷ*2��A�X�A�2�u��L� Bzi���ѻ��TD/W3��F�A6�U?�Os�q��3E
�ݧ�`�Й�./_&b�<v�D���Y9H�����Q-J���F�k�lfV����]UT�_�vnĠ랢�y4����%����ei+���Fi}ku!�L/b�lr�-�Pe_+6��}~�IqV������� y���L	髍�ծ[%%T8��s��S�L����8z��ōr�=�z�Y1���\m�
~!T����
�)aH���0��Vy�Q��z�VG��$���+ m�\ؠl/���!�J��
t o�"��N���F��h`t�w.����T�ly�H�z�����Џ�K8p�ԫyh�t��O�"����5wӪ����2�D�'V�]��L��D5}CɌ�%�B���Y��J�_}w�a]��y�@"=���9�������@q����������KC�{�����ZY���P�{0eޣ[p	h�VHx�����@����}US
�������E���	r�B9�[,ةX�%_U�ZvMG�j�Ŭʽ_zH@��b:�ڰ�����Ct	�l����1&�gjì�J�: �(�,�~�SjN"�^�}��)����@!�d��X՝\�-*®L6�C�4�Kް� ��Cnb�����_{0|���Ír�=Q�gײNx倒ݧ�L�e����
�
.ȕ�`�bM�UFi1Lb<O����-׺ͫE�.O��������R�}P�s��Lۡ�Q-��(z*�����s,D�y��#��G����X��ݨ�(zp�	T��8���H	a~�'Gq����yM��`�#�%2��"���N:!��?��*ҦU��B�O����f�閻��RK@Uy�l�7 ��(\���L�#̗u��*���d�?,6:���ڍo��������Ě{EG�������DG�w�]�`ʣ���13
o�
B�I�/=N������-hl����z;.��[WZǀL`Y��tدw��ϳ{�$�+�h��~{D��G|�ʺ��x @�`j(u����e^�$g��L��(5^F�M�V��ջ�|s��~�8j� uF��q�V����6�ܸ�6���Ќ�Ә� c��a�Jv����~���`�
���QDP�dHA4���U�ך
F����_�i1�����2x�;H�.^$'Y��"�Vy�+�AX/�/�%]��a%����cH���Mt�Cn�R�i�G]8r����6��W/�2���M��A�
ɤ6p�ռ�%����B�����\����̃'!���w��u;S��U�:�p}N��R���q-��3!3���@vtZ��#-x?��t�
J/�i���YЄ�5LG�'�ʚpoُ;��)��E��%�"؍5��i�"�e�����!LE�l ӯ��|�_<��u��|�����b,����=�/PV��F�;�l'US��i������3�ڽU�<P��eJ9�w\TS�ko�׸����-��3�@���1�:ڵ�P��v߬��}F$�į�cٕ���8�_� 
�r J�,#\*6�1K�6.��_TK���tw��u�8��P�&��U!�A��i�T�eI�Ue7�<��� �Y�c@��6M7��C냌 )���!���d��n�>�J�=� ����}~�bO�it@$	N��v6zm�8aЛ{å�x�Y�����ful3�J�TË��r'+8s��9ԟWxt^kF���0��gS�����6�>�VW&��#�.�F.W���<*|k�Z���fg�-����OP�������/����U�2�L>/�4咔��A^h !�@�TH�[�)8��	�_Q��{�I�d�Vf)�ٍ��5+[l���,��v5��������+����3}����I��k�Qy��ZӽWH���wÎ��fnJm�����f���a�
'�d��>�}����ܹ�8Xs%V�U:M%����+./�iv{:3Q5;�a�^2��0�}��6pN����̀M!�w)�{F�!B[t��R����Ic��J�ʻm5m(p~��m%����)R���Ow7I��L�p�^�Vg"�Vwk0�U6Z/����|B��4���1+�� �Ь�F�b��T!'��5▣ ��THwé+iTAR
���N��(44tQmr�yj"..���l9¹<1nv��\�� и��6*�s:eQ�x�7] �zœ�i��qHoE�	-�e='֐q���B�8�ג5l�@��`�V��װ�x�Q�O�WԱ�s@){d~�l�����͈�@���eFA�"O*���K�m�re&v��ai�,=�o�?%}N��|�J�-"x���N�F���d�<@G�a캾"H=����3�e��/ߖ`���3����j0w�I���W����Q�;D������qT���3L���E�-��1F��X�P��o����0���^*��(���&��a�����z!3��m����������T�Q���N�2���(q��Z�E:h\<|���Ce��r��Z��0͵�\y�p�<u�P�2zp��r�yU�ŋ$��=�`��$��Qj@����?���,5��]�/�Fh6�R<��,Dw_�]�e���BF4��r�� ��֌� ;��X�~���ЇK��Ƌ0X�?�]:S�5�w�K�j�����i! 鸧)}I0�� ��W�iŠO7��N0$�s�����9S3�*� ��4�͏s�δ�1I`g":@ d����6VE�� ���RV��4�@/��[G� E��J�Ն��0�`Qq.�}�G43�2ҮL�c��zR�e�lUtl=����־RAU� �Ӟ���%��g�)}�d�p�戴Zx���{jin�}?3����L�e�趀dF�X�ר�D$wu��G����܄����&��۹|���S�BdR���EW���U�[.��-x�����ݍKp+o����y��㴸x��;\;'�H��>I�Ϻ���H�#
i[��#�S�q(_�F��ӳ�9پ޽FCZ�qPt�v��e�!��8����jf���\���!:���^���n?"����.���֜	8!�����t� ���4�D ���S���eHޙ*Ðz���|Pr3��k�P94�K�h�WY�9��l�cR�	��H8}�ؽE�d��3N��a�c�U�t���|���-;'��n,�ӿ��3���FN��\�4�b�Vʫ��wRQA��c��Í���ο6��KӁ*O�F7ө.�w83yǯ�S�2��'8�Zl�/0,6Mf�X�:���J�S�r-ˌ�K�K`��-�e�4%|A�f�a`�;�Yo��@���e���0K�)�1W�TuB�#ݐ6(�������?a|"+)p�����CK�°��ެ��u���=������-�{�3��Ј]�����[`2��8A&�TG��۔���(h�Z_���%�z�_��=��z�b�_�T땛�+���������1�������+�	s�U�������	^��g�d������e�/���c���C���ir�������͑3H*���<���0�%����6������5�c�=�IE9vB�<�k�g[����WJ�C��pZ�>�u��t��Cۮ87�c���wo�ک*!rdϠ��a����K��P*�o��^�c� �=��Je(?'1/��J0�$%�=�+w>�b�����g��f�mn[���7�T0��P"թ�WgBˑae�_�����J��@�ޟ�B(&V�F�G�*�Q-Y4��W�h|T4�_���_���{�Qvc�u$>���r����&9�=�k�����Гn��Y)@��&�)'2WsI���ᑲ8�,'�k��
����;K��#���Dq��j˳>u&�u��NB��sx7|x(=��l���c/A&�\�uj �u٣4~��|��	��u��������3��Ԃ�G�C��H�4Y(`����jh�$���t�#V"�&�U�/�?^1?!���>�t�6+��E��h�K������x����mf{-'i��r��Ys*�|o�O���� IB�n3��⨌D�ɽLE(�����T�砡����0qAdu�K���RfuJ���ER�|����S����O�U���5����>Y�#6ʦTx>d�׶mx��< ���M�=�&��I�����Flc�:	�̳�j���K���ѳ��-��'��e�V^վzN�5����cp�7yʤu\�>�I�?AK�i_��Z�>d�W�#b�x�OPH�I��S��7�+4��*e�*��*��EJ���O5s��=����8W��B�l��%�>����.j#�4dХ?�N8�k錷�������o�A	�r%{�9X��K��Փ���E3Db����,�c�`K�V�%��h��V ����}�r��8c_=l�3���	�^��a��Q9"��6)]!6Z�[�h*�����J�"��	C�+��[�"'�JI�����Dƒ��\�y���gq����wP8����;���z�|[ �w�'��U-���w�B���F���t>f�2�G�N��J��ͺ'sѨ��2EF�	��S8̨=�k�3�JϞ��u�­��ut�����:vWg)$T���%E�-���zw��|v���+��t�Uj�xC>�F"*%}��*���t�J_s��:�HM�e�$�D�"YNoRv�!����X���ˬ��,�����M�ą�t�}����D��j���h
�=�*`Cs���h7�[1w4k�׌����<�j�����աBj�����W@�b\q�yS�
�l��C������/(ˍ��3���k�Ӷ\4_GA�|���Y<�H:82}���V�nI�Z��W�dD�����Pc�'��Wh{��fC{�H�q���p	_����?����7�?�^���tg
�98ytQ�z:J��n��|��*�9���q �߼44���q�����`5_� �v=�ә�`��A�u��2%1<媧
t��<=�?'��)
�ѫ�����l�C��`�_�����b�Ro�WT�k�$Vݬ��Só㽗TD=�����~�f>��2��1G�}HI2'|�6�y�,�Zʺ�����r5�q���4���u��(�w(�l��Hԕ+���6o�?K�E�S�W���:'֠\���uJ7���0�񛲹���S�L^���L�v�p���Vb����2�=+��A�K���bz� �'_x��;�t�}!�0m��z!;r�5�1�iH3)�Ѥ6�[[�µ�4��J�1zS;o�9SzV ·�#,���	�s��8A�����b�|\��Vϟ�mkGUM�L�;.=/g��z$1ڷ�2L"cL�ܗ��ۓ"{o�R8]���B����9�Vcw�f�<��M��X�_0"NQ��=����"��
�MG�P�J��R���V ��GSW���`�u[��y~va�k��]#Kʲ�>.b��h��6��*�=Y},F����d��p��TG�b�G���=³��/�q����GRF�3`8�<q'3n�Ox3��J!�:���� ����"��7W~��Sih�+�{����h;U�@oF�+T�B��{�[4^�P��rUR^>�����cO�L��^����t�{i��y|&0��p=�|�I�{<=D��b*��P"�l��g�=���;K���Pl�Q��]�:-��5�̷�
@:�� ���w'�,n�
#6�틋hN� �\��~s6^����
�wȓB�1m�Y�`+����"�-���vl��p���X]EK���j�gv��Pߒ�VHW'��a�19�0��,1�����P������l"P5ys� %<8�ױ���!P\�VF�0�֙s+�(x�)	������1�'`��vT���Ԣ��������+�"�w�(,�K�5��4U~�m�r�J�8 	���p}�g{�����1q�ŕb���#�3t\�xӝ����=��+���VD��\��?<͵j.�JQ���Hio{&�7�tMs��춁Y��Q�/���|._�Q�yj;hZF,�^hH	EZ>�z���Y�R�ۡY���c���/ӿ���$��=
,�wk��,�pc@��kŢ(Ķ=�[&�Ka³_�ō���8`%O�f�h߇b���m��41��n���;v������F"ٱ�1���rkm��SgKՈؿ%��%pWM�ex�QYf�H���k������+ȟzʺ�4�T܈�PKs��E��O�'��f�E6,m�K�����uxm����V������ �Z�ْ�[��B��F\��0��E��e��:�#ip۠���?ʒԮR��@���sK����{tYs��[:"p^8���� }*�ɛ#3$ش$,	Ʀ���$E��~\o�5Ӎ@W�{�]���s��?h?�N��x�p��-?���2-Lp	[�s���N̓y����?����w�.O�Y9���h��tD�=�L��K���9��M<��B��Y�yK��.�>iv�ޤ5f��C�U&P���'�ئ2�ts>B����q]����v���''`�`I�!h�3X5� �w%��C����9��\��^&�y�X��]@���Ec�J���`�L-�
_6wws2-�����l����Ҷ����G�u�a#o��ϴS�.�4��$�wv���t�!#*�� 	�r@��e����R0�a0+]���Ԡ�;�v��z��^8����L&�wO��J5_��v�� �{�EH>F��;���Αd���|Z7-6�h?��$����k��[պ��Y��|NP��xg�9����@#�>�l* ��FZ|g�eAR��8����9�dI&J��µ,��a sp�s�}UB].iͶ�<?��,���Γ�W���	&�^�8������a��G�[��Zw��ăB,'�J���1d�cJc�@��ą!1�񦨮j�]Y�\�)����l�m*D2�_Sa��Hl
4�/"h<������H^&]ҏ��,x���0$�nM=�zB��u��~wnż_I�|�/J{H`[S�=6F���S��/��l�u��^4!b��M\-��roVY[Y���O�'%�Z����'�|g��-����B�_-��Q��xv���ꆣ���Ƚ��},�B; �K+^�^6��&F
+�����T8�|��E-1�1;6F�.M��
.�`��=%$d"`8x
&��v��.��&���g�f��"%�3�Wz���\PW���8�����㪶@�g�o5+&l�G��)��/�&�UD�q��x�{p��!H�����C{��o�dn�?#�c��H:�A&[w���]ч�r}t����	�����Ao@��2Sw���� +<j4���P�%�Ά�W��z�>�ф�6y��\�R�^�_9��,�j�ߝ���b��ø�S~��l�����] �6�x:�'M6�ӟ���=�?:�g�ƕ<$�+@ê�Z�v��gQ�"�ܨ������[g�b {�� �>�%��)Ҹ��� ���7H��q��c��2_��7P>��`������Gb�b��i������Chʽ��-I��=t�'���D}�3jP��D��-S���XFD��/��O�#\�uR�?���:��t�W*���>��ϴ5'<Hr�WӉH�B�IC�@wf}l�s.w
4���3�J�QJ�)Y���W���X�:�ھ$7fps�nL� mG��dA�gs�d�;��8�р=ge�4[M-={��ﲲK��

���2
p1'�js�9SWZ�{ڿ��+�=����B�f-�'�@�N��B�3j�P-���S�m�ܔ�@<�� @��
����p4g����B�w�\"4����e�2F���R�}�����C*.��e���8N�)-��I�r\�`TrPؘ5)n�o����0p��>7E�Ś���/�B���(߾{I�X���V?��Yz7l���:mEf�K�ę�Z���l�oil�xO�R�.�� �$]�X���v`{��r<?���"�:�P��(�~/ؿ����c��N���q�wB�7A�,�!
O���8K���O���S��w�k��?W��i��� �;�����"��0r���)(���W�*b*�He���
J��L��^��6�T���0��i�	 ]��{o�`����uZ
�Y`]s|5�)��Q��j�ޝ�1ڛU&�3�v|��� ���p�8����l�>��!�#̘���Nxm�AV��=�La��i�E!��kE<\�@��_�r�*�m`f�1pc��k����3�7�.$ϭ���2AG�i���y&��<�R�H����f���7Ώ�֍����6�Z{ڒ� CVS�"�	p�.��y�����s��d�M-�!'�g�}��^�g�4��)�B�d4]�W0�3����q#1i,���%Hg����΋��&3l���=@���4y����;����¸ҝ&E�(�=k,5���NS|���� ����x�j��!Ԋ|"*{�
��\���k5"|!�	�Ψ��j��+�1k�J��e__�o0^�E�c��W���<���pi��~w�/,��?��0����i�J����1���=�\��f߳$��E8+��_�C�@T�z㔬�cG�Ƭ�@�7�u2[��{;�gv~�n�������Cst����o&�Ƭ�5��]��j҄e�=���2WRTs�J^�ed�1X�֟���*�P�$W-�G�%�w`(��³�qt9d�{��]���t���Z6���s����{Ѧ�"2&%�r�.����c�^�f��EuOޖ���}��>I��U�ɰo��u�1�����i��<j�I�P����2��sS�L��]��K)yJ�i�u�פ:[K}����~Iլ&'�lf?�9�D_zC�|;Ne�? ���j�L1/�BW8ȶ`iQ�J=	��]3ww��q�Q\x� aIhVa�2��&z����Af�����smlk>PmӸ�g�jr�t���"W���w�nF�%�1%��ջ�B�w����yu�,�"��W��}���18F�V�B��o��)jC&��k.ʥ�G�⍩7k�/�4U�Vك��l�v�٣�Ꚁ�q=o������A[���Q|\&�;t��g�ʗ�j�
�fH�D�tן�dт9
=,.��R��%+tY��m8�����}��S��rm��}�������� 6�#����s,�J�,�ǹ�O7�ZRk���)�It	hB`��i��C�_��~�s9FJ���`Ϻ�ҕ�Ʃ��Q| �.�Ћ����0�	��E$���[�K�:�7���T�X"P��|~��2��T� �l^t�},�b��.C0
�ʶ\����9�m�JD}�&l��Q�Q��w%�#L�^�P�_���j�s�g*e��]eʪV��#=&)��{�KN��퇏�"��̳�F*rִ6��>�etmvI᭑L���Grr�9Y�i=a��}�tړ��!Œ��6����2�8�yGl8��;�a��ob= lY�9�"	O���]�_OvV�.�=/�������P3��8��+^�N��IS��o���>�)ݽ�t<�k;6�Ն؀)%h���X�]&��0� �Mc�c��L6���o�9vNm�Y������,f���v��US֣ �-�N�)��Q Di�����Y��Kn�	�3r/�Bp�����.>0�:�A_��/;�$(�����Ђ	"�nu�� ��c���%�Х��9N�/k�?���N��JºA���?"u�ͅ.C�����xv.�cP*-�}^����>�ŵ�ϲ�5^��Dd��$�`�\����?��������)�9��@}���N�b���ԭ�J� ]�(aI�.�=ܵ���mdK>'o2ئ,�#�))��m>R���$�,�A�&_��u��Qb#��.Y����A�py�h�����	���	5K�sKZh�9��c�­3�����o�f�Y��мq�`��M�YmrtSx¤$���=_�2!3���s����Py��)a�	i�Y4d��4%���$K�6ߧ���]J����9�7�������ܙ�{�z����	�����g7�]#wW6�]u�U�w�.C����mH~�z	(��&�����ҎYy1s#���y���L	��N୼�Z��_0oX�WT����򸜇��qI<'�V (�4�ƺ=�{Ԛ/�\1�W��m�M/�?�V�d�uh�����R��'k\S�[�ct:�e�n��.�˵\�S:����,��zM��tf�;,Jw8��"�X�"�ѼX�*�:5q����fi#���Nk6���Iu
]WRiH}t�����]����n2�4����m���֕t�8���Z�[�ō����?�cݲ>�G75��y���($�DS�ؕD�=/�\G"\�����>q.?ꠗ=���7����.�^%S�h
�R�.z�ґz)}�\3��B�5NX��1��[DY(h�������L��\Q"d�p�Ǫ�֮�W�Z5��6K��z%�,�8YN���"��ç$=wd�o��`6	�}mh~�u��V]�c^0��o��+��.�!w$H,۹��v��(�R��$<�S��k~xH���z\%����PA2c����_|���k�flQ��1���T��r������Ƕ���.�&%n
��Ҙ�������)�2]u��Z�^��X�ZYyR��������YM�M�Y�SQ�����f-Y�f��2 4���͈������H�}�v�ps���S��_�TR�����o3����(��[{DS���~�b}���vٻ�Խx��w�֧�ޤ��v���U]Y�TFSx���a��
�I+f��숆�N���M�&Q��1CJG]yY�G��α�E	]QI^L�!��M��k?6�N�?��	���!�3�L@�-�,�4	�Y7�7���;]~�֞}jY�g�\�������E<7{{�F���4��/w�E[ocY\�ȆH�L����ZK�Mr�$�����EÍt����S���b��1!�6d&q;Z�����L�|+�����~�ى
����~b8��ji]�cX�q�y�`��pP�ޘ��F?�3�Ĉ���I���|E-vFڥا,~��4YRuc�d�ٛ"3<C�oF���ec�^v�WKdܴ��k�wV�:�Ҏ9�����DO�*S������O?�uޝAog^��+[S))�8M�Ϥ@�pr;��W�;i��@o��tJ�m����/�e�N0�q'�����p�ދv�D�p/��������9 Zh�X��b��O�@���-m�2	5���V�g8X��R��n=E�~c��N�8Qݐ|��M$�׏���vE���O?;&X���q1N�������4K��h�`$�F�b��*��0H��O*��_��w�WVdsiJ��� �?��F�exj���+>j�(z�C�;�x�Ӏ�)}T%�/=��A���6f�my�<��(�ۺ@�Fr��h�KYQPMMȜ@)
���G0��=4H���= ��t/5H/P�8���_��V�(jf9�_��C �e-�PV��UZ�a"����`1\��H��ء݄񾞤i�&4�[�MF	��=�F����b�F�>���3����1F3�ߑ���yc��@��B�W4��{��O��|p�av���v	mkSP�ϡ�$c�����k4���Q5x�խ6����о�\��w�"u�^���6�C�oYб�`Rb���~,�:�7��Ae��坦�����ӦVkKOZ%��[�<�1��.	�l����=6���z#[��NՂ�WJ`�+-C��=�K�b���N��*�Hj[?�
qn�@p�y��v2?�B)�D̜w���d2�Uh���P'@�e�Yam�'��>�P{[W4d�t��Up�\2�/���z
�'��@j�����(�;j�=�(�a�R	�<!Y7 b_�"౳�?8��*���h��Cɬa���+.Z�6 ���YDU0�a��F��?}1d�(gA1���80�zhL�q�?�������!OY�ڻ}v�D)E�)_������4#?UG�wϲ6ǽ�!7~����/��ϒ/*�lE�E�� �*����'!q�{r�����&�t�|a0Tz~�<~�oO/�楸��z���|X���(�f�Ec�z�n/�i��s����0�f�, ��:9r�{�&Wfe���>����i7qB[��?Z>F�2Q�VH�;��R/�ڇ��`RO�/�J4��t��b�1��u��6^�u<�fp��
�谶H���Q�ֺ�XTb䚙��~�L�r�D��z���n��2��&����G��6lq�):��Td��ń��,�W	(��_�"� z� ��e��k�l�^>?����:��-�MVH�:��0��βl���p��q]�I̠$H��0z{,3���Aa �1���|H�z�5=ɼH�$���p��VV�)�q%>aV]5,�"������&�0�Hp>U}��s/h����b�����%�X���qF�C*$�b����9/u��$��_�OH�޹��xƔ�*�w]pF$����:45?
�.SJ�5nM�d�<�k�C�\�Od��Ģ">�=B��#rHˮ�o�,��ypԗ��㣃�U�g�����l�����[����)_0eu��W�;.H�D�JYrp�o�t��),�Ⱦ��TԨ���μ-��Rše�.9Aï�πh��IO�Q@�i�W�42Z�Y�hXA2��TG �
 �ATمk��Sj'��"�J���P�ȏ˚��U�����a4�ƞw�M #ͷ7Z"��H$��z�(���4�`Y������e|H��h��ip1��ZS�y�.� ��gx?��}{��|�%1�ՠ�� &+���k:^�о�u�F�2�}$��4Q%��4E�����/7_�k�����,1j?W��M�M����u�#Qv��U��ޛ�p���}W��i=+\�Ą����iZ�˔�2��S`�}af�ו�)���hJ;Kw@˓ބ>I8��PTE��	�Ҳ]*p�e�-��I�hO*���*~8�j�h�Ǳ PN�|���]��.�u6D�lF�]���u��D>�����>��t���c�tk
�){Tå�`��G	�[(� R��ʽ3(݈>��8����oًE�>���C��	�ב �`�i�Y'�cy���3�z	5�>-��^.<a�$�4��)��/)<��9������46`ـw۰ψ���`y�$(˩�S	X��k��~�
X��%��l���s���ί�hX�|y���T���b�m��ёC�E� `�9@�TK~��e�!S��I�}O�ٸ_Ӛ��rˑ�ɟ3���\AP��z��m�����h@����i^�:u�6h���[Gr�V�E��: ���� ���.��� �hZ"<��ȏP[u�y�[p9�x�@�YX͑��h%R�.������A��r~�>���njܓR8�0N�6P`�ԃ�I+����	%9�Uѫѵ�IA'�\�[t�!��O\���fK���z���F,��!am<"�F� R&����s!j��n����?��lF�7�oy�V_y�Ng_��~�{��*��{�,��x��b�K�{���Ap�z��ղ+j0J���㛭��J'���z��_��>�M�(�b�(�ĩ�m ��U~��FWI@��-*T
9�;�4Ī�
}u��HH�-�~ޙ��<Y	�=��P�� Nc���<�zl΢s�<��6
�5,��a5�:!�}dR��!�X��J����.�H�gXԏ�8�i:�U�F	���1n����� q`I%��bZS��_j�F�m}L��!>
_[*<�p�h*%{5w���B�d(���y~?�%M�U`�G���Q��z�{n4�Q�����ů�m��ܤ�i{sV������]އ�r�;p&ˠ�%�~$�V����H�7@dl��Kd }���-_��ձZ�D�9Ft���T=����B�務���w�f "�#��?�����:��7�u�+���Fn��N��{q��F��FK=�eU�{�ÚI�#����"Pc��<�C��,�z������҃������m5��R羌H5!� ����])�ڬK>��$Ɉ���C��Ȫ]�/�k;���$��2<NyNY�V�&��mD�Plaa�_}f&��qWuG������Z�-ebT��������#���5C2�R9�~�ָ;��8�@�Í���_���ɍ�q��D�߳.A���\�[��Z�6=;�F'��l{ߍ<�7j�<5��>�3r<��+_#���VCg��8��8�v2vͧa�&�ye�^-�؂ �����&��IB�~��+�z�ǎ��̓��x��M���Q�>����Oq��{�3��J�h�X�#;[�Q�ώw9���n��a̿�2��x5�?��j�x�N���T���\=+����ɠ��e��Y�� ��.j���ib���ADP����ͬ��#�벵f>,����7 3?-l��]XZq���<v�w������'��������Q�Z '&�&�xO��鏈��?��4�a���˜]y���*������۶Z���'�s�_tw��W�SXz��B����W��`��Id�$��� !1��љ�.$>���56��zWX��,��Of[?LO��K��BM����zs$%�:��<��\C%!$u��0����2�hAo�r��%��_[.�#󸕢�\��"���e��ap
ٶn�*��!v��ؚGznx�:�������o[1,w �^W��{��4R�ք�#|jiх�O�\�9~�vmZ'+E���`��{��VV��fǛ�?�?�@ w�#�3���	���8{VK���ʣ��G����s�iD��bW܆#���&[��<���ъ��{8��q��T~�J"z���M��ȭx���^��Ӻζ�`�N�_�6L	���#�,M�/��C�z�������:�f��Rj7�������f�<�s�h�\��x�&;|8�e]�:�*�=E�Y)n>��F8������ �mM8�
�%�J�����4�9���'	j�32��\���

��VR�,	(}q����R�C�q�BM5�������~�;��A֘bֆ�|V�Xt��1�����(�*�Ѧ�xft��~?�|p�ky����F/{�h��.��L��?����6����uY�B��~��A&br.F?�_�ݓ���hD���M���)A�A���aY~��VX�K�J���g�y��Hi���𓶘����ЛU��Z�'l? �c�e���zV��S�bU�����bnط�6���鵾:�kr�<��U�w����C�]i޻�Q��bq~/�:E��ڒ��A��ݕ�s��U3{��%�)��h4�RN�.��
�hݧ/<02�e,��wGJ٦�V�Q��C��ڬ��wS�.���$A�7V5���	��3B��c���/"h��� �;��oe%�+\5��R��8@[	a�xPA)�z��nS4�A���& ��������� ��G�m�m��=����s�'-NB��i��H�q�%�NWVaCQs���"��L�����p�������O~=n��}3B��G��
�C����� �j7|�A��G��ED���ĸ�������{qw���\���w�ɧ�'��b�� ����`X���Z;	I�A�vM%��@D�RB�3�8	_҅�����l��F�y*�~�Q���+��@����5F��?��sd+���ĭo��#�Rf�v��R� ���y�s8bl]�=�X;$+�a*������#=�ҷoo�n�������%Y㷮��(<��g������Õb�בh��A��c����F��.��R��6E��ا����ݞʾE��|��q/ɺ uІ�#�֔e�7���X��ys�mE,�?$&tYbA*���_BKM�<��|z�ָ�pĬ�I���dձ�@�7S��D��Ѧ�D�R~rY���g���?�������9�-G����`?��1��t�c��!�	�J���3a��j@#���J�Y&�����T2���k��cj��;@f��H�U}�Pm��h�����,+�:�:��V/���2��'1sy�USh.9.h����z8YNf^��l)�m�5�;+��B����ֱ|	Z�#���㩗�So���R9?{ã�?!5?m
ɏ�O�҆skD���i�	��EH*���ˢ�7MU�����3�� �W��x��K'�f�%�5��$��G�kg����Y��ю':�!�w�f�F3�Q��x&(>\��/��D���U{�8S,��S����~��w������>�52 �Xv�16Q���Iu"x�@��9��i1u��m#�^C���\�퍕{CF��_WX!}�b���=d����E�7������Ԥ�f�ݓT�ǗF�Qs��h�,�B���;ڹ�1��[��R��tc�����F�Ņ��4��*[���T� ��R���[�4I��*�f���^@�ZDN�D��*K�GB��ZK:j*�15	ʵ��]�}U�zN]��xz��C�>����LB�2�8��0v/Uż�L&� ƾ_�,�^��EK؈�|E����Vt�9�fiF�� ���R����[�^��K����\�-���Ԋx��'
� ;�;��9R'K��SɆa��+�߮�;�x��̶��K+q��/J�m�����}5������"ѭ$��XâY��;H]U|@��j��B���l�oz���J%�b�{5)h.ؽ2#���@Z:6�3 bI�^:1'����+<�)�� �_=���M��ҵ�s��U�|�S�y���γ4�L���8��W@��&���k�:�,@���'�Ka]�V�k��s�M�Y��\�����T�e�:�ү�$�sߠ�d�d҂x�`��$3T:�W��RD��ۏ8qK�<do�۱����DN��Guk��
�h,�
���Ym���X���x$$�!3�K4Ty�C����^Jv=�m$��%��=^���	���Avsn4P�W�w���q�q�� +���*��Ư�� =���
�R��pvS�Z5mC�ki�e�/o�8�׫ǽT�� ߑ���+�%c�(%|���j���"��c���u�w1�#�J�J�j�,������32��Ľ�֬����U+ͯ���w�_���O"�B���s�2v�3+���(F��Z{s�Rhz���
�	;����NThU�B�x,�.�uskw�	h�b��te��<b|S���n<]E��'\���W�7� �1���:�}ŁP�$Ѽ�h  � ��U�Oy�"̂$�t)dU]�U����_�c�	x<�����;*(��J�5��2�&�/+)6�u/����/�}�#!`P8�}�	M*9�7�	��(�ܽ��@�k0���i!��mh�E4֪w;��X�_;Xf��m'�"���&ֈ��=;	�u�q$?^@yXD��{H�^q#Q�v`���
eH=���g�E�ӄu����N��e�$��1��.�5��Q7�}ƶ�R��V�F	Ę�
^��O��;J�<0:���x8vA�u���.vP/1�7bA�r�3j����Vg����y�$�/���D�Ȣ����_w�jl���zn����E�L��Cg��؂�Ϋ�M�ֹŌI,V�F��K��_R�Ub%+`�C�N��}��
�_����[Z��Uݵ_W��Ń/����x�9�[/�`G�YI?�zO^��^��Q�Nƒh�Pb�_�Zʂ�Q�\1lyL���4m�NuPj{Xג�^��ٟS^Jq��t1~P"ȉ��/7`6�Y��l�)՟�/K�k�wV���!�Q�u~&���c˄޹;Zg�ܚC?pa�I�v*��{�����,��g��.d�Ċb��я
g���=��Z� �U�Ӯ;jF���Z��Uvϔ��]9C��:^��+65�3�g&�����̻�w��[[�^�1��̨���/4��j��^��% 㓨���O40g��8�X5E�� >�i�/&�o3%���9��j�Y���F�8(Z>)�Z��VR��Z��X�7%�j<�p^�h/�#�dOg�Z�N5M$4[��{�b����B�t;���i�==,j*n&�ׄ�)�MB[O�0E}����JƐ�	����:ح�,շ�g�w����&M�9B�f?��v�p9oG���dkE�^O�g�1���%4��35T�<;��yߣ�a��T�.�%���زh�Ԧ��pDh�y������!�k�L�Џصg��<�;�h��|��2+pW��
���z(:�(܆�z��?M�K$�k$?�x�(741�C97�����>t��u.�zD[?*���A�"n�qfi\eD�[���� �Í��?i���Db;����gP[hb<(9�C��k���l%������j'RP�7�/[�@q�����������֮�غZ�G6��a8�__"g�k����2=�@���*]��Osy����J�Q�k~z/⭦M����p�n�/����3j��)�-q��q\�p�K��m:���G���#9��55�HRn��Q��V��|��
^{�� ��a��3D6t�އ��H|�G��e�:�S��]���o���\��H��TE��݂"uD�N�Gaĩ5���K��f�N���'���d�ӟ� �{��{��ڏ�Ǔ�>�j��7#*�,�ַ�累SM��T����F�G�i����E��J�~e�^uN{7�.��,�n��{Cfl�J�#�/ @�;k�  ����%����\t��w'����[��9��л\u�K�ڵ�aX�SF�*j!)�Rj��(ŋJ�!�ױ6��`E��,�2�,o�1t���U��Y>,ԝN���W
槢�G��;h�v.#LUKA��ޕ���iy)f�}�a��|�.*D���L�����Ԩ�y���9>�����̹k>��S �Z�<��g(�p�e���i t�2n��K�f��=�Mc�љ��h_�+ς��2U�XR��T�&�p>_y��*u�+�`X��'sg�(X:F�l�5>�R��Bۏڗ���ۛ(�|_a��/v%@�����~�G]���<S�4"Q��ĳ���j�Yu�}�7��=�@���N= :o�mmYqH yTe�wޔ�����B�BC�,�|	��۪�z����;s�PD�׿nhφ�l4?G��K��r�N��f:�`M��I+���#�\A� �^~�*�Ĩ�����g��h���L�1���x��V����� x�\e*-����Դ��67�;��J��0��s-��$d��Ӛo$�[�P7ƙj�+��T��Z&��nɀ��tr���2A]�������؛D��:@�YDI��ѓΐgX}�el�%�n��
���H�(��w*o�C�(�!B����'��@Vy�]4�%�D�w�i��EH�K�,!���/�j�/UWg�_2`�F�/�'sw78ӢRy�h0����k#��?�p�����A�MR�����KD���N�0�v��*c��{����a�^��tP�)�G���Q��|��RyE�sb�Ŷa6�]�T���8��U��?�"ܷ]�B����E�ܖ�0U4)��U���չJ*V[Ҁ�ޮ_:�P�r�wy�&L�7�q������h���G�2��w>5�'�Xed�D&�Lgl��u|-3H�o���ۂ����Bٿ.��6�Ɔ�����'��A�&��|��o9sXӸ��j��R��|�4��bZE�d�a������0(L�r��Վ-������F��K�O�i/~��E#�J2�3��T�����1-�x�T�bs���O�j�����l�픮�9�X��?]Ŏ��d�i�Z�i��Qʵ�KP��N����#(za�ܫ��q�sW�eԥ��I�V�U�wZo�{e@pG�(�Eɹ��wM�S�_�o�bf��~���4B&�!,�r���mX6��*Z-)��lF�Q�DJm������/-B�����Q���Mĳb��7!6G	��:���=��_㺅I��bu2��ߑ�����ܔ�7J�*c*|�u�ں(?���1	�ڦ�{�ˆd�%�J�s9�\�#��J���l�բߨ#"�9�U�CD���uFa�U�An8�۵`0
��(F���E}VVj4Q�l�����y�;�E��	׵G�3r��d��*��<X�I��}���[�7��_+�����rMsY��\�R���_t�bT_���VE��S���}Ԣ�ț��	*�K#�_�Tb��{�T.�hG�;��h1�|�ab�)��G)���"؋�jl�/	NǠ_��|nd��(l�R�a�L:H�@V;�V��E�?$��zղ���D�j5Tٳ��Q7��&���pl�peՕ���V����w9O����z���P��F"���6���
ւ
��A���6\��)�,A4�W�^!��6� Ȫ#��;4|��'�D+I�3����!��؈M�>�Tt6���L:w�%�{�:�y�B�dv���Q_�gϝ�]�j��� �"�6?��� ���h����9y�i�7��[����f(���h��y���η�	�Mx��(����:����W���MxC{E�*��Ya7���+e1��V��զC!#�2w�Y�_�k�ҁ_����a��>�>��bs��o�j͟^�Ũv0 Z��K�w7�Z� ��Ά��;�L�����Z�;E��	vjC̖��=_���Ug8?������
;�����W�ŕ,j!��;,Wi�)����g��n�¹����mZD뵱/� �������l+KSK��"�<vD�=�O���77�d;���%�cN}rI��O4Y{��$Wn�Hd���4)8�(��x!W�%ϏtG!K[�K'L��w��7)̸��n2�iRJ��R���I!Ω�������ҕ��V����¦҄��M3���D�G�Q-�-��d���?V�2�l
vM�Do�9�>��M0IC���>!�SV���֨I�}����QUܪ��n����E=�5jy�z�U(4����*���	��p_r��7@tb��Q5iF�󒭱��%�1K�/vugŉ�5^�zƱ�wl�"wH<���GT���j���a\�JN�����,��g)�r�D�����ݑ �h�����?U�����[���E�� QF�DT�W��P#f8�`����k�P�\�WL�p	�@�o�HH�{�>��: t���T	.��빼��ؗq'�Z˦y�)��*ꙵQ홯�vK༝T�F�*>H�	��Y��Q?���+<�@�HŲ`=�۝��9nzvQ�~�a��y��n.�W���ÊQE��d�@�ט{��;�<6z�.�L������Rn��P�s�^�&�czv��3=8�C�)���n=��~�z�O���N57�0e��Y�T��d�RCN�/VW\��!n������:�j܈�v�|Qh���Q>�J��h���>דU\ۅ���l7��y�S�<��{�Ⱥ���4>X�/4��t� ���#V���O��ȭߖdui%���"��B��)���$A٣�xX�<��K���Ea*�#�����Jg��2�d܋p�<���S�+��;r$��߆y0���}�t�\[d�\$<��>5~}�X�9n���T��!�V�5Ȝè=<	"B��'��`3���5������n�7H�Th7�%���)|�%w��[i�Hv���f&�_;�j�'��[Ya�4��&6�e�b�=��IE�
�E����*_�wbM�0��M�٥���	�+���8F庀ţ����ٕ��^�/��MT�J�P|�*�N�B�M�������#�œ>��0�Blat������zz���ܸy3����-,5����&5���c�(����-����sv�x�Ϧ�]���=��SxA������A��bɠ<�L�r�4b?=@�<S�މK���)}(WsƱ�`e$)�$X�YZ}���}Mz9}��V��V%��A`�;\�|w�`��eDA<WO��'emkq��!��Rݽ�;�j��<b�j=�^���k<=F�^pj�8i���]5�v��Ug����WE�[�z��})Wc"/���z�����ׁ�I�37�� pP@
�Y+6��N#���!Ѐ���c����bV�X[��>$��7xT�\4e�̨/tl��3y�)��P�3z�>��cT%r�G:�
R��^��n� 䴪su%x"~��R�US��rv�z���*��y��W����ښkc�q���qlq��7�:��s:��h����z�%7$�e�G���m�ߊqiԸE�}+4qx:r�SM���e�F��83���X����j����y�U-v`���OQozo��1���	,p����� \�i�[���t.ܼ�v�h��D(�3bwhG�ɫi�ji�*�Lu^�u�դ�����V������qe7�^�9	n� 7�(��%��8)��
��̦� �F�qH��Zs�͇�M���a����U�ՐPˤ���~���~�RU�1[`W��I�+Ձ��B��m�J���B�������UN�7z<�d\0��3E����\���ה��Å�k����C4�_ �+�/?���'B�V_eϖm���!S�M�Β3�"'t��c��S�䣶+qi�	�,�*�O�p)��5�W��o�+��q�x��i�X�v�јax��Q=�y\_��@<z.&��ԷǙ���s��ŷ�a,~��A���79[�3O�ȬПT�����Ԣ�����+��~��*_YmMhG6$[��&��'�$�;�?^`�� |�=��WqJrӢj�@��,�?�S�Bo��T8zI�J�����ř���Wg�3}��Ҩ.K8����,�гEѻ����c���q��e{��s_��#���=��{Q�BN����X	[�Pm��yO�K�N�v��-�y��I$�#G�U�0��x���� �����HJL��(霉qq�R@O�B��� ��,�o�������Z��� �yVS�;�!7�x����߃u}Ô���!��גB��?+�~#�d���8Ӵ�VH���T���i�ĬYa\7�D<Q3���cAE:x�uOG[�@hb��y'2$�����&^�!�CoH�d2[G *��r}1􀝸Z���d�Box�g��A��&][��"S�M$�T���H�ԥ�8�0���r�k���83��P�ޅ�wH�-��X*ڛ�9��0�P���s�D�taOB���0������
�'5u�_���6�$�]�=޺N�5�M|�i�Z�p�,���� s���;�ȣ��BC��p!d�e}��9*��	�v���΋c�s��B��?Q�U&
Qf.�p{��`x���aoG� �[����f�K�s"��u�O
dO �Ⱙ��LY.5��7?��pqq������l{��+������[;�d�
� ."{��Q�!x�W��@�N�4�՛p^! !��C�`���v֟�Ĝ�=H��mz	����Q5��'j�	Ӊ��V��:�sE<O�r[~��=�t�/D��-�2vD��o$H�'���=���W8�p�Y�����//�*�j���Y߅�ZÕ�����������rcAB4�?���)*:�V+�b-��o���e�+�7_8�4*,�N �4���ѡ����/�y����dB�좒��T���H��=Z�mQf�wʕa@����jG�"�hc"�����W8f�����Z���(C���'X/�O�s���?8�'>P!Di��Kh�/��Dq� ��\�MR}M
]ܩ>b�E`s�q�Y1/hB�dE���Q�O��}��ktj��|��I�;x9� ���y�@ʮ2�M�����O�S��OƮ�W����a�RT�
�C
3>yCE�@)E8p���-db?r8a֯����`0*�\�1�Y��Cٖd�ǜ���s��-�в���׉�ڼ��֩�v����cO�v��1���ٷ��͔ ����f��8�p
Ӳy=��4���ϐ�S$z=����[��l
��m1s[�<2�BWz3��7S�t�,��<x׏ޖJ��S�x�蜿��N���I #�Y�܅�a�<}��
߼���Y��.�������.I�w	�P�n����H�ȼ�6����R{�͡x�w]�oO:�`T�%�s=���S�&�
�s�b�f��O��S�K����5I�ն~&�t���j,�*��"�sb~��uf�MNb�׿�U�����y3~���JЃ�����XD��������\�_��z�Lf�C1��bDNm2�'�t�Ҍ]B']���f�ྱ�żݩ�ȑ=�_��-I9t���gY���PM>��z%���\�u����K�u������u�rSadE��^-a�X�ȯ���Ԏl[Op�ZB��̧g��ʑ{�Y9:�PU�~@��g�A{J#�Y����(=�\�Rch�����g�]�߃��+<HowX�I>IR��M���q�=$uw�Ӫ"��E� ~�VFEv��6�"�*�ćmq����}��L_�����'Hn�=�5/��oY����v���4C���H�bQ(�ݍҿ�w��MȦ���y�����e<[�35@�|�����mU1J��)���0��(S��>)�cssM��u:G=Ea�M9`#���\U��
�V�P���g+�hX�U�S���QS�|+� �o	����L��X
���	�c�$ ^xC��*T<�\��}�[6�X����e@�	�����b�)�
��1��@E������\D*��E]Pqp{����o�0�Nj䮪]�#�r<�S�����,�oWK:FPY5�V-p9 "���tL�V���]�-�!gY�F�t�s��r*���S�Q�p�+��@�<N��?D�Ԋ1j�DR������%�4:��Ǟ������X�w���Ćb����G[)(�]�ٕv�
+~���:�̦�7��":�,���(�T�k��e� ޘ'�~��+j�zmDE�R��s����k(��`�<$��<�E��,�ͫ�?��)#�OV)kC0�US�?�Ö��SU��wH��=NnW�D�Pv�ʿ��թх���\��QCE|^�(?G�T5�Jq���[X�F]L��;���C2��Ӫn�\v:�#/�_u���X��w����@\�l��%�@�K�UMk.���<�B�)�1WAk�3����8��څ���*FĴm<}��A�l�x�6x��8Z3���#砾A�1 M/��2�1ZG}�У	�B���vC�e�V�{�+�E'��5�0_�X�r��\8 ��$���E��n�U�D��LO'�n���f\~eS���fn��Մg����G��a�l��d0��NE�m������ ����z�U�^a��tI���U��*��-��&C�}>6�Ɯ�����;s��?�������â�?��K���l�&S�������._�D�ٌ.2�΀�Y=Ƀ<�3�d����Li���Td��j�8J���^���8��p<� �4/}��v����KT2���({��wW��
�c�pƎ�"
�4�.�/�ӯ@����N>?Y�6� ��Pm�n
�=�K�>��b���>*[��򗱱˙�� ���w���u�4��MBIX��93L:��:2��կ�*i�e�1Ṱ+�*��HHZ�^hݤ�d������G��¿��-~�U�����z���x�Uw���z���x�O�2�#nį!(���C����0)�ON���r��'�pk�Ѫ7�9(h����arЈoe�)����^iRI��W���\l�@�;Kn*�A����#�����@yDԦ���W�\���W�d�)�����7�%�!�L�K�~�L����Pc�hw�#�m����G<WY��X�D䋂�_�'n*qw�;-s1�;՗;|�(������� ��NоD���O9Ȩ/��a�����@d�����hpa��Bt7ԜF_��:����y
�1�hf�;��U�J�.6MЙ"
]Yo-�s���%�nb(:_���G�����#�_�$q����b%�ՙ��v,����\n_�Ƒ�->ǽ!��ɰ'ݤ�a~C���;�c��3*�6�{ϳ���pD����L���k�t�t��e.|��!�f����2��dx�q��`A�C�ȫ+��3t��XUX�+?����ઓ�Q�T:���m���m��+�k"a���/Y��Q�ĢIy�I���ư�A���3����E'a�41�@j}y������CF!�D0+�} �-Y��Uw6��$�K& ��n�'J�$[CW��&�n6��P\��"��w3N���hC��zUA�I�V��B:�F�3�\�M�Gy�;Υs,'OE���_����1+.D�{��-*��f���)�8�x��<��I�`^��ߺ33/�foT�6�7��y�-^���b#�}t��ys!����
�rm� 	�l�H���B�=����f�8��L`\�P�CևO]���#@���NJyj�&RIVN��͌
�dK��uG��xg���	�TAh�ASt�͒>xO�[h������C�����{��=
������.� �'�>�I�Ts��r���0�Ȳ�B����
-�LDf6���P�#0�\},�(bI��_�n��m�_�8�5�S�����ŗ6�i��;�ELuf�JP��&􄓊0_�,w n�s�a5� |�־".�Ms����e?��֫1���Ux]�|1�6xGB;���X�C�i���V�Z�+�:�H%�y�������(7�50N��S����Na��߯�p�N��˧�U��6q�	'�ܨGs�܉��T�����9{C��3��۵aSi�S������{S��Ku
�FWV��PI���;c=��/]&�a�������fT�g�M�I��7l8)]W�3:����H��Żޢ���s+J%5���
N7n�"�j�ռ�`J � ,ٚ��$�8�3s�-�j��),��X3,pQ�p��L/b��L�OX^��nz4�r�Ļ|K��+zUˣ�m���A�|M;���t�x���4�$8����H�����!NM�k�1<3 �F�T�%��/T�{��S6�_:����p6��𷈶�r���O{o�5��|���ɤN��ߎ:!�p\�B� vI�a���;�A����Y��>�!i��?���'�˵��{�yN�� �lpAB���:@
եq<R��y"�㵑ȼ-ʢ\j��n��H��(����ZT�*��{U�䯽��.�{���{O�I��?��.�E�ɀo��w����hU�[��}�C�c��Z}�\i`�K��?�]/�_�6f����B�}�B�C`�Txm�\�yS�Z{���v���N���3J��2�j��/$X7�:���R���xK�V�k�9�z(���J5H�f&�(�XJ.8�d�KǊk�)E�W�^�.��m�髭�����+��rV�o�ӵ�Ty�.f�
	�6�ͮ�,R؅�t�P�i���@-���;]������r����$M~�%m<H�Rc��0Z��>�Q�,�����A��38,]D���C_4�ٮ�wL��
=�4�to������u����!��:��� a_��n*s6�� �<gz4B�8J'=r ��u�æ�cϝ=d��lǠ�EOtO�cNo(s���b���澺_�\@��"q6B]$�<�NF�2�}\���+��U�IUG��) \��ax|_[-�J��oNI���s��O��m��3�, a)Jb����I�*l1}���Q�I ��N^ӍNL*��H7�V��e�;�j����Ρ��8.dԷ
�k&�z��piN!�ծ	3Jb��@��n�����>�pt��w34]Vՙ�s����	���%�s�pȨ��R���/ָx@���\'�v��H~|���f�r
��'#;�*E�sg_���GU�f����ί#�>	jA�;�_~��,j:BƓ���{{���Tڍ�!�o�5#�DBX�ӡ:9�R�1���f�� ��n��_S!��9lU�2�ƣ���lXj-�:����3ӡ�}�V�:K��w��Rď�*����u���D��o�_7�Ѱ%�]�W�S�:���"��J��c,?�i�<�js�I/VV%v���H�ӧ�[-�曢��ٚ�c
����҅I4�M�˽x�k[{�X$\�Ai�o}�:���Z-ebr�9ށx��P�%_���TyEh�ĲxS�L][�rH˭_�u��R��oq�'��j��R(�.e�Ყ�R����'���ʙ�%���6t7�~nZ�b����0{���rsq�wC*�G�2c��h��fw��P�D\
�tF�-T֮	8=wp�ݭe�2����p��{�2����X#Y+gm�6�9\:��ӾdZ�dK����@�Fn������=+�g�W�߉�y�K"���7��q�9W�E@���-���kV�a�u�^P���x�s3�etؙD�_��ȝ�|?�H�1�)�?� K���D�WYT�ߺ�s��x<��a��Q*���/ �f	ԃ�W��s�dyyݵa �[U�CH ݕ0�������cR��U�y��~=f�e��V���X�\����׻Xe#(.��e���[���9��<��  <�"E�+���*YZ��������j�Pai�%��L)
RE�i�R��:�����
>1|k�I��J`�/�p���>p��
��_d�-q��@`�#fIy�S&�u�����g
Y@gl����G��,�k�Y8�mB!N��V�X��?-T� �}]�Əҝ�"Pڹ?�N�C����OaAg=9�*���z��9!-ܞ��\,�n{�H���!f��f!�^;%E�ڌ���h�0|^>Z2��!�Ҧy&6������	�
L�8�&�l�wzH�w��<�"}����={g���lE���Dg#�@���Apt�����I����P�N9<���k��O�Q�9��v�S����g��a#)�}���e>f�AS�(do��<�wu�֠'����W�}	V�LO|ۚ����6�n�3�$�l�O���A	lt?�a�����a�����%���\��	d�l����T���__%��)��n�H��1���ȉ�ȼ^O4�ʰ�|#��2N�E�e�>
��4uF�}�Џh=��ƙlN�ד%�<�E�A�Jǒ�`TZ�g�,R
��ЅQڦA^?�Zu�%1����&�u�Ͻ��e{n���S��:�<e�@��D�d�1n�I��I����e�o��D����M��t>	�LU�:��'�H��ə�k7_S �*�k���Y=���BC������ͳ~{���3����Dg��U�h=4�����WYTE��P%#f��$�"U9x��5�?�[�PYyE�R�e�F�<ͱ�9v{]an����R� ��9�������7Gz]h�D������^�c'c~��j�پ�5?|�Pנ}� �͖�ܐv�Y�W�@��UzS�V_!8��P#U|�DH��D�u��*�Ы��('�P����&!D��I3Z�"P�V@5�
^s2�8�<�;,�ք5�#�b�]#��SDɌ����9	0h�)/�C�{��֡��E�tɟ$e��(�@��1	�=���h}��2�BGjp��o�X[�E���V������K�����ゎ�ر���M*�a�v20AL�c~DX������;؟Q�O�V����:lXK+0��	0^�?��>ʦ蟞e�Ź�?s��S��KX$�W�{�c��[{,���pi�LV7-��3�$�2s�́�6v*B�o[Ԥn6a��ݰj^o�s~۝���țh��Br�׈@�a ͖`�8]�pm���us�ڽ#	��$�c��yS%��ҝ�9T#!N���\� �ї4ro�{K�`�z�eɒ�w���Я�x텯�S~@��V�'�i�v#�s���z��u���J�TVcݣ���P@�WAMi��Б��`ARJq�lz�����y�	EQ/�V�b�H���8�9h�P|LDs1ue��/N� �x���ߜ�k�z�A"�&O@۵\<��N�qo&��a	;���`h��V.i��]�*�x1Y�{�s���D���XR���f$À���e�B����P��((:(E3UL�w��	����H��T���<��sǆQ���M��v�
m����3{�9T!-$JH�38R�A���V��KD�G���Ӈ$��� a��ϭPEX3Q�I��8sL�e!z	��y?+1/���-���u�� c욊<���M1^�'hJ�MQ5��������)�D��%�^=�i��r�Ǭo�U};MEl>A��fюOn���I#R������G� ��\_\%���On^K�\�S�U��ʑ(�:M�R�Yo�Ҽ�ٿi0���������%"�$����h{ �~��*��e[�d�ۙ��yWj:,�L��&Ӭ@:����t3�A:4m���n�Az#�����w��-{
���V-f���,�Qϡ@��6XB�h��%d�#Ko��5@��[��K�Y�����l��O��$�JM����<�N[-sh9��K��=���m�Ȕ�5�x!pWǀ@/�an8�@H���{���_����@��cǗ��f�$���W�.2�q.����� �rJ��+,����ƙ���~ >S���/�A�ߙwE�2g����y!Rj�}J����o~��d5ms�0%4pu�fuD�?�	�C��M�xr��B�]�zr U|S=����C��^�B���RW�6t��qhOY��B��m�{l��Y�B�pi�4���/П�Vfϐ_-�����������ע"�2�X�Q�0x��(L�̈́gN��J��������� +U*%��6�k�!>�!H*�ل$���������E59�$w�u��i�q1��$__�?����&~N>�b��
pR��ՎE��_�,�X	�xպ���(�i�pz
|#�4�Q�/G9��2��^�IN�X�������m0�:C�1ͥ�;���ż��CxcM�v���ih�A�6ϻhMKk��'H#�
_y�
k��U{�2M�~].�;?�`2��1���b8XS�u�8���)q�a�3z� q� ���%��GZ9������{b��|���&��8�n�àA�0Ҡ���T =�m�s���3�>f����N�`��G���B`}��/h����F����R������r����V�.�Κݦ�6ⲿZq�-�� kn��Q��`?q?dwϿ{�Q���2���C�܀�h��G�=��/}#$����%TN��vY�V��S��^^�B!"�#�q^P.RR�Яe�Y(9r�J�rj�y��AH!�ڿ�ͻ�J����^��?���g�BtT�"���oO:���4���Q(6�B�W �I��2��_��W=Uw��P���*���b�H�j�����F�i�%:F�,��e�7�6���͌|�?����'����q�z������q�2��f�<l�lt�&۫e'�H�m�J�^*ZV9�Ʀ�n��iķ2�y\ٗ�<U�;F�k	���W��$���0ȏ�S�T˯��Rǁ�t?���u�`�U=�o�윇����)��S"Ł!ρf<�0`�����ѧ+~�:Aȓ�&;^y�C�khp���:�;ꁠ�|/�2����_��(����1�BŅ�f�!82�6L�KSH��ٻ�;6j@.*�1D���3�	������@j]�~`
�0�`GG�ܦ<���ܴ�m�{m^��'(��?av/��'�6\�=�RUJ�6�P��h�`3� ,�Ɩ�ZېJ�f��_��&S���Gf�6��U�5�'?v���������O[��uWf"A�����U � 	�]/E�5�41]��lC�	ώqE����������Ըx�n���_�EA�恼A[��$*��=xf��B��U�Ç@N�� �I(�x_/��~��Le��(�9��N���n��壡Lrd]͘3��~;���ƥ@���i#�xV®�,��#�`�PO5��n���)�����(�?��R�a5��TCC����j
4(�,Y�kB����i?K�{�e�^~�6�ظ+mr�u�3L)�(Ȝ�mڲ�v҈T/Hen�Xc����K����b��M��^�~*6*��[�[����"9)���fN��E��X��rj��c«�A�WE�vR��	��_]�Y2v��I�����/[
����\4P�����۷8W�~�OlO�b�8��])N�m�L�/|��.��qK�����Q�1'�
a���A�V���,��^&~qY��nO}3C��<�����x�L�{ᜣ���X9ڥ�����o����v��lj4	S���PU��k��f[���Pq)�f�A B�D4�<K�������ʩ =e�Խ��?����1��[�,���*h璚��%J�+%fpO�diaX���Y�i7��� y�ʂ��HnS��_v���!����g�� �S* ���
�y@��P���ȳڃN�ǘؘ4+�K�˟
�KF�����R��W>��AaT�qw�te�ύ!�'g���}n�1Rc�MՍv�0�l�zB �vr�F\0�D�
�hG��L�A��1�5V VI�l�K���5_�Yͮ��ֱp�{$�zSD�lЎ�5��[̘֔�$}m��'1�Y&:�b�2��`��S�9.��)��#���X.�F�-����1����lf��v��"˔֥�]�cZ&�B��qˇ��T��}u�����.T\��C���E3�ʨ������*��X �(SczpH�\�|����T�X��Q�DF{%P�j�i��5<�E���eb�S�6<��L�I��z�DE�LȾ��ițs_��Zf�	�xS�e�#�Z!�����������b��^,���L�G���R�Q.3%��҃�ؗm>�����߭&�jf)��b<Y��(9"
ib	g��~uY�\��8I<�{��n$����+a=��'��sL�����o���ε��N�Vǋ���<4k��6|ט ��	���c�  �2;���p'����\/j��D�b�+�*��>�4u���]z٨�Q[ �$�Z�a��-��56���5g���jw��~),�_S9?QU��!�?���$Qa⾉Ĉ,#���~s��7TN��;��㠫H�D�m��:��f���C�@;Ts¾P.���:f�vl�������X������[��'i(��M��X#��&���4� ޾{�5�=�1�����O��`��"����$[��A$�ᩊ��S����q�7rՅ0��`W@h9���+�6��ˊSx��/�5G[̢$���Ev�-B���/(�#�q$#��kF�g�k���㞊7��-Ɛ�4RC���)������Xx�]�Gр�R9j����x��tF�&�o�\����>��b�M�h��p(F��u�nb�zd�n_�'	�>��x/3B�i�qJiPK��g�Fn��|��,O�7�8��wћ�'��"x��6��C4�N ������f��"�d��
���I�o�x�Jr�f��Q�������ag���j��]G��6��;��*�(0�B���{��Ւ�cf*B�-��=�FKW�{��'(EG��?�3H?�	�z�8�y�=�� P�~b~���R���w�m�;�y�������o*1!�Qsf�{�4��	+�	�ɮ��%&Zb�iC��a,�f20�\��P6�͗u��]T6����~/ _�9K���njAws�֣���n�����k���~ӗ�Г��Ġ�̉��m�B,�U�Y�U��;uy�+yQ-p4[Ѷ�k`��~��z��hwe��.�v���I�M*�L���Խiqx0h�VQ$x�`�s�J�j� ������� k��k9�]��Պ���{�l��F�9liJ5�6A��ۊ��K��=��ld�BR�^]5W�[ql������3"�/2���Ҕ�a�-p��	OL
�/L�3V�����A�0�[P�y��W��Z����u@�4������xB?%���r��9���b<�k��C
�������_��;9��}�h��5�XWX�����'�%�*72F7=��3�����TSZki��N�F*�v@�2�W�*^����$�����_ $+�������៧���¶�x��^f���9������_�m��
�f��m7�8�2ߴH���� �!ö,��޿d�;i�V���B"#���j�&��%?�l�_T�d� ���#��9{c^Tǣ.҃�b�,*F$�i�4�Ʈs[�<�y����i5��pe��JM� I�{j�>S����5�f��{���j>���r��>J"�t�@���1̌������3a��9�m�}�C�~�*;n9�@9Y�5�� ��e��g�ȉ3a��w���b@��{�8a(�X������'��L��d�\�6wF�~d=.��)��ؗ��� :���W�0'�����#��_�Ũbn���ޙ�$�.��¿�
�� [�#�-���N(��7��,@�Np�4f�������&�.�0=�?�rR�7
T0�6����}�����z�e�b,��o��F�z�u�6���>d�&g��$�w��_�hz�d�@�A�|i�e��g���UEf�nhN��6~��5�[��U�� V6CVkP}�&�ԑ�/�[���uw�mn����/N\k0R����s�x��dz�d6�$7����&m�(�Yn+�Ɗ�t�L��G�>Of� ����!�*����qN�/ױ�p�[���|��d�31D%��TżӖn�#�K���*���E��j��܎/4����(����~�S��STA*�LĐ�%N�C�9�>�i^�Y�c-�7t˱�1}�?�<&	B�4a��J�	��i6A�����!���;})+Lq�E���F�c�h��z�j74�K��=R{��mwN�&��Br�sd���e|�L�@��)�e<*�U5��[+z��?<�N�o+lߓ���pѯ�����ˮ2��
�a�q�`ə���T�L�,�D��&K�G��[��{/�0�w�>!�1����XE��|!+7M`������j8�v���}��?�t�u�xuI���"R�mr4�'Uţ��_|�����<�ꌻ/;�Eu՚�D�M�*�n���{�+X�-��� 8S�10�(=%�H�鿰%Vɗ�+*k�K�8�׀�ͪ��E�pp��i�R�6����l�+pq\�.Yy?n��ǝ����,ZE�jb���1���~�9|#��*�1�ΰ'�4�}�
�o��Rbt�u�p/�&w��;Z!�����Z�!��i��[l�F{/4���z�/�M��?v��	�k���ǔ
��uG�q�R�ఇ�rS���R���m�������]�Z7m	��,O�����l0	�=o���l�G(x� �m}	�&h��.��NL���tI��,C�0�M��?��E�+����P��k%q4�
c�gТ8����d�`E�G�ʰiw]I��t���E�JcLʄА�䍫�Ԣ�xU�XH���_���_�jO���p|c;�k� ����DFI������B�$����8�yj�I������)5�X}�+s1!d��>D��Уi6�p`]�(=����������)���[Oe�hݪ������p�	�O�Q��
��c67����gx�������L��*����.��g�ގ�sK����	�p�߯~#ON�]�oӓͺrA��0�5�[,}�X����Tr�9&���m~߂�/��ȗ�ttq���?A�ͣ��R�R�{X�pB���j8}M�T�N�Z��X�M����N(��nu[9h�h�G������@���?Q���A��0GU�����:PRH�V�4nLXB�K}� 	&g9y �]�Qϲұм̯���
� 8_�v3��!�EX��*�)M�%w@n�Pj�?6A�D��r�+`�fB�{�a�dN�L����`�v��<X�n]�o�98�pD�ؠ��T�2��]�%�6�pl:��k{��υ:��1N�ܕ�H���PB9���O���?P�Z�v�ɝc25&��m�^;5�ִ�������}t����!����;�����n��"�RuE	��d}1�G�4�{�%B�N�c!V�l۸T��J��l�tHJ����mГ���[���t�g1A�M#8�d*B��Ҥ������65a=?<G�s��'���"�CIG�H����*UH��7��3��j� ���c�ɛj ���B�\��^TC�L�����T,�xQ�,��e(��[o2��ӱp��
�{�"'������݌'ԺQ��9�C�k&��H�����ٳ��r��5Y'��~�ȸ��+�� ��4^ϓs�D�/�mfq@���/�Y>�	H]9��p�ƍSe��*,/���!uBxІ�#u��5��Y�ރ
��B�yQ�
��Օ�X/}Đ�2E��u\���ry2^����/����?�xn|���M~�ww9�@"�D}�j���M���ڢ"�_�3U�8��hr.�a�^�~��w��vI��90��6�*u�S�C��;k���m�׃ "��S�/I�����eO��	�p�]���!`�K�,�����?^=l̞)t�GNuDxrg�b�G��u���G'�:�W^lu����cn��V����m��+��*ˀ��D���S���~�4�Y頌Da=mk�W��o>���Ƣ�"�k�U�M�������M��{_�+���b���}�
�J�w���T��È^|�����]�5���\�mu8.��G�j�;�P�a�}���Oe�	\M>�l}H f��� �U.ʹ�]�8;g��q�S'�V�޹���#BY��jFY��|#�\촔��4�4<w%1]p�{42��!D:(nK�������{K,� h(J;�I�{�79��N�Z��h$���	��a��ZӨ$�o�s��ֲ���h$܊�D��b�wc�zpr��!��fB��j&�j�dŴ�>�\$R�� �œ��`=�-�C�G�Щ�mneX��W�,�2D�͗:�X`~1����su[b:Qj"?���ݤeV��U��b��
h�����0�����t;�����!��ƽ�(�%�����4�]?`"7{#�Na^1�%Wp�	�h	$[Yޣ���L8��!�{tPA�,���ҿ��lF3B��!�v�u?�C��G�sgFE���J�Ľ!U ��ڼ��KGo���I�.�t������Z��}�0j��φ?^��W�����x�PgW�N�l<�=�?:OT���vU>5�|�&U�?�+i��V��'7-,�K����5��S3Z)=��M̛;�����+�I.�@��b&���v��y��3��]s��B�\2�c����b�D!|�t��A$��S��8#d\X\�"if#�6�k�E܆���b��T>�^}��v��Y��iE�3Õ�>f96�q��q�_�����2�T����iEb!I��g�TJq�&w���=���}���#�{�������zp���|ﱡ�	�@��s�C���ν�'z�0g-S�h���ڕ���1���P,>Kh2�����E�B�r�����B���T�[��@\j'	�D�9=��G�7*h"��b���ɴ�Wӏ��vd7$0���dF�@o�Ga�)̞�o/���g���&m��y�2X��ڇ���jd�L����ld��t��p����G���x��f����^8)�>��6F�v��Lykt�������T&�1�;��HU��t ��2�K�>;��قi"I�vPn��|�1�������V�)h(PY>�/�
+���L�!Åd��T��ޞJ9�`7�h��l�)����{f鼬`wd�7j�o�.@�4} ��p�ʈA��c�TN�^T�}Hx����GVo����h���2ԁ���|��M��~�-��=VU�#�f�d{�πX�Ói��_Η�����@NFIF�]_����75L�7L������xl4-v��1���w�����*6���q��$\{���t-v�tG�W�D�v�7���ĖbE�
��҃��>10RI�J!�fW45���o����&YK%U1+��
�Ļ��x�j屸��2��iv�F��^���eN� z�A��9@�0��goC���c�ܻ�[�U1䉐La�m�J��
��-�1����]Si�<��z����*��}e��T�o���������x��!A�ya���T��G��ۋ��C_E�{�J1b�����}�=/b�h���Y���題&*�
1��:��3{λҧY��v1b��P(=.�H"�V:�꼜�WK� ӣ�w(�r$ӯ�VlE��g�;ȟ���8�Nh�o�LK����^�|@&�Gh�h<u{�'������r�v[��t-B��]�P��g�[�qBf��%��(�UT<�:�ƼPs"5V�R6L�4���13[��i���5jt�v����E-YC��8��2!,��n&�ܾR��bv5UV�����"1��v��������e�41�ߟ��Ȭ+9���y.��i�y�w�D�
G��`�T��.�> ������*y����Og�$�I0��TsQ�Z�J�ff��j��"F��R%�T�T;~^�jE,����!k��@t`�JF� Xĳ�%����O�52�Mz�M�O�YU?�����ފ�5�+<̠�Ͷ2B=�p�������n�+�v_f,�ª�W+��"�5�j/V�w� 8#ΚY��6@kA	�^ł��&ֱ:������;oZC��
�Xc/O�q!W�b�<�z} ��e �@v���"b9�r-�����DA���<?��*�C��T����ԎO�[a :g�m�	G��X����f��N��s�U��ɩC��I�$
ٱI��q��YGVoo������3G�M�j��}���	~Ne״�|�{�hjDeQ��2q6v�w�K�#9���UL�&`��u��4c������k�,����I��`B��J\P_���]��pg%�(�Z�ᙟ�Q����_�8L� �]9����S�/��S�A��� �I��^<|�*^ٕ��ѹ��/��aQ5�O,-���89 ���[mc�/��L1,�]*h(�8@A94�Ȉ�Z+�a!��j7�Q�T)s�)8e��+9���??����Dͼ�a��me���a����=c��ӥ�ζ�($�|,;��I�/ӡL�E��5�>��n�C �����
�w-�zά���1��X̚�A���2^B���u�C� �8��bl���8~�Z�@�3`�
M�����cv�� �:SMp�)M�%�=���FH��ѯ10�<,x�=~��I���F��̻7�Lc|R~Ck?Ҁ���(у��y�|V-S/5]h�»p:l��4�D��d8w�!��U���-��DR:5@Z�L} A����W��o��k���9�� Uqɑ�Zɼ��╈(�l��u���p�b�x�����I9�_Ok/)H���b5�%)=�b*3h��+��گg��M.a�'>bD��'�S��ؕ:&J�5���a�670����s�O׏���n�`��y_n��LǪ���]�:��0RFHh�K��\����j����
�r�:�� �4�Cy� 9!}��߿ڲ��n���"{�M�ޟ����>�$�AL�tXq#2 �z��Or�.a���N���S�r~���N����G� GNiZG��`�y9N�6��*��_�'�}6��8�h�B=|Q�Օ��������
��ޓV������>��|�� 0Hg�<���EӁò�f��<i�as��QK�� r�X�0{��\/���{\r�p1����Yյ�a�<Yn<�o�����Q&>((	ϽDk�$���B��А�k���dgIx:w���c��A�EP��,P�rUFH�u(�fX��<'�C������	 >�7�pfb�&A�yр���"j}�������q��(�]�7\u�9J��\b4x�B� O���̙|$ 7�ݭ��Zا]��ȁ����B����~��S�uKwo�ZeS�;�c�N0B��Z�TdwT��b�GӐ6]6���*��=��Imşh����͍��A�(�en)q�i ���P`6r�#���8y:2	oI,+�i��'`c�+���!;ED�3 ��υ#���IdJG�8s�l�or4���gQ6Q���`1�~=tP�Br�"��"����Z���g%��~�LB!t�	���N��l����c-2H����y�l��M��G��p\�?�|G�Β��;:Wά>܂ܻ�����e�;蟒j�8�j��f�����mD�C�=ݮ�8�آݵ�W��'N�(_���ѿ�c�ަO����vT� ������RiaX�JD�\p&Ň��ƅ�'��=�v�D�y��6��JD�;hz���H�aŝ�>'o��������P�a?���'`�m2[2HwK�0,�����]��u�;�{���W�\��DY@F�� q�>����~�--���/%�<s+P��&|���m�$��[U�qT����8�6�q��NR��㩮in��候o"n��6ʽ'��n����i:��߀WZ�w��E,�u��\؋�j�����s�'ہ�?����K��
L�wp�q��0LFڰ��"��_�%}����r�5�4�Y����K{�y���d�W�!R�ҟ��*�S����R����B����:�\<گ!�+�&�1��6�$Fo\k���x"��= M�ԐC��k��P���f�Ea��\U�1�]e׫}����e�SA%&cB1��`L'H��F���b�Wmb�O�a*f�iO\�B�ŀ@�9���{��wD��8���\s�/�T��w������h���zp$����P��٘����m�L0~�Hl6_�b��h
�&qa�1;J�
*U$!%��7�v��������;W����M�KD� ��c?�A&�'B��Job�$	gزz�5"
�(.G� X�^"�(��_��3�R�����ޜ�^�o��8yI|�Wy;Xw_�,�g���B{r4UҒ��Y��K�W ����UJ�۵����,�<Ut�����*:��lL�p�1*����&@��}7��>Ӳ	���<�3���\�k���� �LD��j8�0�����J	��Y3�\'5r���[��2��n&��gE��=?t�9}"�I�����EE�s��,��&Ujo���G��^�V쎤�9tґ>��ω��pqt���G(�5���<�ߌ�p$x��;������%��kl��9S��+�Ǩ��.d=ƞ�r�Ï�<�Q�u�$�Rzs���Y1��1b�ǃ�7�U	����j��*�)�G5*�	_<z�~:��5���2�S�Z����$�q�G���c칞�4�S�J��X�Ғ�;Q-aV��8��IqN��m��D�8�qؾ�r�@(�s$/��WM�l��2�^<`��e����[��l�9�+�A�x��#�
l�s�^����-�2�/_}�e����o��,>۟�z�HNs�+T���;z6v�9%�����du'8�ǒ��)=Q%!��v�^%1�^�Z�oD��Q"f�,|l|���\T�H��W�����!�??�1��x���nQ��F�䆵�`�Ԇpf����gž���3�SFs[�}j����씊Y��&��v�W��1�.���۽��Mv��͗���'��L�� ��� 4�5'�t)Y>��V�����N�oNH��O!;���7_%:l�a@����ĝB���XH���{���`�����q΃Rh�i"�.�ϲ��?N.���sv)lnZ��h@Ģ��%����G�!j~��I�Q3%�C�0��VD2nryW����p�p�R�8Τ��<w0��m(�UDt�ZD*ŝ�����q@"WיּKK�_�hĢ�UK������ti�j�Y���d"�&������5�&/z�Q2;ϼzX�yF��f��m<Ȝ�̬)��#��fN��ʯoY	R�!��Q�.��(���a��<�%�m�>]�WABYюk���M���Ғ���:^mui֞. ����.xf����dv����+[��o�������8@��B~?��+
�G����m��)H���n۪ (ν
q�J�5c��%��l�vr�;<� d�U~�+�i{�?�*o�_nn�9JS|�Xu��7Ch���請��Q8jS����^&�Q��ys
����>%��Bnw,Њ�K$�{�:P?�M��	�SC�4�@�Y�Ǻ`�p����sL�_O��㜮����E^
�"��V�6-�����(u�5���"+��$���k(���D��5�ϵ$m0��~��y�g1����\{y�$c�-�ds�Qx���|'���ڐ�7����-�wi����Cj��5�$��&�8~EQ,�B�Y��!>o�T�M��q�3�����+]j,D��kT|�AV�$u�	��W������X�G��F]=F�Id)yj����1�H�"����l�2(��>��/��T��&���P�qN���X�ݲC;b�	S�U_�n� �6g��6�`ۭY5rVu�&t
����IOӏ�ݓ���G��Վ�k��E�vrX�A�}4e����?�A�g��D�{�ӥ�uX'F�|����D`��D½0G�`D@�>�0R6E��vŲ�}^ ��T�K0KD����U��UL��@1�e���Თ~�Ϋ�Yn�޷�څ�*<�Fo(���0?-�쿍	n\n�wv?���l�6wk26|b�u��b��b%�p���S�r�N�X��o�?�t��V���)����692�mޒR=�oޡ>x��,�C`�Ag/��m�W���r-��urWO������&��KԞ���tc�Ӝ�e����i�&�d�sϟ3���R�?>�Q
7��d�P���X�I��Z��R۵����=`|Tǵ�BO�K���\�<�~�3��o�*�b�Z���0#�3&v��%�JBD�z.*?���vj�*��`~+8�ONZ�/�3�q����Xn����ИY��������x4��c���Sp��u����"��8����Q�������0�]�Ԙ��s������:Zb�+��B��$��� (9L�B�s��� �:�|��z�&�]JZP���u������\Xr��;�bD��Q���:����!&�G�Y�+�LJ�5�4E��� �>�_��5"�*���W�W���1�M=�
����S�:u�j�����H�Ы;�%��U
�!?ӵ$ی.�~��{�)�)�[0���R�������X��u���0��(`0e��f�S�rm�	ȁҕŃ|Kh��|��$��_�L�G�bI��`� 
N\t��j1&�7����z��E��ӵ�}�p��.�[9c46,W��6wW1CsO�LcS�JY���]{������*��yn��QfGY�����4?-�H3B�*��)j�����ɻCi�������?a�AƯB���e�����«�
\Yk�c��?�����H��
>{�!�$�w݊b�@�R����gm�ݽ�T�F����.�a���3�g��d�� �(�NA���������=�B�W����v'g��bS$/����*&y� ,��C�/  �`��F���2�ǳ@����rC�Z]�W��<�67�IG_n�$>��C\���)� m���� j�2����'�bY��&v�W�?��jE�A���e�|Hr%�\/�h}:���@���z��;� 3�xӷ���T�~��bDc�~�4�i�򚼍�?�H���ӵ>��b�d�]q(������d�k��P3�|�̇5A�n)k�8.���i��TIY��7�o�4���2��ƠP��l�^���O]��t��'��0p�W��ˆo?O�#^�����ͭ3;rƟ'I��~�na�����AŐ��Soxz����t�%G1�pvo���mpba�W0V ����Gj�x=�U��ʜ�T���̟]���w7l�CV���y\~�2�IN9����<u��GS��Jhȥp�@^{�p��RI��������$��n�c�НK����Βn�'A�vv���A4�fx���e�� ��c���8 ��p��7voOؕ��;���ވ�fZ�y^M��9f,piS�R�U�q�d���(́`�)qMܭ�����y��a2u ՝n�*$3�0.�-9��R%�:�NϹ�d���1'	8ӥJj�F��L~(����;��ڥf="�0��؞}|�$ЂC����N�(��c�П2������?Y�ՙNʴ�~�ce��wK4,�Lt1��C���5�v�>6�+���<��ɖ�Z����Ȅ"�f���iԹ]3h�#-^��e(�`T��� ��WES<��#Ǚ�����d����܄�]h���+8q���oi��^�IF"�8�Xͭ�xB1g5ʆ�g.�B5�i��7���`�U��N�@-B���f�m���8��r��-�J)�Ӧ�v��}ђ#���z����a��[ �3\�є��Dƞ��}g�����ȬU[)PU�:�d�wE飳 MJ��Pg�6ڽ�>l�q���5����9�|���悖��I�ӎ��P��8��L �q���y��h�k6� �������O�C#���������<�Ӏ�~	�L��r��U\�r�u4�_�$ǣܟ9y� ���zۦ�4�O4%�	��MS�O�����05kP:]6�2~5�z�h�ા�c�D�2U�2[�)�(6(PbVv�$�����\/E 8Cҹ�Z�u�!(�U��mu����[��/ /WFT��� ���6��q�n��&��,V�J����MW�!�"�)�p�ͥ��'lE�a�Vo+�̶��	4[ax��U]�	> �D3�]���C���]
~�^��:ۑjR/DOJ�ɴ��Z� �6�y����T9��d�`�
�D���NO�|j���i�H���5_}����vꈄ��ED	o["90bЦs�Yx4|�`�o�	Q,�k�sD���=΃���@� v����M��;e���-�5��`�����(���#�X�SI*���З�����������,+��������s�4����% q�>+�V��ŷ�R^Q-�m/y�����"y
z�����"
�-{��ܷ��Ox]��~3�����h��n�����4q��l��Qk�c�db��$)�Gx����(BcVJ8E��U�E�W�����na�D9\kJ����P�k�+&c�1��)fm�6�2x.o�&ǳd~;F�CUZ}i{n��U-^,h�:֞�	q~����^��z�oKLv�q:���ڋ%��2.��x	R�5S���F�U�x�r��N�go�hfHhDs�0�j���(Z�2DHe%�1(F��",�?��Ez�\�&��0֣�;�SÏc.��Ѳ�#�^?Q������)W^ط(�Ϗ7�y9���ɕF��I�@p�ex7V��eK�=^�G�ĸ��ڊU:`���,&�
�p|Pz4:\���Zc�D�%fH�R�$7�.�_�_�w�E�|J�E�+��N���ƈ��f�!�z��M��R��@](�Y����K�!�AS���I���]E�I�@��u<�e�:�=�������N�e
�L�9��鳔�G.�@@���IQ	�x�"�y8"�� k!OQA��4�"=?����j6�'#01#���qA��g# ��@�~�S��o�H������9z���?*�;.��n��h��h�֍�!Qp�\�W���U���\���qF䝻:����vv���$r����͘\u?L�{�Mo���P]S0ɢ�"��'�^�X�z%�OE�/��(hex�A��g�����h�q�XU|�T�p^Aq|�y)!
Κ	�0s���[�_��$̲ ���XR_��ݑJJZ��a�	iY��h��t�Is�%{�LNtĖC�6W�m��~��~i-� ���`f0K�4�����θ���Q��H0�#Dr��p�*?��IR��9^[C-���L���mL\���@�K��g��4��~D썌��HytC��I
$�ZI�k�
��O�Hg�Rc�y0ˍj~��gҚX��b�9������*���6��qc�eU�P���"��9��E?v���*d,6Om�kmy����X�hϟ��;(�ū�F/ti*Ʋ`�+���xe�g'2 �������d���.�,��t���Lv0��+����1�}�*�{?lZ,����#�?���dg%�26l����X?���WyJ浥V3u�����W��w��~hH0^�G�X���k-���d��!�pDRb�t	��|� �;��Ǵ��B����0*̌խڿ���"� ����`�Sy-+|�(P	���8�hg�Ϲy��&��I�}Go=F��"��cͬoh�Y��z;�TLhX�OkrD���FF�h�$.y�g:</+h>~�����P֠.`��E���g�6�l� �b�f[����y����|Z�����c����'�pm����i�|Z,x�����]u�u����#pࢅ�C�P���*��s2e76F��h����1ŕk�}pG�Ē��{�-�/��X�@��cУ��-d�y��W���I���t"D�~�����T�ԑ_�3�\�}8ؐy*+;�U�@�2�n����}��'$���2{��m
�C�?���}��.w�a7�B���7pz\��1IԽ����{j1�اL���~}8�999�	橔�y6�49�/�^Q��H;�ab�a1<��#гw�%|jE�g��ƽt=Y�F�����(��(���mG9����o�k�V��.��6W�c3�IvuR�8�7�V��1����"]#f��j1	!�7�c�C���D�U+��)�d��B��F�x�0��bǎ.����٧�ηe����~Z��F��O�'��_C�}P���GD��D�s7 I�C�ֈ������=���6\v �
/D�t�JtS�W�R@"xf�{���շ�����l�֩�c�d>�H�g<�љ�;�1������2���-[X03��6=�N8�v���%�g�WM	�q��3��ԋ�*���]iR��N�n�<T(�<m�$�=��g\hL^M;�s�X#�IK�z��B�q�J(X�M�~��kf���rqU�t(�������I�Ɣ�Z7�����vǻf�L ���R��R6�E��uPV7�k�b�LfT�{O���G}�YX��a<^��Z)�
-�x��I��I�_��.Rygd�.(jN�I���s�Ab}��w�nsq;,�V������3�:.�T���&�+f���F�RR��ֈ0]��E����91ᆊ�ɫY̊�}����v�-#Dy��M�������Oz���4�W���v>�ʞ ӈ_b^#E� ���K����������q:���Fx�{���s��g4w�'4b�������@='�����H����n��M����v��|#��<�.霰����˃n	������g�?&�J�Z�0�C$g�֒Z0���ڨ���T��O�s+`Hǹ7�5ډ��r��/��9ɡc~�'�L=E�7V��=�1��V*�E-Ô�8�K���+�C�D��HP����&����b��"*���Cr���U�d�)���j�lڔDQ4R&�i�)��ҧÊ����1�K�۩bh	&��I�&��Q�P�J�)���:�LW�ez���*�N)F���,���FRHyN�k��x��:�_�T 5B�K�妕l2淘����r�6hށz�nW̍vE�%����^� QraGl٦A�*�7�;eW����eY�J(\�¹�{�UE�#9Ş�	%��vmK���a댹hv�9CJީ�q(�\t�׮����wm'��""Br�	�zN�龄���#k��t�HS}�r;V�^ j!(7�Tkոǳ�4�4��5	)a���qk�ǡTE�M��_lL���n#�0�: ��M0�tK�"v�aJ�C(I(96hi��3u����g�k�E�_y/ ���j�`0�!%4��h�N@ ��c��jK�U*C�c�˶.ݭƿ����2njhz��xz	FLy�YB&�A�Ӊb:��_,���ȣ�x�3�"��\Q�Pl�!�R���������>�!i��We��	����K�8QM[ȧ�GGeG*K������5֝�{�$N7��`h��A8����[���9����#@z�A4�X?�O����=��T�\�[H�r��'>O��ʻ��OV6����O�9B�8i�?\���]9��>�ţQC�
�fզ��7��o�2)7>����)�����V���M�:�[��`<�g�m�$-y����S�������u��]��{�8�p��)�u%@*��b����,5�ʵ@�]5�O�^��[T�,}���r���=Hc�6],Ǧ,X+3ԇ���*.�2��c	���(nv1�h-��&��2��g^���fᐓ/$�t�������
]M���%��+����Բ�e��YF�дk���~�yj���ܷo��~<�)�J��N,kIF�%�m� �/��j��X�/c�y|+��FoZP̭h�#cq"���âpt<8�Y( ���!S
)��:[U��?�ʤ�oa3F�~"�'������č����8�������I#�il4A��?��������7)�x�҉��F05�u�˗L�s�d��;��'tZ��x�H��� +�e^�&���\�hm��CU��2����.�E"=�6��hDa��Y@A�L��,>j~8`�@����Ő1k�+��*�c�����fq���i��&��q���@P"����cG�+�i�D#њN�d�ֻSO�8N�n,ƾ&��U���ҖXF���룹����v'#d�DP))���`��X�`C�~�/��u��cU���ȴG�{+&��\��N�p��t>� b�Wj�0
�WgF��'d_�\s0��'T)i;�i�n�gT4���4�t+������Q{���ra��J�8RU2#�?iߨ�r;�����?�%�#�����aL�La�<N��v`���)�捬���$����܍���'����qCmQ��U�cǢ��>�O���׺��3#{�O�N
�i�(A�k�C�R���4��;SEw',ӈ�CR�*J���˜wElY���>8Lϛ��m��!M��*����H��&��6=n�*y�xh)�DEK��RD��4s��n��ߔAw�鏒4�C��ދ2�Z��5�3��A[.��{O:d�c�X�g��������<������p�L���_�z~�Bۉ���Q��ڜI#ãtJ|�A�� �����S�+E�Ep��w�팰H�4���^���n��i8�Oq��k� 4~,�9�%�.=Xw)�E� ���J'"�[��?�@����u���3�?Ed��Ŷ��=�����+2cȪ2"�aJz���d��竼I��&\ߤ3`?�����Ǽ"k)�h<u�K�:��^�)��o��x{)s��Ϛ�ȳ��'�a�� �<��ݻ?V�5D��b���t��rp:�?�dY��a�zp�ۃ�a`�of,���}�ȩ����f��
W=���X
�1yLߴ(�o�[����Jߤ�j�O濡(��Üm ����iQ./P%����b�g�l����Tf�]`{�s����!^�gU|�ݪ�3���|K�G̚S��܇�ɽ�-�`�,�s��C�g(��ҍ$'*�(6�xf7��aM�K�{�F�FWA9�}�	��,Jǝj=V�����(���kLY���տ�[O��n���7rZ�4a�'!�6�����,x���B\t2�Oc���A�X�驇 ۩&Q�^H:s�bW�U�zeF��֚�3`&�˽̝K��I��ga^[���C�&�E:8D>fCHJ&��?�t�5���h���O!�n^DVL�4���p���7ӆ���y��t]x)���KHQLQ��q�N'H<��K|�r1�;�c��'tI�����W#�M�"���ȍ��E��Iɘ�x�o�2L)romiŖ� 7@��o"�VH4�:�����_?�˦�=?��S�H�8��a�K����
�0�u�ؔ+�r=Lڲ��b�Q��m�='�-l�xO��^�L9g�Ǝ��[�/)w��햱��{�Q/V$��-����,�F�[O�ouYd?�lpbX�c	��݀�.�Rݢ���ͮ�DV���`���q8��-bw�ƵJc@�镶չvh7>�^%��;����bϼ� C�ho�$.Py��=*��ܑ�h���D}�eŵ�ЯP�5J^����e��x�$�/�mUF�>��(�-�s�/��0�O`�G��H�& z�[**[)I?gh3��R~�ƾ:#/�T��|X�~�Z�6�?��<-�&.ח֣�`:$�Fص�	�2Fc��c���UW7��&7K�c��*i�� �}��"��>����H
�"L��4�Zd��O�y��3U��(�uq���{eA���N@0/s����wt������l3q�ۚ�2��p՛lőoi��Z��y?D��i6w���z�h�bh��e/����`��}q�*����=k���\_��%~%�"�_�Vx�͵� ��K%���|4:���R�T ���ط�W��$b �.���*��R�n�f9���/���]��D4Q[�#jÏ�bsDDQ;l�W�t$�r���S�|�7�y\�6�&!��[�T����Z?h�^�%��������u��?��Gk����{�!���Bg�k�W�1�g�T��.�	~�0��M��oQ=9N'���
�i,���zP�yv�y��Tt[SY��Io1�6\~/+�x��@�;ʛ��3P�:�Br��5ꌰ�C6KK[��۵�4 Nh?��I^M�_/Yb�����c���@3)'�J�y�V��֫�9�P*�u���%�l\	u?A�P[�	e�ו�D/m��b��o(_*���N�J��ĪhPX5@�X�2�!;���]>��,��O�ܯ�"��hٔ 5�'��+�����;���S40�56�p��gMЦ�la�}g#E�݈���#4�B����q�&�Gϱ[��kc[)�A�,6	���O�o{u�:q^�;������*U ���l�Y�,k�;9�^� x��n��N﫢��R�m|(^_�n ��q�Ր��/8�r#Fg݁20���8�*����C�,<R�~�9�|#�����,G��Q|L� ��G�F�'fXn��Q ��X�XXo,�Pީ��NO�Q�Q�t �=R�mz��-��c��1�0�e�
���Y���i��敧־B�V�/���:dI��hZB�3�N���h�ÃQ�[���vtG^E{Ջ�8"��ߟ�E�KIP.��ʉ#�C�i���?��SdJ��� �ĈL��������|.ZqS�����0]W��+����-o�r��;t&��xjɿ���(�뺴��]X�ra�����Ec?w���j?r���_��E����+�$���S�sa�*�hfVrVRJ����Jq(�I�42��J0f(ώ�G�=��+����9���W�c���:U����rb��/����+ZS	ɲ��W���.�>8ֹ�^q� y����"��c��ɡ�|,�����C��H�F�c������Tl�řd��y��o�SZ���I�b4�t�yin���5!Q�v�F�fD6����
$�����3Ll63Nʣ��~� ,�K�V��0���v�a$zV��&k//S�s�7T���D����,�;�t�i���e�p�)@�w�ִ��(F��ֲȭ�:�CsI%k�j����**3wǮ��e�kx���)%��l���b5� 遲,J:O)u�[l-�����5�J�:�$�������0�̥��C����e�C���Y��'{���ATb�|n����n4f����}:V��[���S�g�(��T����f��s_�d��j8��k�ص~�����F��ތ���,%븆5ֲOJ���m���`�$��P-�9 2��L<�:�?��",dH�>�w'k�O{����0�${QC�`Y�x�w�B�A��b%��d������Xh�*����az	QD!��	��� ��
g��|�wZ"���Y���l�J�cMc��:ܳ���Rx-|0�H+%_ǭ��w�<��V̮�p�n�LX(��du"��4o0�BD`zf�=1�$�+���Tct��q�k�����'va��+�!���I�73<�.i�����0Ϥȩ���ӯLI!&go-s�=q��ML����w���l�]?�#!��BDW�HJ����֋�S�	w�F )�p 2�>h`�4�	�����6�>`�ƹ�.i�Җx�����a��g����NA���\5��Yr��4�
ɘ�q��+p��B�����^"G 
6��}?��)���^�����X��C�ۼ�H	��j S"�)�#�V��H��2�9��!2�SqF�
��?@��Û)��^A~�}>d��f&��GJp�2�kЌ��t� ���D�T�@��X�����Y�]̄���g���.���V���0 ��()o��H&�H��h�ܔ_�q�_)[A;pFP��f�JdC/)�;*��W�\(�q��ȍ��\.�m5=WmQR�&C�<����������'3�Z�M���gB����,�\��6�<���\���V�I�tK��$u�XjrA�.��*2�?Dx�,�4����J�m�ob��HXA�^��P��q9�Q<��qL����p��,:S`gI,ů��Z��n5�����+�����H5�_�ޓB���خ�92��9���*y8|���Nn��ۧ��bU�,���[j:�!��P���/���nBT�s�0�׌��"5ɛ�/q�Rӂ��N�6����;��u��$2GëPp�������gAuckJ��� �aq��W���J��QX�t�0��|�ɰf�v�Qz���匉{W.�NYc�d���R<̏�v���H���l_�;[���Dy���hq�>����{E ���-e.�x�'��$�dB�U[��4��Z=��<��|�>�(r����L���d����~ vsD�3D.�C��*ݟ��"�b�'�:�7�1������M8�JO&���럌����������]�����:��BJp?wH��P�^��X�x�[��r�X���GI1���$�&<��%�U��-���݌(����:�Z#��u�<��_����q���n���k<��>*i\-�; �R�P�(���:)�t��kJW*��h�Ҳ�!�?	��@.6\�,Il�%�p͌;���Ǣ�G�HQB�Lg��q2e&��X|�����b=�GS�Z�>���.���Y'k�k6�iړ��`L;6�<"��'�y�%��<�r:ު0�~�P�Р�,H����9ek�ׯ��k��m¡���7�O&\�D�Hr��g�!��ٗ�a|�����XPL��)\��lY2�ɔ��40�
����W�<�`�x�G�q����J��t��@2>ό�#�J�����ז�Z==����?;�����!,�����F�$�8.D��޳H̅(ɎF�Z�	�� >��J�����J�+����ʙ�Ȑ�M)c����V����<��x?�(l��{)�
�KI���k��V��DS����B}5�FB���^���Ha�ٷ��A7�֍�j�	2���Q��^��
�x��˂�zln4������wv��2%R,���_�@"mp
R�B:��Y���;y5����%:��K���RP��tor@mh�����S_ʌ8�X�����`F:9�O��!Q���f0	ƀ�B2IX*ɽ�b�ճ��ސϠ/8c��S�jcL*v�
$�q�WI1�w?���5ƈ�>ڂ[�`��"�pN��%�� �N�Xt��&R�ǹ��n|%�-�~���v��t�*��#5W�**���'�UH^;s� 󦮥WO�����fn�9<D�G��U~�B?��{kߧ�k�1n�7�\K;p4S}1���H�0��?�r)َ~�DAT������$�*! ��t�������`�ĐhL���>/W[�Щo�ʱ⥺�19���n���\���æΧ�OAm��CG6�cy�CVE�֜�s�����|$���v��
�eK�$c�R��C�@��F��=n=����mE�l���}��Q��SF��#�:C;(�zU�%?��Uȓf�Q�s�������m�^�J&��`����ʱ附օ���U��
nrn2� -
�6��3o{�����<V{P�;��xzE���'c}^�C��M\�H/�_��]uݿ�_�U�)�^|c^�=�z���@����+7`c.G�R�����ed��4��׋��A�V�;�K�dMf`��*��cV�[��\��XM-�6����?utH������׭x]ܟ��Qd�o������>��^�ǲN&�Q��?��2� 7��̀7�.5�餿�����Z������1���*� ���v���'�z7��̄~?O�������� &�v�|y[^LCplu����B�}2��|VN!^���k��ι[��c���P�g��x��m��oDC�__�N�མ�{̕Ǡ1��M�<��3�ͤti�7*`�9���^�O�{�	F�m�Yb���­:��9>�l@�p[h:Yu����]E�<ڦ�X��o�Q		���J��-O���J �-=${��`qŁC��@#�l�����*���#��5۶�3���Jȥ�ބ.(��5�!GP��5�+����p?�$RČ���������NZ�?���剮L���V����C�섬V��k�0�sr�t�3��s�8�g��"Ω�;�o���BC`/U�ɽי`Uh���
U���,�[��-u<�r�*��XY>�(ȀA�?W����g��Z��#�"z_���hWޓ�!�����sWҿԌ:�%F�ѩ������T�Bf�����˯ޘ���;q���p�M�}�FU��g�ϣH��NR�R����;;�K* ����\bTӦ��f��M���n�_Nı�Fg��?�K�Y����P�����:��͔O���o�ytF-2����PqV��`X-���T�?�u�:[n������#4+[|���4�F���9\�p���
")K�� x�Q�BMI7\i'v��k7�C�M�p����z^F>�X\�Y�'X 3��q�b�*.�D��RL�)�C�����[��rK�߱����Dv<�jQX�S����f�^�ĥ��Bn�7U6�z�^~2M�|�w�.]bRZ���9b+Dܿ�j�:P�O��
��P�IL$	��W�YQ���j	jU����̰���7�@�f����Ĩ094���W�{T'�j	[�Y���Ap��@mXEb	�G3�=�c��SZ�W�.<l���t"S�6�]y�� S`���۳L| W�T�:'��S2ȯ~�%<0ⳬ8�k��xxc�r��x�B�%W" i��$&�0���h[́ru��B����є~4Տ��6��pF��B�ŗ�_�َ�n6���z�i��>��(�Ȑv߮c�� B1Ƥ޶�y���bJ��U�`l�LtʆKT�ƍP�ERp��8�=�H$��ّ�CV>�'������U(����h�㍧jo�Tt#E�wx� a8�����Q���}��"Sd��?_`��	dǏ�ѭj��@��e�c��psظ0�Ǽa����>+��c4���㭈 P�=���|mu�e�	�����cbA|ǽ'�R�pC�?�Ú�&+X��(]�Uř,���Ġ~��|{>��G"��13��E����2�>p�p�Y��I�Q�p��x��tF��?�*��Փ� ��补y�=���'�1�����H��<��d�p�y�:���AKh�W��Lȋ��w��.=��x��:�l���ߘ�X�s���5 l`p�gY�i�,)p��S��q��ӳ?��ˠԽĐ�s]���x�oo��G��<>Q��Ɛ�Z�9�3�s�Zx�/�I� ��Uf{D�{������y ������޾TD�Ɋ�E�i����AJH���z��aDצ���%w�a8Ƥ�	Z���\h�U�]<�H�&<�b,?�f��4� e|',�m�k����w봃�᰿^��r	r2���י'���|��O���������j�7eReu����:�r3����Oٔ!���/gٿ�,|�x+�dXN�ʐi�|+K�@J��Ox��_��Y�2�2�\k��4s)̜�paF�iA�i�Bl�[Q�y��I,�2�����H����������nL�g�%�z��{�B���~5;-6�������Lݶ�)4ƻ�3$��d���q��;a��`��!�	�z�����ף�q�C<>=zSVЧ�^�5>9*��,j�2���Qt쐽 Km�x���J�y��T�dv�s�u�i+�ca�jn���Zm�*��g�B������b�\��H�ۜ^�b^9� ���I�Ztz_u̵�r��e�B壤���n0�#kךIv�O���뢱2X��W3�/����:[� \��T5"�Zqf1h�3��]U$g�0]��2�qKwWV�t��K�U���;��r&��q[�Ĥ�����M:g�T=@D/���$�嚸}>��ZjgI��a����C��oQs�'�Y�2g��2�*{Nb�Z�e�FYp��d�\h^L�5��b�0���-~��e�)�2�l�W�ك.x�<��v�8�*RB�|v��~��r݄�n�@�����	�UEp�v������p�F�[�J���[�9)��L#�)E1A;<l�Z��$��諎�<g6s��X^�Ur��%�Hs�l"/~�͇���l���7|ڧ���3f�2X;�$�vR�M@Y��'�MF@��S�D����D���� ͱ��[�&o��hԏ�L�*ZU�?��I˱m�j`NOL�5!�YR%L���Q���|�d�IOk(~�|�%�0	�+\��zϦ	B�.q�OJ5��X�Q؆��P�N^ུu���dR�b��n���+Ʈ��n��.�ϓ��o�k��YX��`����ow������:�.�Z�`gf��$J�5�gSxP�0�T',5�3��s�.�靸g�&��(w�`|���Ly3�4b�d���mi݄��-�n�+{�ij��P��y^��P�lQ1?�p�o���Ai�~��!���6H-��|���	������z��)���2�#�U���,%>,�Fd��v�F�yԢ<)��L�=#�Uʟ0:��.�37��H7s��u���>�G����X�T�:����#Q�4f^��'�G@�$li.��-������HN�J�)���f�h^�W
�ð.I�~�c?6���^[���;�:�Q��7Ǳ�Z�\\��a�tH��;tMk����&s��d3��ž>���7T#����K�����
%�=��k%5�Too�L�}��W��>[�t	�X���/��8'N��I���JH����jy�It�]_c�U>?0�L��b�����+z�1C�#ҵ�����ī%kȰ�Q�x�݁��5�e��%�&�{:Kx�%mvX�>b��6hB<�TR}JS��>���kO�_8lR��\W��u�-"�6����W��# �)-�m�.���¬]���u|갽r~�,��i����w������nLGs�Z��#�n�T$�㑴�1�����A�h�D-�ǘ��*0�A�\� ?���WUhT�BWq	�`�E���Nw���"m��\����x�^���N%�H7�{W��l�i��bjj�|(�:NpT�u�@�u­Z�蔜��xu�e�!8>9@��A��p��1wnf�F�m��C_4�)H�c���"�#1o��B*������7.ʮT`��I7�6�t�O��o�؏�i'&�:��#893�;u�"�BʓC0�A/F�1$�j�~��� �J����s�Zv��"5Nb����Z�Ś���0nL��Xm�����$	[:��� ꩆR�2>L�Z :�aN]��'�P5�2����"r-���*X�t&�ئ�T�����h+Q�V�ntI
7��]�s�P���2�My��wEUM�����ɜ�e$�5�#s;��}�/�֌�"�ўx�npD�M��[��E�����ȏH�,C�!�z;�Ԫ�~�Cc�j�eQ ��v)t�I߂��U�P��'��f��K�a�]'�AT��V��sI�>�6��N$�}<�P���hE1��P����`E�J���**��G#x
q��H��E�cK���yux-L%��mp��F4�~�K�3|n�f��#GְtJ�Ξ����,��w�׌Rhf�����T��$	�bu�ɶ�h�~��.J��%Q! �R�d`�>��\�	��k��
 ����؎wcWzs�oo����d�.�� ��,�m��������.�.1�4���8������=V��mp�zLzb��	Y�#u�h�MA��A�f
rԆ 2��m|)9��+O\߂f�N�t����$�&�������!6�j-}i~�T
�ـe��ib�"���VB��6��"�\ WRh�Ĳ�8��k�V%	�E��غZH����݌*���:���P@��U����@J��]���l/���s�čF���!����~1F��������{����F� ��7�D9�e�Q��Կ�	]O�%�*Yy��r#8S4���[�~����
⒔�b�^�ל/4M�=��D�E�NlƘ;�N8`��L�6���Z��f��ɐ�m�=�w���k�wB���9�Va�'�r���@ќ�Ƭy|�m9e{c����	O�T;��y�V�CleE~��L���`�gFC):�����з;b5sd�/�=G��4��� ��DPt+�m+��6�y���S��p�a��� �ё��]C�D�v��dd7��n8M���dR��:��cv*פi*�>���̖E�~���$�?��+�3��g��9d�H �9~i�V���6���(Q�v����ׂZ(�j0�A�A���������Y��a��9��UEq�ZK�l#�$?t��u!}
:�7��Ī��MB�C]����N�c�?�+ׂJ'�~��$�9lxp?����FB9"�Q�J�ƌo�j��b���>/�I�1���d�Vg��}�G,l��i��x+�u�evV�X4��@P����]�]3'ySu��],�Y�]�U�E@_,�"��C�6S���nV%"��!�g�,X����dV�Xڿ.
��г�K�ʗCx��V�4a�&M�]�[��0mJ���( ќE�e"D�}m��ϓ�|�s��p9��]R�^�@�ۖ��eo^��J���b�I����%yh�N	��+�-+��'A������2'��#�K}�-�T�@���8jϔ��1�n. ���v�����d�엩w䵜B�6�����7��I��<z�:kQ��gF�A���ب.��h����h� ��V�������̩�q	�0ԛ66�s�ny3�ﳰ��]7�>�7;1M�)��o�C/���Q1ꧩZ�q�mn��?pQ� yK8[�j>���kݦ��UN�J)L^���i~RS��i����ן�D�L��y�cL�$�É"o� �Lg1�Bx(��19a�G�d�	p-��O%�c���2Sۦ,L��gu����9Z�׵p�Q�"�2��8,���\�Y�`���N�ڟDd�8�_3S�z2���I���%O�]ph#��!��m�5���\�i**?	+��q������� ���g�%���Ԗ[�1��9��9���j&G?Y]�
�'���*�m�'Uo.�'���b�j�V��C||�S�#N��~�w�r�ZH�M3��͡���v�r����
ʯ����!�@q� %�AL$�^�A�vO��;0j�qN��E�.���:���Ԋ,o��E��o�C%��ǲ|TX�3J�U;���߽̾�E�"�F�(�#�]��*y�kYY\[bm��u��G�"�khG�W{�ʂ��?�J
pf��>
G;���ӄx~��OK�K��8`��b<و�?-ֵ�~F���]�#�tpTP7z0�9eu+��^�E2�6�����1�	�4��Qŭ��dN����ZU�@��>�k����$D�n�<�� �<�#�|�?V��K�;&h(b���@���q�����~"��J	fC��̈́���%k�^����Uo�'�A8c��!��WM����o��kf8��������DȾ��F�����CkU�6��X	wa���%(�g������׶9в.W�w73�V�j�n�"���;ǽ�"k谷N�\��s[�w;�:8��D`Úk{���kw��Kn1s�2F�3 ��V�����/�e^f1�!ܣ��mW�Ԩ��@���zO:��]+#p�v��JO�T36���t±/m�PIn��I���8�4�E�Byr���@�M"�)~��ne���fSH�K�Y�M����#	IB���� �U��K���AW���� ���ޕ�DkB��.��杻O��T�B��C6y�s�����%J���j��lcz^���6�s�>�z�#��0�=Q�f�ƫ��-؞EoD�=�]IA��lɆ�_3l�Gs9'�I7E��(h ��d�mwl��$����1���)��5p��ZO�r4��w�B���E�i-Wr�P%	e> � ��������Q�.I�WC�k��˿��v���;S�A��wǰ�1�n:?�7�Y!n��iT��&9�huƳ���W��L@֢��9M�卵��)�����'�޹�� �߳��b�he��/w�� 
t������'JZZT�J��d��F~�Y���4�b��2:TI�娘���l\Pc	륟�*�l���-P�q4��'
�����]����d�����L��������.�f��U�ldmFz�R��+M�p��@�m�;\=9��x���4�4	%����1��.�S,|j�8��X�N�����	{y�ޜc�R�S7�_#�N�]K��k���e�͈���W�����4�Q~���o��]"�2|zqo�y��يP���7`�[�)�j˾:�i�\z�v �� ��6;S���b��b�O��0�;f�(_��Tk}!�$O��+ҕ�s�����I��r�e�;��roR��̷��|�{7Ɨ�4",?>����m��ߕ���9��U�<Ɍ����hR�(�{��x��(��~M%n�B �:]�5]~�앁8���2+� ʹ#��_SB:[|UHo�c��:o�R���e���"�/^�X0�l3����#�˾��}Ѭ��k�����1$�U�E��B���Q<y)<{v5��, ݖ2	n�Y`(7��A'|聋^#V Sv���(���zb����_���0�h��E�c�EN'�W�>�$�����4_�@YE�n��6Caح�9�#iR�
0�~�D�^8��ŀ(��dmLB��f�rz�u�]�D�ꎟ�BWT����kv�7��b�t�}�iK����!ѿ�����F<t#Y)���B~>k��ۨ��L�����'*�6��luL&<x,k�X ��UY�N�?�c@\��T������ið}�VΨ�ٙ�Y�6X���.��/ƌ����;�:>�Ld�h$�j��Xz�x�1_;*�k��5�/�B߸�>r)ؘ�r8LA�˱�<;Lv��~g��������'Y6�=������1v�����LfR�2��s˻�g��T@p��a��	�M���zB=����cXY,K_�F�������O<r��0�V����)����/��q��	~em���A�Q-�?��Si{�PRj��k��	;�����i,�)U����JG�Ќt�!���H��@��h��z����4���N���t��y
R��_�,�Q.��;kpf.�)�,t�%}h~��?rm�sE�B-���`��K����-p�����R!��EhfNU��nǀ.��cR�ln�����0��bᴷ~�\����!'�����%c�TP$��ot[�8�E%U5�ӧ��0�0�aw�C@�եHї�+�kʹ�l�\�~����3䕶Qmҧ�
���b����񸰐L�Z��*�p�6�~k��s�-�Fn�����9=��|����Dz�b0;ޯ�&o[iR�p����WP��e(���@���^�=��_9X�T��Q.���TP�MJ�tqp6���ߓ��O��m �~hhvɼm��Ri�lQ̀��`ԣ T�O�ǹ�r�*����o�p��Y�O�g��S�O����i@z�:�*U,He�`u���^R�5�%&��4�m������]��=����j����+H#2���W�V0�Vt�����t;��NsS��)�IX[�|�%N��MfSϓ����K��E�Ք�-�ǃ��|��N��cn��0��C$����7j�K=���r�6��>���PٛaH������f�N�-e�w
�A�G*1{"��Zj��(ȼ�k�]���a[YN��\![�ak��F���٦��f|I�Mi��S�NZ���5*H�4���N��(����i'��LQ�՗�&�@/�����䞳���{�5�\���}2�$�r�� ���f��U��ѧ��W��'��i� �A�Ad��_z��� a��,e$m{���5Ǐ�b��2Vdk��������0��g>?x?NP���*����������'`�r��o��(�,X�i����jn>G�a�t˯��� @� 
!�&^R;z1�{Ètڲ�}�	��Y-��{O���b�Ή����?��m�ob�׍��ӡ�H<�XSЧ�7a�W~g����l�t��O��H�F��j�H���@~.ކL�0_�#�m�9�ܴ� �.�9T~�	X�MbQ�lJ����_��[�n7	��e�v.Y�yqMJŝ7����w�+�nb���{4�z��q*r"���1-���e��CAQT���Jy<����%�Q�H�ߡ�R��h��5�4��=���{�y�։���X�^��	� 0��U[���Ԩ=Mo2���[�(ۉ�Zh)�c�����>kг��q#��5�{�m��zW0�{�����)�u�cМ=���i�f��2�<4o����p�6;z�"``No�o_���[Z�Y�O
�f�T��� t��n�/��B ���<t<�-�����K�׿�M#���� 浜�|YC_gv�1�px�q��K��iIKe�̉i�N�-.�/ߊ04��	�1���ϡ77��V�rv�������_)�`9�sDk����}Ӻ/h��d���$�N���1�~v��^"�MS�K�	C�Fh<�����ԨO��|��vU�j��"K�L��ed� 'ʘPu	��p�z![��gP��i��=��r&"����x٥�Q����]�xtc�R���+�K!/����(����A�5]W�Q���L�G�'�j�!^�a�3�a�
5���<F��yL1�Z�aÚ�0:�$x�Je�c��^��ڷ�nY@+��ۏC2-0���#8�(D��H2H��>�{���:�X��<m&^ͬ��т{��<�(�$���	5��|���_�%FS������yߓ���j��niC���:�w1`�0��5cHd�\�2v�)�L�;[B@�G�A�m�Q+�ه2�T�[�MZ��*��y:'��g��>-flD7�UVj�ژ0�<�����e\%�)C�uϊn(0����M#b�>۸�K6�1�&I��Pƾ�wi!�|�m�O��0�N���5muTY��=�3ba�)GƐ�c��k(r�q��!�r�2=<� }�����ޒQ}�J\��:Ϳ�ߤ�z���^�t������6�'�,�t��� �j	R�����5B����Ʈ�]�pԁ���� {kEF2�����Cԃ�����B뎂��~V�[)��?�x-3-5�d(�4��L}�~���������!D6>Y�5�g�Jz��t-�u�m��ᰐ�[7a�� �ǲ��P��H�6�Cac.n|�%����+	fx��jn;(��\VD��"�0i�*����Jb~x�ޙ�]�t�	P�N�m�4C0��za
	6s��i�&����)����g�
����ueGB�j�a}Y3���40D�M�p&��U욝4Ci< �;=�W��HsS���
#Oɦ	�:�Z��P�� ��aņ@J�'�M�?d��#f�P�/be�pzgp;h�6uR�Zo?�<_k�0�PT�F�1j�V��x�Q����)�#�6�v3d�>_��UlXo���#g��%�p2[z�o�����c �G{G��wt���2��-w�W�#c0u�$Å���g1��I�%k������F����9�����N���qh;V���à���tjS���q��ou�3���0m�{=��_az�5U�vD���[�&C묗�@��dUv�No1����|<H�$cg��
��qdk� ����������hU�t1����3n� X~��������h���0qfC�>�*� �����:���8��]xѝ)Q��7Eދ�pN`q��`�܊�Y�2y\4HyxK��)pn.�`�ό6v�#M�)�J.l�%c}�>B���4� �O+�N�ȝ׭u=��3�dǗ$C�����:��s]�����%�r���j��b�����Q�bb������A0��GR�������Y�*2�T�$a�������|Vt�t�MQ��y�zA��w�@q�z��)���]����{��Y�%+
���<HƎQ&̯�җ����5���5�<�]��7���<��)Yo�{``/t���"�b�FAh������3� �=䮃�Fld��u0��"
c���ds���_^�A��;�ωT����RA<j����z�^���X�Lu%b�ͳ\�GÁ�����
e�x� O-�q�-�E��H5E��p�ù��L��,F���x��eA�4�Y� a����ȥ]����܁ڝ��U�24�֝׃p��M���������(pO�LFe%�I��4`|��U_����SMY1����U��tK^�����_/���C���S�OY_�sy�(,vىOXs���z��pȸ��̠c;D/g�YR����'�I�9At��,�k�� !��O�D'�cIgϤR}%s�f�:s� ���d�Co�Zj���o�M��:�q %Uȭ��u�RΤ�h�>���;b�⯣M�v�l��4��Şy	ܕ%�[l�Gs�t���^X���g��} !(�6��<p��y �����������1�vYG�t�v�_�,[�zZm&Sd}�ڋʭ��� dn8@0�U%*7ۆ�nNڊ'���|̦�ᆍ���-��[+�C��~�E�;�H�l�N��HU@��Q�q���B,?J�l�^	U��m�������#<��A�sxC*���x:v��eT�Z{dDV���B$Բ��~'��fn$�E�w�S(�5�8�k�_�&�� �7cxJ-_�<��Tf��0�����(A�!!NC5�E�B�q���Gꅷ�ל��`�e\���Ƈ[�S[��fWp���2+��kv)�"���G��P|�m��yO�����ϙ}�J��
3�����r�Ϡ����<9�@��b����p���	t^�ʩ�����O�Q��j1���ͷ&VǶ���J~����KH ����黎�;q��-O�/Ω��jEu�4�G�5I^���o(�����U�w�x��!���_���M�9�)��?�5d>��i�LxMϚ=�� G^�i��
7Vx5�WA�_8HB�>������;�+Ћ�m�e���M���eD��/��"�g�}JR�����=%�Z ���n1LR��`��/SVR����#>�H���	�b3B�]׈�<n�B��s"�ckl�F�+��	-�oa��׍�:q��'��dw&���������\�� ��X��M�5���ђΖ���.��ݻ�yr�;PL��)C9�<6�w���(�/
�Cz�	�'�P�I�+t��ںI�L���Z����%��Yp:�3�s�K�9.�� �U���T+��;��5oPO���·�
�QU��h��$Rn��������*����T����Y��sW��s��k'ĸ/����Rt�h:x���W��_��<	���<�A��=��c	��	��E��y}�h@� 叼�x��G}��f�"nF/{Jn�+��6�Y7��$}B�C���,6��'�;��Ӗu��Y�ܠ��Jxs�AT��P�A�)_� �Z�U>N�v����?�cﱆʆ����IoT2���J���|��p��ü?a�C�;�_xJb*�}�EB��	�o�}�{�,�G2��/f�D5.�5֯�Ի�W�O�b3}�/��)�U��ja�X�좙iZ�E�u4��˘�OYW��f�c�Td�[�~z�����n��[dU�5Ӄ�&�NY��0��e�tbӱ,ˀ�Gn*�'�#���U�QݷNlk@SN-U'�����d��i惡SBA��K��"�j�~b�E���+�i�٭bP7�2�h��g�U����~!Œ���]��cZ���dI�Xn��� ����0��2� �.� hr��a/-9�a �G6�xX)9=wK���[	q��Ow�zo���;�U��tT32V�{�-F��O*��bAr��}�ň�~��+��K��wB<R��5P�9�>mpإl�}��8~/쐠w���@Z�v��\��P�r m����X6�@,��8s�e|Iv��k|����tP��J���p��%sֱa�yhZ��ց��1'�u�N��0�S1��v�����h�wN��~��������|2�sjVᠼ���a�k�)����,\՝��
k_ ޵3G����l�U�j�W?�X�~�pnt]���|WG��Z��	�}e\��ӎY�����Sj���{M���`f��b�4J�{5z�aM��\pA�?$r>��<^������Z�K-�Q?`P-"u~�}rRMe���� ��j�rR�`E�L9@A���J9Scy��=���S�6�3;�.�����\x>ˣ�nO	X}�	�ŷo>�ԋ�8�,)B	/d���h��W"�lV�G�/]t\����oR��T�THi�'�	z���aa�$��n����p{��2yƦ	��;�p��ɶ4>�6&�.Tw�*G5��VFE�B�j���R���t�(xi�x����2�3�X:� R5��
;6l]_@r.�L�bv՗��0�3C���>�o��/c�]΄����k��!� �`����U��e��r�
���>Ґ�	ߌ��"~fe����`ʖKmզh�<���|y�ز�=	��?���>ھ����� ݢ��x
��MϦ�\r�ջ����zr�P2�к�������u��j�n*��Z����񫁆���
��S�����y)�S���!���vW�8;�4umt�$:���
q������g�cV*�s�te�G
���{�� ��kOQv,��5/N���=�
�}"_ę�Ӗ3w�2�:_��o���x�P��XSz��>*�K�ض��Fu�ݥ�vE��{����B:��w4E�+79E����~2��zm;Xy�r�82o�"�ܐM��j�{Zà���Q��v��f�iձ.=��ݪ�d�K��3�zuIW-Dd�����8K�6��JA�����%r��_@�R#F���?�-���-P�0�I�m[a-(��b# �}�ź�C&��(�r;�W�������ª��qz�w��QMb~��<i�nN�cHU��W'�J���m
�u�������];�G��Q��/Xd�e���Q���a�E��&��Ě���c#���KEOe*�h�dNsP]�^Z�����2�cv�P1Qv�j�>R��ԜڔW/Ke^K\��"v1��L�R�T���,d�{�9�x�/h�p(�B'@��&%W����@nMy��֛��%��D:���p� h���dT�1�p�Wm��lpl���sJ�eP���Z�����ok���[i�?�SH�P�K.�m�/�^e�ɾGb��t�b� |��ϋo{�ےhob�_|dQp�����)M�GNbV�58�	�z�������+�#��;���wl-�>�K�H��gy�����*�+��x�S������3��q Q�Ŧ��9M\�:j�m�k�%�M(C���%�1j�'%ނ|��KH�P��yoS�%�nh	Xy�r�y�H�j��t\��{De�
F�/�ZЙ��ӏ�����]��p.3*�	��Jr��>��G�T���M���������a{�9�?`�A�p��1��
ҡ:�`�Zk��.h�i�b�;�Pz��F:�,[�'�HG�j�ƽ��w�J�}�Ź��a}�~�5�U��X��!��Ê?K
�S�'P��];��	%Wuf�)9��0l��K��}��y�|V聎z̎d2\qq��ó�{"6����yT� �^f�Msx�3я��rwK�q�]YF�b��VM�8�*8�2\�����~Ű��OJ� � �s�L�< �:6�~O�����+�������I����@�m��5�9ǅ��D���*P(嚽J�e�9��"#*�}��"�[G���;+JRX����w�^��Y�R�$�8���f���J������f����`�K�J	r�ފ���'^O[]���VF��	Э���u�T=PlV���8zH�������8��ͽ�2�uzL��Wk��#��^t�.�yV2%�i3`�"��	Z����+�)���h��N)6�c�S5D0D��>�#p8�X�.KAHv�ɯ�`ߪ}̮���Ѿx����*�Ŝ;ȍ
��(@25���Ѝ�O��a�v^o]��]����G�M��!M�8�۷($?1\��kҡ2�v��W3��W�NnY�b
J���s�\io�q��ZY��<�E�}^"�P69g��(>���O�Ɇ��L����%_���M<�A^li���r��6y��0]�����?r;�&���3�g��l_{H�n�8Q}�fʏx�*RZ��I��f�P�`%����m�!Qk�zA�E����D�P�1%ƶ���d�nG�s$�r'1i\@��+�Z%P��i�5��o�pp�B����S�&[g\����L4.3''vqN�?�ܷ��j.- 
o��p�.u+�\n��nk����v����b�*�E�8��0N��5N���/��Vu��QUrў6\G����um��;�"��M��V
Id�◹ޟ) o��{1\޽Ɠx]��1p������$��d��>���w���x�����v��ܑ�P�G���L��^ɬ[��D�]�P��XE|�V�5���vdhr�_g~���#H�c�^7=������D�t���ӖM�0�6�H!��>�aIM�J��ńA�c;Qۣ��v0d��u"���v�o5uFz��쥼Ա�/���ݍ���e��v;�^����x����E�*%�=���j���;�wo�)�{�n?"��辰�[��1���Goc7x� ߫|�K��粽��ف���u�K���B!��y*�`��}K���R�� l�7���..V%$ڨ�"��N�j�y�Z4�b��5��t���`[�~�"xfmu�(Fl�B�������k��.O����,�x�cHv�����a�s�����ğp��� J��)HA���ϦV�]�a�p��ҺN��i�6�OC���LU	�hm�mQ�uS)�r�����%3��������������Fv���-A��^]����{�J�T��A3�I��C��	[�b<9c�.0�$�	���U�fݎ{�Vk �
<4�m�SHn�!ks�
O�	W-�3�T�q�j�oS���)��0t|���fF�=���܉!xa�oS��pNq�'�C��YL$�[�E��oz�2$��6,۩�	qi$�,7���b]:^C�܂(\�<G�駐�Y(����`�π(C��,���0/6qcb�*������= u���9���_�P1�B?+Je�F,s1a3����l'bQ�3dܡ�7��9�c�\��Q����-���􀳂w��ۖ��@}r�J�e��O�M�&6��{<��Q>��b������.Z'�h�"r��L�Z����8�ө@�±������ˢQR79#q�xK��ƭ�L�.��j.��+{q��X9�s��sx�r����� \Kv�	�໚��֮ _Q3!9��}�}��'FXr��L���ɼp��Q	$/W�Nԧ�S��#G矿/��^���W���W�o�c���3i�bb�$U�lubEX�?J����r�^Ec��`ȯ�4��4��,k�2iw�#.����5`Uz�rS�ObΦ�A]\��xy\��7	-�Y[�A��nN!�'m?9��Ѧ�Y�iPAs�Z`����l>����km��'�O])��kk��K(��ұ�ĮܦM������ދ�6=^i-��&��º��G����q�C\���H�^�[��4m�-���&�b�������Grg��QҺE��4 Ծ�ȇ�ƀ�c��t�w��Bg����vD��[ G>Yᙃ���e	�ۢĖ�B�|u���6���5#M��`���53�=�b�s����H�J48(j�?WH�"��z�Odݫc�4SR�ȏ%�2��M]t����sNq��9�#����=>�r��4[�O~l��Q:˝�����"�yO;z��솠�/��N!V2�C��@�G�q�F���X�C�����
�O���z�&�.!ش�e � �P�f-R� 6��X�+�[�/3{z�	-�R�B�?�˗4m��.(��
p�>�ɵ���3n=r�rhhr��]:A�A��2hxn��w�0�'h�*�w�b��hfMQ�$�^���%��ט�BX�o��Ȳ��D�~&B����xw$�X���t�xu�'��k�b��;=��L�F����K��-�:�R�G�w�	k��Ё"��i�~���!�{Ҩ��Ȼ0�w���S�M��3BH���#�nv����F�C�� "Z#�W�Gs�L���YM�X�Ә�؂�TѺ���{�_tN>i
��3��-f����W���X��߬��XCR g���x2N�+�ⴙPt�ԍ��	�6�OG�`�+�H����b��{�Z�ה���m	��Z�=ח��[]��+��ϳ=8��z�Ԫ�E �Z!75�v��?���K|��]��ѻA�9L�t�z��e����S-"h��@@�;jh����|٢A�`K0��G�U!���_fĐL�ۺ��&�j�X.3Il�kPm@H/�l�r���G�b&IF�1�RYPd'�D)L���>�۲2�]���ϵ�}:h���ƕ�Ѫ6Y���N�n�:w�4���'BR�|����o��M �A�_�S ��.c�-�Q�H΂�
Z���Y���� H&	k\E}Z��/
gM^x�*��K�.S}��CBE�i�e|:��"✐"	g�fg"��B飨�s�d%y};��0Z�y��o�S6��Z�xߖ�M��(�.�T�$�}�=J��R���b&�U�9���`c��ڧ��Ȕ�%�sg�:���s7�i�����ݦ�/��U��hY��濫N� $3Pz��nDSYHf��!x5��thi�(��W��~�fB�
iEja�#]k�P�<e��D!��h��wN+V�K��J|�۫��j����L�Q�[WCq�MHi�;�����MQ= ц��I v&.����Ĥ�J�~����}ʇ
1O��
��)Z�t����I�R�U.�T �]�}߉��,����O�%tr��kc(Yz&P�ͧq�L���[\�}P��k�Y�
+�P#�P�d-�0�>��`�#���3E^�8��ɍ-�����d���\,���(2y���	�o&�%�qB�: ���8-�����9�BLk�ڡ��|�����f9����E=L���A�����4��%x�P
���/��e�+@ڙ�t� p���dsBo�[����T*%��F<̨�����RgK4f2/ ��?O��z��u#�XA�K��|͎>e�0@�h4�:+;.(��+F=CaT���Z��%%��n9q6��톆z��ǒs��v����.��,����˴û8����>�Ŭ�iGL�Wj�Ț�ۂ-����A��1yt���~RJ�� ��_t���A��ɇoÑ�a�%�!+^|V`I�g���>�g� %�..�Q�Y�^}̏�BnXL���`6@�0yt�Z��n	Q9��ŅH-ɣWKG疌p�Z�1�~�"w ,��,EJ��-߯�ּ4ͯ�b��|������t�鉛���֦�m��u1��c�}��ocV�^���'ߤ}|���s�jt	�<��kL&�z�����Ex�-c�o�P.��d�1S��U�>'��$΍QSm�'�iMp�����r�G�]�7�N4]��g��0YC*�����m鮍x� ��E���tس��x@�]#z����fD��~�+��c���Z:p���A�4�F)D13g����њ_�e=b�2\k�Ϛ�t�Z���FHM�P1ʪ��/��M�s���e�lTNU%8����LEV@FhIq�8hr�`�ި{�*�A��`���%�p�_�K��+�^�ͺ��
��wCۆ���*@N�ֳ���U��0][���F<ZSy���#�YV��݆(lKPE��N5��O烀\-�?�f�GŦ�6L�h�IȽ���o�֐��LJ�&6���PbզH�d%ڤ�=f�zR��)`=�+�iX9�Ro��$��� �f 	Jε}���n�����t�90p���i�@��
�+�̰N��gx�G��}����6 ��9h�lFA ��v�n�aΨ�R���fO#�͐lQ��am#>;.��z�Z^^o��xL��2�+-�*Эf%����-���NS���cƌa��ƪBa�.�p�ar�TGD�y�牭ϭ��+�����G��-�p(�VI�+��	�#���}��8�0o<n���U��m%{�J��j�P�,s���`HN�g�cz�V7^�N�������s0Pm�a����I�$b[�-[�0�_�ֻ�N��ژ<�$��ɹg8 =�0���Ӂ���VK7�9�.�·�F%�pC=]���<ז'B2�اQ�8�����TfM���4��H����tV��U��V��P9m,!Mq��<�,��j�y��m7��Ay��I?d@|)˟P�cYҞ��碻��T<V�hD�Q� �km�d�)Π��N�t�8�["�Y�"Ll��̠��g���e�@��|�-(q�
J�LwÖ�Y�&�4Rq@佼�����(pX���I�P�Zh
h١�0���-��}������t0�J���g#C�h��P����E:��l����Kv��Dg�j���EF�)�� ���"Q*�����$��-&��9���7�}��2�>2���X��7,�%D��k%E�~��b���`.�O���H���5�ml@���s����+y��܍�s�n+�q�jp����С�2�٠A%�� �$S�$�8^��;|��Y�9�n4�1�� ��Z�M����4�b[?�����1�5�&��&��k���c � z��m�4;%w*��"O��&�����l�m�Μ���������c/����̇O��6�م`��B�4�Ɗ�y���#EGq�9�~is$��"�;~˒���l�$�chj~�Ğ�&�S��5:\S�R��]g����ŀ��Z������҄��ՄAY�OT����ʜ���� �Z׋����QQ����{J��E��|mɄ�4��馳.ܶnv˟����V�����ѕ�ݐ?
m/�K��l�俤{rR5��%g��ʐ3�ɨ=�%�`P���-ﰧC#0�^$I� ���ʢ�Ț� �X|���`<����l�I�����Dmߞ����=�N�|7�7f�SW�dp3Ϻ���[-�E4O�9�(���\�JW��d7��d̝sV�%�ucS�R(W��^�W|"��U���`�Ur5�S湵�t�vx�͢G�-ȹḷ���s'[�;z�r?��Ñ/���%l��B!H�4G�dA蜗'?M�&�`04��I[�4�yD)t�z5��{�\��Es���E¹�7p[͙f,�z?Ţ�F^��.9�qQ�vE��܎?��g��s�6z�=X�dR�e��s^ewn��r�>fC��9n_�{Y�T������\R��P�d heM��Yi����g�7���F����|��A7�J�q����;��fW6j�;���"���l��#۠�!��Ө~g�?���ɪ��ܥ?1P6�Hd*�iѠ�eUr��8��ז�
	��K{�/����V$��&��2��{+?7p�?�.f��������h��%�)�㭈��o�&��~�2�1�q�v��f��cU	T�T�h��  ⚛�pq�d|^�N�����y���1�:������[��~�4��?��#�h{���T�S��^p,�*�p��>��IØ���BՒ��2�r������K�k��A@�N�A��3h�fX+���'0�ӏY�Q�q�k�@��?"�/�GDv�F�c�2	��U�a�A���|�1l�65v�^F\�1�'��<c9���Oe��Ш��Fs�t�vλ�Iz��Й���G�Z��r̸�x�j�:������w:R^�%����7��ډ������<[7T��Cc�Ә�/r��c���w|�D�e��K:|���`O#/�[���f���Q AM�1�8��������Ź"�,JJ�z!���q����v��ݲ�����A,2�t$�H<��e�Ά�i�іX��+��T��U���^hWPb� ,����\!��ގ�rvk���GF}��ZPcv���\s6i��Բ��l9��~��*K�l�̍�.�&���j}��9���X�L82�Q�T���ȋPT��:���خ�U��5���N|�9�lk�u?��r>�J��GN����{�A�Ы��+~.e^��V���p�����/,����8%�r�b��9�ZLO������oo+`�O���p��Ul? v��t� ���l����`�Y*�C9i*��.�I��0t� 4w�{�.��UE��{~E���O���`�іۃ:��i���e<��R���E���A�M'h@vF$)�x���[)��dM-Q�Z��<�Y8`B�JKf�k 9�#V}��V�L�:��V�v�\�2���2�RR�8������[xt'�͌,���b��5�9n{�%��&���me�@Ԩ�ߚ4��������M	�}l��������<y��Kj��Y�m���H�a�I\�x�ʆ ���G�, S����s��`�B\�6b���	�Pq���bM����'V�0�����'A�+��4�T`N��z �f�ԣe
�o�u_����-����� �'>	���)La6�%�[v�l�l��O��o�Y^�&=﹉K��, �sX��p}�l�f���'wmdчw���j��"��-����)z��f��%}F�EDe]a-{@��uI�d�UH�J����`�w�+f�����Ԅ�^�y
H��c�g<#�@�_�9ޮykNƘ��30��*\]C
���P���6E^�bU?��A��J�����Oe�8<`-�Ċ�V�h�j�l����Q��g�$B�e~x�*6��_��wirq����5K�S����[/i�rP�c��"�p94�#�`��
Ð"�H����L+U����U1���V��η^��=��c.�[A�N��2ƶ�����I�m�3:��Z^FU�����{Rs4.ۊk�D�h�+�}�),�\���i�e�O�����l�_;#�f��A7-���Ϧ*�|���s��p!�4�p�	�"�;�1S[0��_;QX���:-CE�G�p�����G�=������j���9�.l�mNZ3t�F�Y$�~�IP�t{=�AqG��2��(p���fB���"vͮJ��V��˙N�7�d�1+:��m�&g�#>��p)�:��M�1��,i[�jlU ǤEcyF��l27Ib����=��@l�Z��7�6.���2����ӿ�ɗ,�~�?_]?f8&�bؽ@�N��B0�q(\�	B������ߚ�\1k���m:�F�;��@�Y���!��T�&9����W	mb���!E��ǂ֔��;�,6K*N��%BLi��r7�X	��m7
ceɌHO�q;rt��엾U���r[�LP�19��i��o�%Q<�o�|�7-/��B����)T|�d�(i�"�� ,�y?�/�gvU*�F�dC���^���.��Q� �oX�2%���8��R�!.��^��g౼EJ�m��M���8�0J�T�`x�Bo� X�_4��0��Oa����������D�T$+wJ�n$��Ӝ���T*�-�%|��4^�a�|,q���9>�GOܖB���T^��Dt��bn��#��&m2�����Ӓ��Z h�Ȟ��.H�gta�i��_1-D`�0������F@��e�6)^O�W�l���wL6S�O����8�`)l���ϑjS@
������^���ݟc@�R����o������Z����"q&���R"'V-;kFQuq1����\�����HNwF2���|/Vu��7&<.J���_'��Z��V��״!�)�C�6�.�ҳ��H�����U�Bo��,����uJIbZ�ض+� �m�'��r&�����!d�s)�>�댋D4xd�h�fj�����CZ�x�*٫�^��}��T�{\v9C "���L�ؤ֩������	�Wy�#)�Li��)[����F��}��E��y�"�,~dI��u�;Nb�B(F�/�y�Z���
�������{o�{+�H�+N�Ю��T{7-���"8��O�]�Aq=�������5��w�r`��ţ�v'�*!���S����*YYi��f l�h�x����J`�e�e4�N����P�󛡚e^VD�|z��9yJ���x�DT�<^��bI�GJH����g��׳c]�q2�aT��9��~{����x��f�_)�ɬ�@we�t�6���ٗ���p���kQO��[�l�lVs�[J��M�U|Qﮃn�����͔f!��lY*��Mh��G&�!L5ƴ6�1�֡?�J1~ז�5���Bb?E�U��#c������t�?d �zFRf9�^&�dr#�Wc�����Er|�0{xg�^���&�����m��0��0l���jza����l8����=)B�Z*�W2#DN�z?�(��n����/wsp5N�"T�'��]E8�Q����,R�2�U��A;02P����c���zsP�������:�D����`ܪ��M���u2BD��N�;WbP��N�n2��Y�g�e���y/ʲ�.��~���}���
�>�5�L�e����3z���6=���n�nh6ȟc��gh���@��gLA�릇+���C�!5���Q�4�ߢq!}S�Қ.ڥ��?L�Rȿ�����r>j)3t(L��	��J��R��h�L���rp�~�˔t#�p�˕_��"��K6$�g�*�5���{I���(�ڸ������Zן�N��!���q\��/N�з�O�w�A�o���mb{�^ؒz��<XY��f�����v�7z�)��,U�	��;��?c��Y�!�%q���d�Pv�Gi;�1�YA�t�d*����p���_g)���f#��ԯZQ.��5䯴�%)r)��"l���G��?�(W���@�)�T��{;�W<k�CW����Ἐ3�B!C�
wo9�� �zkz��L3MiH�tJi$����º�5�\����ޮ�k7K3��ۗr 8�m�8x����?蜻}2E�졔��Hik���}1��{̷�Cu�vA2�#��jt6-�K��,ʓ�$ϡ�%���(3a���ME�/e�B��Ѷ��E�����{0S�>?�Xgd:b8K��3Z��]B���Խ��Zo2�Y{4�4�s%�O��24�<��tE?�H&+���ݜb���.�VBʍ{x��7o�d�[`��ia
'��9i�%�ʑܟ�Üz�K����W���!�P{<��A�:�g���.)���/ɿ��;76h2�r�o� !��w�R(GyQ\�T��b-�`H0t�
��2�J�g���|�V�jk0|%�".�V˱<��V���)��s�/��(���y�B8U��vM��Vw����N�?�����{=��H��2nS��C�MUڊa8/��5J(�9p���*�3;LϢ4 ��ȶY1O8�&ǖN�X�~�*+Ҷ�\
t�.������n���趹�y�u"�[zIҲ~��L�|㮉�����K^��/4��,k�e�{&}��a�)pWPл�ķ�=���eU��&%�!��4^�ݎ��8}(Ї����=��M���f�}���ǩC������_���%��`|*���7��)�Oja]��p8k��D^��SAUV:Qfm!�S�A{D!W�C3*m���Z�sп�2�X'K��~j��,w"z;�F�v��2{B�l���3[������ˆBP��^AS�Z�ŀ�4%�vk�z���l��u
D�Ǌ�'��΀^*?���%jr���*�Y��"�Im[p����8t���#�s�6��^N��ŏ!{@�&��&9�M�-ǹ����g�	�M�S���ſ��J�ɵ#�g4\_��;�#�j�� �7�<�hvlq�pE�L"�"��>�p;� �6�M�&��A�.��^;�Yg�a˫�n����z��	u�$�Ԋ��;������r��B.��i[U#�A/��t����ԉ���w2�鐻���Ć�0�@��
v�	��I]ۃv@XGϋ3��=B]`�x'���$	H�D��z�E�����#qu�j~���]U-�؉��CC�j��`.f�䑔�~�Ӌ�y�ȼ�ws�[7��r�����Aw�d\��E�Է�,����Uk}�����Z�Ow�i�t�,�%F4��+#& ���6H�4ɸ�d���U���\T8U.%�=�B����y⠣\�&�� ^ϼ��I-WA<sF��%hF��݂EeZN��u�i�A��e����}.��ṗ��R����%��If����(����U����}�;�$�7(t��^���^(ŋFܑ���>���a�����h�!�RZAs]����&:�U+��Mx��S ў��]`Q���|Y�?�Vܭ��۳gK:Ϗ��٦�3��YL䄜��ߨ��:%B�W�S��G�Q��:�{��.�ZnZ'�Fi+�� ��|�mBpX��/�@���51^w|��5�V�wN*�"'DRф`V��ە����7�'x�I_�)�����-���H|���wVkt�zdA+��TC�]�v�.���^C�)���M�z����K�ke�&�w6��hGf�$@./�a��{N�U��}^��m����{Z���*�^,�Y�y����Ʌ�ˈ�R��E:�� ƽ|�֢O����0ӄ���b����s��(���cW��ШuA�8�@b�F�IHRO+�����:Ϸ����T<��j$�寊�����m�PQ����!���� 9=W������P�>a��fX��w�CE���窲S�6i�#�*�$���5�|��G/u�kl�YY��z���/��H�'��|��ǌ~�����F��7.�> I�8l�@�YK����2�+:*J�!�M����y����e�y���w@X�H��P�V���k�r�.衼��	�j
#��:! �u�z���l�c�r��]��k��CYZ`�@���ί�	S�75D3F_��v�l��E�;>[��d%qMr@kggf+��������
�)_��T�����(��-uH�	.�UA�}�xH�c����V��-�C�L�Pٻ���y���P�@7~�MS�kP�������W��E�!&��
Eax��b,�e�hH�l�24<��}���U�+�y�TϿ#����q�T�_�:�W���iĕv�1[�T�BT��޻Zr)�ls���r������4�F��R�ա�%��х��Hrs����IrE e,i!S'f�V���s�4������ȓZ���Lc�ܵ!p `y��$��6p�;�m��"�x���^N9p�#�L�d�����X�-غ	myK+�ﺩ9�����s{c,LW�q���2P��u�#Q4H\��bqu8re�lA\x��:�y�D�vn��Z-��6��\X.#���>��0j��T�K稀$�S&ZC����m�������d���E��`��9e��J��u˕s���	 ����:J]wk�|���������;�m�T]Y��翮�o�f-��0�28p�v~����䘻M�׈�>�+��.��e��$�P�-\�b �H��򮿃�ө�&��&�-5���W+K zxх"{�a�0'"h�����Ƶ�z��������7$Z��̿lԊ�j�aL`���z�������B�E��i�*A���\pu5[|�����a�q~���<?4j3L��A>�z_8���ߠz���t��?�,�I� ū���\�B�2 z[9M{¾�(l�����G��z�B��f����!PQ#l�����/�4�I�t����أ�^�(�;x�fT ��7��$�;<[o�κx��!���Кo��`�Ï�F2���,��w:5�{r�H�o1R^����ROS�w����gh=h�v��5o�f?Ãx&��~AQgm'�2M�P����5՘Ȏ�U��G:f�|F�"N�a�������|�� ��WCu9mQ���&eRt��<B)�m �� U0?�5W����o�f����>�DP�yC�?� �8�PF����* G�M|�Z+j
K��G�-�1�q�@����=���yY�^˲�6�1��,v$�R���AE1�o&&�\ĭ�>*�Q�$��N��>����~�}���:F9ډ��Q��Q��+Qk��viP��ѣ���>~2���^����N��֔����2�h˱� ��s_m�