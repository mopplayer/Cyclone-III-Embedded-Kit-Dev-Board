//megafunction wizard: %Altera SOPC Builder%
//GENERATION: STANDARD
//VERSION: WM1.0


//Legal Notice: (C)2011 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module button_pio_s1_arbitrator (
                                  // inputs:
                                   button_pio_s1_irq,
                                   button_pio_s1_readdata,
                                   clk,
                                   reset_n,
                                   slow_peripheral_bridge_m1_address_to_slave,
                                   slow_peripheral_bridge_m1_latency_counter,
                                   slow_peripheral_bridge_m1_nativeaddress,
                                   slow_peripheral_bridge_m1_read,
                                   slow_peripheral_bridge_m1_write,
                                   slow_peripheral_bridge_m1_writedata,

                                  // outputs:
                                   button_pio_s1_address,
                                   button_pio_s1_chipselect,
                                   button_pio_s1_irq_from_sa,
                                   button_pio_s1_readdata_from_sa,
                                   button_pio_s1_reset_n,
                                   button_pio_s1_write_n,
                                   button_pio_s1_writedata,
                                   d1_button_pio_s1_end_xfer,
                                   slow_peripheral_bridge_m1_granted_button_pio_s1,
                                   slow_peripheral_bridge_m1_qualified_request_button_pio_s1,
                                   slow_peripheral_bridge_m1_read_data_valid_button_pio_s1,
                                   slow_peripheral_bridge_m1_requests_button_pio_s1
                                )
;

  output  [  1: 0] button_pio_s1_address;
  output           button_pio_s1_chipselect;
  output           button_pio_s1_irq_from_sa;
  output  [ 31: 0] button_pio_s1_readdata_from_sa;
  output           button_pio_s1_reset_n;
  output           button_pio_s1_write_n;
  output  [ 31: 0] button_pio_s1_writedata;
  output           d1_button_pio_s1_end_xfer;
  output           slow_peripheral_bridge_m1_granted_button_pio_s1;
  output           slow_peripheral_bridge_m1_qualified_request_button_pio_s1;
  output           slow_peripheral_bridge_m1_read_data_valid_button_pio_s1;
  output           slow_peripheral_bridge_m1_requests_button_pio_s1;
  input            button_pio_s1_irq;
  input   [ 31: 0] button_pio_s1_readdata;
  input            clk;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  input            slow_peripheral_bridge_m1_latency_counter;
  input   [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] slow_peripheral_bridge_m1_writedata;

  wire    [  1: 0] button_pio_s1_address;
  wire             button_pio_s1_allgrants;
  wire             button_pio_s1_allow_new_arb_cycle;
  wire             button_pio_s1_any_bursting_master_saved_grant;
  wire             button_pio_s1_any_continuerequest;
  wire             button_pio_s1_arb_counter_enable;
  reg              button_pio_s1_arb_share_counter;
  wire             button_pio_s1_arb_share_counter_next_value;
  wire             button_pio_s1_arb_share_set_values;
  wire             button_pio_s1_beginbursttransfer_internal;
  wire             button_pio_s1_begins_xfer;
  wire             button_pio_s1_chipselect;
  wire             button_pio_s1_end_xfer;
  wire             button_pio_s1_firsttransfer;
  wire             button_pio_s1_grant_vector;
  wire             button_pio_s1_in_a_read_cycle;
  wire             button_pio_s1_in_a_write_cycle;
  wire             button_pio_s1_irq_from_sa;
  wire             button_pio_s1_master_qreq_vector;
  wire             button_pio_s1_non_bursting_master_requests;
  wire    [ 31: 0] button_pio_s1_readdata_from_sa;
  reg              button_pio_s1_reg_firsttransfer;
  wire             button_pio_s1_reset_n;
  reg              button_pio_s1_slavearbiterlockenable;
  wire             button_pio_s1_slavearbiterlockenable2;
  wire             button_pio_s1_unreg_firsttransfer;
  wire             button_pio_s1_waits_for_read;
  wire             button_pio_s1_waits_for_write;
  wire             button_pio_s1_write_n;
  wire    [ 31: 0] button_pio_s1_writedata;
  reg              d1_button_pio_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_button_pio_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             slow_peripheral_bridge_m1_arbiterlock;
  wire             slow_peripheral_bridge_m1_arbiterlock2;
  wire             slow_peripheral_bridge_m1_continuerequest;
  wire             slow_peripheral_bridge_m1_granted_button_pio_s1;
  wire             slow_peripheral_bridge_m1_qualified_request_button_pio_s1;
  wire             slow_peripheral_bridge_m1_read_data_valid_button_pio_s1;
  wire             slow_peripheral_bridge_m1_requests_button_pio_s1;
  wire             slow_peripheral_bridge_m1_saved_grant_button_pio_s1;
  wire             wait_for_button_pio_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~button_pio_s1_end_xfer;
    end


  assign button_pio_s1_begins_xfer = ~d1_reasons_to_wait & ((slow_peripheral_bridge_m1_qualified_request_button_pio_s1));
  //assign button_pio_s1_readdata_from_sa = button_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign button_pio_s1_readdata_from_sa = button_pio_s1_readdata;

  assign slow_peripheral_bridge_m1_requests_button_pio_s1 = ({slow_peripheral_bridge_m1_address_to_slave[7 : 4] , 4'b0} == 8'hc0) & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write);
  //button_pio_s1_arb_share_counter set values, which is an e_mux
  assign button_pio_s1_arb_share_set_values = 1;

  //button_pio_s1_non_bursting_master_requests mux, which is an e_mux
  assign button_pio_s1_non_bursting_master_requests = slow_peripheral_bridge_m1_requests_button_pio_s1;

  //button_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign button_pio_s1_any_bursting_master_saved_grant = 0;

  //button_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign button_pio_s1_arb_share_counter_next_value = button_pio_s1_firsttransfer ? (button_pio_s1_arb_share_set_values - 1) : |button_pio_s1_arb_share_counter ? (button_pio_s1_arb_share_counter - 1) : 0;

  //button_pio_s1_allgrants all slave grants, which is an e_mux
  assign button_pio_s1_allgrants = |button_pio_s1_grant_vector;

  //button_pio_s1_end_xfer assignment, which is an e_assign
  assign button_pio_s1_end_xfer = ~(button_pio_s1_waits_for_read | button_pio_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_button_pio_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_button_pio_s1 = button_pio_s1_end_xfer & (~button_pio_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //button_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign button_pio_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_button_pio_s1 & button_pio_s1_allgrants) | (end_xfer_arb_share_counter_term_button_pio_s1 & ~button_pio_s1_non_bursting_master_requests);

  //button_pio_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          button_pio_s1_arb_share_counter <= 0;
      else if (button_pio_s1_arb_counter_enable)
          button_pio_s1_arb_share_counter <= button_pio_s1_arb_share_counter_next_value;
    end


  //button_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          button_pio_s1_slavearbiterlockenable <= 0;
      else if ((|button_pio_s1_master_qreq_vector & end_xfer_arb_share_counter_term_button_pio_s1) | (end_xfer_arb_share_counter_term_button_pio_s1 & ~button_pio_s1_non_bursting_master_requests))
          button_pio_s1_slavearbiterlockenable <= |button_pio_s1_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge/m1 button_pio/s1 arbiterlock, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock = button_pio_s1_slavearbiterlockenable & slow_peripheral_bridge_m1_continuerequest;

  //button_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign button_pio_s1_slavearbiterlockenable2 = |button_pio_s1_arb_share_counter_next_value;

  //slow_peripheral_bridge/m1 button_pio/s1 arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock2 = button_pio_s1_slavearbiterlockenable2 & slow_peripheral_bridge_m1_continuerequest;

  //button_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign button_pio_s1_any_continuerequest = 1;

  //slow_peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  assign slow_peripheral_bridge_m1_continuerequest = 1;

  assign slow_peripheral_bridge_m1_qualified_request_button_pio_s1 = slow_peripheral_bridge_m1_requests_button_pio_s1 & ~((slow_peripheral_bridge_m1_read & ((slow_peripheral_bridge_m1_latency_counter != 0))));
  //local readdatavalid slow_peripheral_bridge_m1_read_data_valid_button_pio_s1, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_button_pio_s1 = slow_peripheral_bridge_m1_granted_button_pio_s1 & slow_peripheral_bridge_m1_read & ~button_pio_s1_waits_for_read;

  //button_pio_s1_writedata mux, which is an e_mux
  assign button_pio_s1_writedata = slow_peripheral_bridge_m1_writedata;

  //master is always granted when requested
  assign slow_peripheral_bridge_m1_granted_button_pio_s1 = slow_peripheral_bridge_m1_qualified_request_button_pio_s1;

  //slow_peripheral_bridge/m1 saved-grant button_pio/s1, which is an e_assign
  assign slow_peripheral_bridge_m1_saved_grant_button_pio_s1 = slow_peripheral_bridge_m1_requests_button_pio_s1;

  //allow new arb cycle for button_pio/s1, which is an e_assign
  assign button_pio_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign button_pio_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign button_pio_s1_master_qreq_vector = 1;

  //button_pio_s1_reset_n assignment, which is an e_assign
  assign button_pio_s1_reset_n = reset_n;

  assign button_pio_s1_chipselect = slow_peripheral_bridge_m1_granted_button_pio_s1;
  //button_pio_s1_firsttransfer first transaction, which is an e_assign
  assign button_pio_s1_firsttransfer = button_pio_s1_begins_xfer ? button_pio_s1_unreg_firsttransfer : button_pio_s1_reg_firsttransfer;

  //button_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign button_pio_s1_unreg_firsttransfer = ~(button_pio_s1_slavearbiterlockenable & button_pio_s1_any_continuerequest);

  //button_pio_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          button_pio_s1_reg_firsttransfer <= 1'b1;
      else if (button_pio_s1_begins_xfer)
          button_pio_s1_reg_firsttransfer <= button_pio_s1_unreg_firsttransfer;
    end


  //button_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign button_pio_s1_beginbursttransfer_internal = button_pio_s1_begins_xfer;

  //~button_pio_s1_write_n assignment, which is an e_mux
  assign button_pio_s1_write_n = ~(slow_peripheral_bridge_m1_granted_button_pio_s1 & slow_peripheral_bridge_m1_write);

  //button_pio_s1_address mux, which is an e_mux
  assign button_pio_s1_address = slow_peripheral_bridge_m1_nativeaddress;

  //d1_button_pio_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_button_pio_s1_end_xfer <= 1;
      else 
        d1_button_pio_s1_end_xfer <= button_pio_s1_end_xfer;
    end


  //button_pio_s1_waits_for_read in a cycle, which is an e_mux
  assign button_pio_s1_waits_for_read = button_pio_s1_in_a_read_cycle & button_pio_s1_begins_xfer;

  //button_pio_s1_in_a_read_cycle assignment, which is an e_assign
  assign button_pio_s1_in_a_read_cycle = slow_peripheral_bridge_m1_granted_button_pio_s1 & slow_peripheral_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = button_pio_s1_in_a_read_cycle;

  //button_pio_s1_waits_for_write in a cycle, which is an e_mux
  assign button_pio_s1_waits_for_write = button_pio_s1_in_a_write_cycle & 0;

  //button_pio_s1_in_a_write_cycle assignment, which is an e_assign
  assign button_pio_s1_in_a_write_cycle = slow_peripheral_bridge_m1_granted_button_pio_s1 & slow_peripheral_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = button_pio_s1_in_a_write_cycle;

  assign wait_for_button_pio_s1_counter = 0;
  //assign button_pio_s1_irq_from_sa = button_pio_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign button_pio_s1_irq_from_sa = button_pio_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //button_pio/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_jtag_debug_module_arbitrator (
                                          // inputs:
                                           clk,
                                           cpu_data_master_address_to_slave,
                                           cpu_data_master_byteenable,
                                           cpu_data_master_debugaccess,
                                           cpu_data_master_latency_counter,
                                           cpu_data_master_read,
                                           cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                           cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                           cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register,
                                           cpu_data_master_write,
                                           cpu_data_master_writedata,
                                           cpu_instruction_master_address_to_slave,
                                           cpu_instruction_master_latency_counter,
                                           cpu_instruction_master_read,
                                           cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                           cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                           cpu_jtag_debug_module_readdata,
                                           cpu_jtag_debug_module_resetrequest,
                                           reset_n,

                                          // outputs:
                                           cpu_data_master_granted_cpu_jtag_debug_module,
                                           cpu_data_master_qualified_request_cpu_jtag_debug_module,
                                           cpu_data_master_read_data_valid_cpu_jtag_debug_module,
                                           cpu_data_master_requests_cpu_jtag_debug_module,
                                           cpu_instruction_master_granted_cpu_jtag_debug_module,
                                           cpu_instruction_master_qualified_request_cpu_jtag_debug_module,
                                           cpu_instruction_master_read_data_valid_cpu_jtag_debug_module,
                                           cpu_instruction_master_requests_cpu_jtag_debug_module,
                                           cpu_jtag_debug_module_address,
                                           cpu_jtag_debug_module_begintransfer,
                                           cpu_jtag_debug_module_byteenable,
                                           cpu_jtag_debug_module_chipselect,
                                           cpu_jtag_debug_module_debugaccess,
                                           cpu_jtag_debug_module_readdata_from_sa,
                                           cpu_jtag_debug_module_reset_n,
                                           cpu_jtag_debug_module_resetrequest_from_sa,
                                           cpu_jtag_debug_module_write,
                                           cpu_jtag_debug_module_writedata,
                                           d1_cpu_jtag_debug_module_end_xfer
                                        )
;

  output           cpu_data_master_granted_cpu_jtag_debug_module;
  output           cpu_data_master_qualified_request_cpu_jtag_debug_module;
  output           cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  output           cpu_data_master_requests_cpu_jtag_debug_module;
  output           cpu_instruction_master_granted_cpu_jtag_debug_module;
  output           cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  output           cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  output           cpu_instruction_master_requests_cpu_jtag_debug_module;
  output  [  8: 0] cpu_jtag_debug_module_address;
  output           cpu_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_jtag_debug_module_byteenable;
  output           cpu_jtag_debug_module_chipselect;
  output           cpu_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  output           cpu_jtag_debug_module_reset_n;
  output           cpu_jtag_debug_module_resetrequest_from_sa;
  output           cpu_jtag_debug_module_write;
  output  [ 31: 0] cpu_jtag_debug_module_writedata;
  output           d1_cpu_jtag_debug_module_end_xfer;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 28: 0] cpu_instruction_master_address_to_slave;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input   [ 31: 0] cpu_jtag_debug_module_readdata;
  input            cpu_jtag_debug_module_resetrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_cpu_jtag_debug_module;
  wire             cpu_data_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_data_master_requests_cpu_jtag_debug_module;
  wire             cpu_data_master_saved_grant_cpu_jtag_debug_module;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_cpu_jtag_debug_module;
  wire             cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_instruction_master_requests_cpu_jtag_debug_module;
  wire             cpu_instruction_master_saved_grant_cpu_jtag_debug_module;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_allgrants;
  wire             cpu_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_jtag_debug_module_arb_addend;
  wire             cpu_jtag_debug_module_arb_counter_enable;
  reg              cpu_jtag_debug_module_arb_share_counter;
  wire             cpu_jtag_debug_module_arb_share_counter_next_value;
  wire             cpu_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_jtag_debug_module_arb_winner;
  wire             cpu_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_jtag_debug_module_begins_xfer;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_jtag_debug_module_debugaccess;
  wire             cpu_jtag_debug_module_end_xfer;
  wire             cpu_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_jtag_debug_module_grant_vector;
  wire             cpu_jtag_debug_module_in_a_read_cycle;
  wire             cpu_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_jtag_debug_module_master_qreq_vector;
  wire             cpu_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  reg              cpu_jtag_debug_module_reg_firsttransfer;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_jtag_debug_module_waits_for_read;
  wire             cpu_jtag_debug_module_waits_for_write;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  reg              d1_cpu_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module;
  reg              last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module;
  wire    [ 28: 0] shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master;
  wire    [ 28: 0] shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master;
  wire             wait_for_cpu_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_jtag_debug_module_end_xfer;
    end


  assign cpu_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_cpu_jtag_debug_module | cpu_instruction_master_qualified_request_cpu_jtag_debug_module));
  //assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata;

  assign cpu_data_master_requests_cpu_jtag_debug_module = ({cpu_data_master_address_to_slave[28 : 11] , 11'b0} == 29'h1001800) & (cpu_data_master_read | cpu_data_master_write);
  //cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_jtag_debug_module_arb_share_set_values = 1;

  //cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_jtag_debug_module_non_bursting_master_requests = cpu_data_master_requests_cpu_jtag_debug_module |
    cpu_instruction_master_requests_cpu_jtag_debug_module |
    cpu_data_master_requests_cpu_jtag_debug_module |
    cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_jtag_debug_module_arb_share_counter_next_value = cpu_jtag_debug_module_firsttransfer ? (cpu_jtag_debug_module_arb_share_set_values - 1) : |cpu_jtag_debug_module_arb_share_counter ? (cpu_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_jtag_debug_module_allgrants = (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector) |
    (|cpu_jtag_debug_module_grant_vector);

  //cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_jtag_debug_module_end_xfer = ~(cpu_jtag_debug_module_waits_for_read | cpu_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_jtag_debug_module = cpu_jtag_debug_module_end_xfer & (~cpu_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & cpu_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests);

  //cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_jtag_debug_module_arb_counter_enable)
          cpu_jtag_debug_module_arb_share_counter <= cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests))
          cpu_jtag_debug_module_slavearbiterlockenable <= |cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu/data_master cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & cpu_data_master_continuerequest;

  //cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_jtag_debug_module_slavearbiterlockenable2 = |cpu_jtag_debug_module_arb_share_counter_next_value;

  //cpu/data_master cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted cpu/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module <= cpu_instruction_master_saved_grant_cpu_jtag_debug_module ? 1 : (cpu_jtag_debug_module_arbitration_holdoff_internal | ~cpu_instruction_master_requests_cpu_jtag_debug_module) ? 0 : last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_cpu_jtag_debug_module & cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_jtag_debug_module_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_cpu_jtag_debug_module = cpu_data_master_requests_cpu_jtag_debug_module & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register))) | cpu_instruction_master_arbiterlock);
  //local readdatavalid cpu_data_master_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign cpu_data_master_read_data_valid_cpu_jtag_debug_module = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_read & ~cpu_jtag_debug_module_waits_for_read;

  //cpu_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_jtag_debug_module_writedata = cpu_data_master_writedata;

  assign cpu_instruction_master_requests_cpu_jtag_debug_module = (({cpu_instruction_master_address_to_slave[28 : 11] , 11'b0} == 29'h1001800) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted cpu/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module <= cpu_data_master_saved_grant_cpu_jtag_debug_module ? 1 : (cpu_jtag_debug_module_arbitration_holdoff_internal | ~cpu_data_master_requests_cpu_jtag_debug_module) ? 0 : last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_cpu_jtag_debug_module & cpu_data_master_requests_cpu_jtag_debug_module;

  assign cpu_instruction_master_qualified_request_cpu_jtag_debug_module = cpu_instruction_master_requests_cpu_jtag_debug_module & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (|cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register) | (|cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register))) | cpu_data_master_arbiterlock);
  //local readdatavalid cpu_instruction_master_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign cpu_instruction_master_read_data_valid_cpu_jtag_debug_module = cpu_instruction_master_granted_cpu_jtag_debug_module & cpu_instruction_master_read & ~cpu_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_master_qreq_vector[0] = cpu_instruction_master_qualified_request_cpu_jtag_debug_module;

  //cpu/instruction_master grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_instruction_master_granted_cpu_jtag_debug_module = cpu_jtag_debug_module_grant_vector[0];

  //cpu/instruction_master saved-grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_instruction_master_saved_grant_cpu_jtag_debug_module = cpu_jtag_debug_module_arb_winner[0] && cpu_instruction_master_requests_cpu_jtag_debug_module;

  //cpu/data_master assignment into master qualified-requests vector for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_master_qreq_vector[1] = cpu_data_master_qualified_request_cpu_jtag_debug_module;

  //cpu/data_master grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_data_master_granted_cpu_jtag_debug_module = cpu_jtag_debug_module_grant_vector[1];

  //cpu/data_master saved-grant cpu/jtag_debug_module, which is an e_assign
  assign cpu_data_master_saved_grant_cpu_jtag_debug_module = cpu_jtag_debug_module_arb_winner[1] && cpu_data_master_requests_cpu_jtag_debug_module;

  //cpu/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_jtag_debug_module_chosen_master_double_vector = {cpu_jtag_debug_module_master_qreq_vector, cpu_jtag_debug_module_master_qreq_vector} & ({~cpu_jtag_debug_module_master_qreq_vector, ~cpu_jtag_debug_module_master_qreq_vector} + cpu_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_jtag_debug_module_arb_winner = (cpu_jtag_debug_module_allow_new_arb_cycle & | cpu_jtag_debug_module_grant_vector) ? cpu_jtag_debug_module_grant_vector : cpu_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_jtag_debug_module_allow_new_arb_cycle)
          cpu_jtag_debug_module_saved_chosen_master_vector <= |cpu_jtag_debug_module_grant_vector ? cpu_jtag_debug_module_grant_vector : cpu_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_jtag_debug_module_grant_vector = {(cpu_jtag_debug_module_chosen_master_double_vector[1] | cpu_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_jtag_debug_module_chosen_master_double_vector[0] | cpu_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_jtag_debug_module_chosen_master_rot_left = (cpu_jtag_debug_module_arb_winner << 1) ? (cpu_jtag_debug_module_arb_winner << 1) : 1;

  //cpu/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_jtag_debug_module_grant_vector)
          cpu_jtag_debug_module_arb_addend <= cpu_jtag_debug_module_end_xfer? cpu_jtag_debug_module_chosen_master_rot_left : cpu_jtag_debug_module_grant_vector;
    end


  assign cpu_jtag_debug_module_begintransfer = cpu_jtag_debug_module_begins_xfer;
  //cpu_jtag_debug_module_reset_n assignment, which is an e_assign
  assign cpu_jtag_debug_module_reset_n = reset_n;

  //assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest;

  assign cpu_jtag_debug_module_chipselect = cpu_data_master_granted_cpu_jtag_debug_module | cpu_instruction_master_granted_cpu_jtag_debug_module;
  //cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_firsttransfer = cpu_jtag_debug_module_begins_xfer ? cpu_jtag_debug_module_unreg_firsttransfer : cpu_jtag_debug_module_reg_firsttransfer;

  //cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_unreg_firsttransfer = ~(cpu_jtag_debug_module_slavearbiterlockenable & cpu_jtag_debug_module_any_continuerequest);

  //cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_jtag_debug_module_begins_xfer)
          cpu_jtag_debug_module_reg_firsttransfer <= cpu_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_jtag_debug_module_beginbursttransfer_internal = cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_jtag_debug_module_arbitration_holdoff_internal = cpu_jtag_debug_module_begins_xfer & cpu_jtag_debug_module_firsttransfer;

  //cpu_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_jtag_debug_module_write = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_write;

  assign shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master = cpu_data_master_address_to_slave;
  //cpu_jtag_debug_module_address mux, which is an e_mux
  assign cpu_jtag_debug_module_address = (cpu_data_master_granted_cpu_jtag_debug_module)? (shifted_address_to_cpu_jtag_debug_module_from_cpu_data_master >> 2) :
    (shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master >> 2);

  assign shifted_address_to_cpu_jtag_debug_module_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  //d1_cpu_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_jtag_debug_module_end_xfer <= cpu_jtag_debug_module_end_xfer;
    end


  //cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_read = cpu_jtag_debug_module_in_a_read_cycle & cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_read_cycle = (cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_read) | (cpu_instruction_master_granted_cpu_jtag_debug_module & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_jtag_debug_module_in_a_read_cycle;

  //cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_write = cpu_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_write_cycle = cpu_data_master_granted_cpu_jtag_debug_module & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_jtag_debug_module_counter = 0;
  //cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_jtag_debug_module_byteenable = (cpu_data_master_granted_cpu_jtag_debug_module)? cpu_data_master_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_jtag_debug_module_debugaccess = (cpu_data_master_granted_cpu_jtag_debug_module)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_cpu_jtag_debug_module + cpu_instruction_master_granted_cpu_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_cpu_jtag_debug_module + cpu_instruction_master_saved_grant_cpu_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module button_pio_s1_irq_from_sa_clock_crossing_cpu_data_master_module (
                                                                         // inputs:
                                                                          clk,
                                                                          data_in,
                                                                          reset_n,

                                                                         // outputs:
                                                                          data_out
                                                                       )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module high_res_timer_s1_irq_from_sa_clock_crossing_cpu_data_master_module (
                                                                             // inputs:
                                                                              clk,
                                                                              data_in,
                                                                              reset_n,

                                                                             // outputs:
                                                                              data_out
                                                                           )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_data_master_module (
                                                                                       // inputs:
                                                                                        clk,
                                                                                        data_in,
                                                                                        reset_n,

                                                                                       // outputs:
                                                                                        data_out
                                                                                     )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sys_clk_timer_s1_irq_from_sa_clock_crossing_cpu_data_master_module (
                                                                            // inputs:
                                                                             clk,
                                                                             data_in,
                                                                             reset_n,

                                                                            // outputs:
                                                                             data_out
                                                                          )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_data_master_arbitrator (
                                    // inputs:
                                     button_pio_s1_irq_from_sa,
                                     clk,
                                     cpu_data_master_address,
                                     cpu_data_master_byteenable,
                                     cpu_data_master_granted_cpu_ddr_clock_bridge_s1,
                                     cpu_data_master_granted_cpu_jtag_debug_module,
                                     cpu_data_master_granted_descriptor_memory_s1,
                                     cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1,
                                     cpu_data_master_granted_sgdma_rx_csr,
                                     cpu_data_master_granted_sgdma_tx_csr,
                                     cpu_data_master_granted_slow_peripheral_bridge_s1,
                                     cpu_data_master_granted_tse_mac_control_port,
                                     cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1,
                                     cpu_data_master_qualified_request_cpu_jtag_debug_module,
                                     cpu_data_master_qualified_request_descriptor_memory_s1,
                                     cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1,
                                     cpu_data_master_qualified_request_sgdma_rx_csr,
                                     cpu_data_master_qualified_request_sgdma_tx_csr,
                                     cpu_data_master_qualified_request_slow_peripheral_bridge_s1,
                                     cpu_data_master_qualified_request_tse_mac_control_port,
                                     cpu_data_master_read,
                                     cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1,
                                     cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                     cpu_data_master_read_data_valid_cpu_jtag_debug_module,
                                     cpu_data_master_read_data_valid_descriptor_memory_s1,
                                     cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1,
                                     cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                     cpu_data_master_read_data_valid_sgdma_rx_csr,
                                     cpu_data_master_read_data_valid_sgdma_tx_csr,
                                     cpu_data_master_read_data_valid_slow_peripheral_bridge_s1,
                                     cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register,
                                     cpu_data_master_read_data_valid_tse_mac_control_port,
                                     cpu_data_master_requests_cpu_ddr_clock_bridge_s1,
                                     cpu_data_master_requests_cpu_jtag_debug_module,
                                     cpu_data_master_requests_descriptor_memory_s1,
                                     cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1,
                                     cpu_data_master_requests_sgdma_rx_csr,
                                     cpu_data_master_requests_sgdma_tx_csr,
                                     cpu_data_master_requests_slow_peripheral_bridge_s1,
                                     cpu_data_master_requests_tse_mac_control_port,
                                     cpu_data_master_write,
                                     cpu_data_master_writedata,
                                     cpu_ddr_clock_bridge_s1_readdata_from_sa,
                                     cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
                                     cpu_jtag_debug_module_readdata_from_sa,
                                     d1_cpu_ddr_clock_bridge_s1_end_xfer,
                                     d1_cpu_jtag_debug_module_end_xfer,
                                     d1_descriptor_memory_s1_end_xfer,
                                     d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer,
                                     d1_sgdma_rx_csr_end_xfer,
                                     d1_sgdma_tx_csr_end_xfer,
                                     d1_slow_peripheral_bridge_s1_end_xfer,
                                     d1_tse_mac_control_port_end_xfer,
                                     descriptor_memory_s1_readdata_from_sa,
                                     high_res_timer_s1_irq_from_sa,
                                     jtag_uart_avalon_jtag_slave_irq_from_sa,
                                     pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa,
                                     pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa,
                                     pll_c0_out,
                                     pll_c0_out_reset_n,
                                     reset_n,
                                     sgdma_rx_csr_irq_from_sa,
                                     sgdma_rx_csr_readdata_from_sa,
                                     sgdma_tx_csr_irq_from_sa,
                                     sgdma_tx_csr_readdata_from_sa,
                                     slow_peripheral_bridge_s1_readdata_from_sa,
                                     slow_peripheral_bridge_s1_waitrequest_from_sa,
                                     sys_clk_timer_s1_irq_from_sa,
                                     tse_mac_control_port_readdata_from_sa,
                                     tse_mac_control_port_waitrequest_from_sa,

                                    // outputs:
                                     cpu_data_master_address_to_slave,
                                     cpu_data_master_irq,
                                     cpu_data_master_latency_counter,
                                     cpu_data_master_readdata,
                                     cpu_data_master_readdatavalid,
                                     cpu_data_master_waitrequest
                                  )
;

  output  [ 28: 0] cpu_data_master_address_to_slave;
  output  [ 31: 0] cpu_data_master_irq;
  output           cpu_data_master_latency_counter;
  output  [ 31: 0] cpu_data_master_readdata;
  output           cpu_data_master_readdatavalid;
  output           cpu_data_master_waitrequest;
  input            button_pio_s1_irq_from_sa;
  input            clk;
  input   [ 28: 0] cpu_data_master_address;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_granted_cpu_ddr_clock_bridge_s1;
  input            cpu_data_master_granted_cpu_jtag_debug_module;
  input            cpu_data_master_granted_descriptor_memory_s1;
  input            cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1;
  input            cpu_data_master_granted_sgdma_rx_csr;
  input            cpu_data_master_granted_sgdma_tx_csr;
  input            cpu_data_master_granted_slow_peripheral_bridge_s1;
  input            cpu_data_master_granted_tse_mac_control_port;
  input            cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1;
  input            cpu_data_master_qualified_request_cpu_jtag_debug_module;
  input            cpu_data_master_qualified_request_descriptor_memory_s1;
  input            cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1;
  input            cpu_data_master_qualified_request_sgdma_rx_csr;
  input            cpu_data_master_qualified_request_sgdma_tx_csr;
  input            cpu_data_master_qualified_request_slow_peripheral_bridge_s1;
  input            cpu_data_master_qualified_request_tse_mac_control_port;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1;
  input            cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  input            cpu_data_master_read_data_valid_descriptor_memory_s1;
  input            cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1;
  input            cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_sgdma_rx_csr;
  input            cpu_data_master_read_data_valid_sgdma_tx_csr;
  input            cpu_data_master_read_data_valid_slow_peripheral_bridge_s1;
  input            cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_tse_mac_control_port;
  input            cpu_data_master_requests_cpu_ddr_clock_bridge_s1;
  input            cpu_data_master_requests_cpu_jtag_debug_module;
  input            cpu_data_master_requests_descriptor_memory_s1;
  input            cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1;
  input            cpu_data_master_requests_sgdma_rx_csr;
  input            cpu_data_master_requests_sgdma_tx_csr;
  input            cpu_data_master_requests_slow_peripheral_bridge_s1;
  input            cpu_data_master_requests_tse_mac_control_port;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 31: 0] cpu_ddr_clock_bridge_s1_readdata_from_sa;
  input            cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_ddr_clock_bridge_s1_end_xfer;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            d1_descriptor_memory_s1_end_xfer;
  input            d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer;
  input            d1_sgdma_rx_csr_end_xfer;
  input            d1_sgdma_tx_csr_end_xfer;
  input            d1_slow_peripheral_bridge_s1_end_xfer;
  input            d1_tse_mac_control_port_end_xfer;
  input   [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  input            high_res_timer_s1_irq_from_sa;
  input            jtag_uart_avalon_jtag_slave_irq_from_sa;
  input   [ 31: 0] pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa;
  input            pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa;
  input            pll_c0_out;
  input            pll_c0_out_reset_n;
  input            reset_n;
  input            sgdma_rx_csr_irq_from_sa;
  input   [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  input            sgdma_tx_csr_irq_from_sa;
  input   [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  input   [ 31: 0] slow_peripheral_bridge_s1_readdata_from_sa;
  input            slow_peripheral_bridge_s1_waitrequest_from_sa;
  input            sys_clk_timer_s1_irq_from_sa;
  input   [ 31: 0] tse_mac_control_port_readdata_from_sa;
  input            tse_mac_control_port_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 28: 0] cpu_data_master_address_last_time;
  wire    [ 28: 0] cpu_data_master_address_to_slave;
  reg     [  3: 0] cpu_data_master_byteenable_last_time;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_is_granted_some_slave;
  reg              cpu_data_master_latency_counter;
  reg              cpu_data_master_read_but_no_slave_selected;
  reg              cpu_data_master_read_last_time;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_run;
  wire             cpu_data_master_waitrequest;
  reg              cpu_data_master_write_last_time;
  reg     [ 31: 0] cpu_data_master_writedata_last_time;
  wire             latency_load_value;
  wire             p1_cpu_data_master_latency_counter;
  wire             pll_c0_out_button_pio_s1_irq_from_sa;
  wire             pll_c0_out_high_res_timer_s1_irq_from_sa;
  wire             pll_c0_out_jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             pll_c0_out_sys_clk_timer_s1_irq_from_sa;
  wire             pre_flush_cpu_data_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_requests_cpu_jtag_debug_module) & (cpu_data_master_granted_cpu_jtag_debug_module | ~cpu_data_master_qualified_request_cpu_jtag_debug_module) & ((~cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_read | (1 & ~d1_cpu_jtag_debug_module_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_cpu_jtag_debug_module | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1 | ~cpu_data_master_requests_cpu_ddr_clock_bridge_s1) & (cpu_data_master_granted_cpu_ddr_clock_bridge_s1 | ~cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1) & ((~cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~cpu_ddr_clock_bridge_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~cpu_ddr_clock_bridge_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_descriptor_memory_s1 | ~cpu_data_master_requests_descriptor_memory_s1) & (cpu_data_master_granted_descriptor_memory_s1 | ~cpu_data_master_qualified_request_descriptor_memory_s1) & ((~cpu_data_master_qualified_request_descriptor_memory_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_descriptor_memory_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & (cpu_data_master_read | cpu_data_master_write))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_data_master_run = r_0 & r_1 & r_2;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1 | ~cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1) & (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1 | ~cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1) & ((~cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_sgdma_rx_csr | ~cpu_data_master_requests_sgdma_rx_csr) & ((~cpu_data_master_qualified_request_sgdma_rx_csr | ~cpu_data_master_read | (1 & ~d1_sgdma_rx_csr_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_sgdma_rx_csr | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_sgdma_tx_csr | ~cpu_data_master_requests_sgdma_tx_csr) & ((~cpu_data_master_qualified_request_sgdma_tx_csr | ~cpu_data_master_read | (1 & ~d1_sgdma_tx_csr_end_xfer & cpu_data_master_read))) & ((~cpu_data_master_qualified_request_sgdma_tx_csr | ~cpu_data_master_write | (1 & cpu_data_master_write))) & 1 & (cpu_data_master_qualified_request_slow_peripheral_bridge_s1 | ~cpu_data_master_requests_slow_peripheral_bridge_s1) & ((~cpu_data_master_qualified_request_slow_peripheral_bridge_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~slow_peripheral_bridge_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_slow_peripheral_bridge_s1 | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~slow_peripheral_bridge_s1_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write))));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_data_master_qualified_request_tse_mac_control_port | ~cpu_data_master_requests_tse_mac_control_port) & ((~cpu_data_master_qualified_request_tse_mac_control_port | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~tse_mac_control_port_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_tse_mac_control_port | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~tse_mac_control_port_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write))));

  //button_pio_s1_irq_from_sa from pll_c2_out to pll_c0_out
  button_pio_s1_irq_from_sa_clock_crossing_cpu_data_master_module button_pio_s1_irq_from_sa_clock_crossing_cpu_data_master
    (
      .clk      (pll_c0_out),
      .data_in  (button_pio_s1_irq_from_sa),
      .data_out (pll_c0_out_button_pio_s1_irq_from_sa),
      .reset_n  (pll_c0_out_reset_n)
    );

  //irq assign, which is an e_assign
  assign cpu_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    pll_c0_out_high_res_timer_s1_irq_from_sa,
    pll_c0_out_button_pio_s1_irq_from_sa,
    pll_c0_out_jtag_uart_avalon_jtag_slave_irq_from_sa,
    pll_c0_out_sys_clk_timer_s1_irq_from_sa,
    sgdma_tx_csr_irq_from_sa,
    sgdma_rx_csr_irq_from_sa};

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_data_master_address_to_slave = cpu_data_master_address[28 : 0];

  //cpu_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_data_master_read_but_no_slave_selected <= cpu_data_master_read & cpu_data_master_run & ~cpu_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_data_master_is_granted_some_slave = cpu_data_master_granted_cpu_jtag_debug_module |
    cpu_data_master_granted_cpu_ddr_clock_bridge_s1 |
    cpu_data_master_granted_descriptor_memory_s1 |
    cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1 |
    cpu_data_master_granted_sgdma_rx_csr |
    cpu_data_master_granted_sgdma_tx_csr |
    cpu_data_master_granted_slow_peripheral_bridge_s1 |
    cpu_data_master_granted_tse_mac_control_port;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_data_master_readdatavalid = cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 |
    cpu_data_master_read_data_valid_descriptor_memory_s1 |
    cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1 |
    cpu_data_master_read_data_valid_slow_peripheral_bridge_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_data_master_readdatavalid = cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_cpu_jtag_debug_module |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_sgdma_rx_csr |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_sgdma_tx_csr |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_data_valid_tse_mac_control_port;

  //cpu/data_master readdata mux, which is an e_mux
  assign cpu_data_master_readdata = ({32 {~(cpu_data_master_qualified_request_cpu_jtag_debug_module & cpu_data_master_read)}} | cpu_jtag_debug_module_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1}} | cpu_ddr_clock_bridge_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_descriptor_memory_s1}} | descriptor_memory_s1_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1}} | pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_sgdma_rx_csr & cpu_data_master_read)}} | sgdma_rx_csr_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_sgdma_tx_csr & cpu_data_master_read)}} | sgdma_tx_csr_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_slow_peripheral_bridge_s1}} | slow_peripheral_bridge_s1_readdata_from_sa) &
    ({32 {~(cpu_data_master_qualified_request_tse_mac_control_port & cpu_data_master_read)}} | tse_mac_control_port_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_data_master_waitrequest = ~cpu_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_latency_counter <= 0;
      else 
        cpu_data_master_latency_counter <= p1_cpu_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_data_master_latency_counter = ((cpu_data_master_run & cpu_data_master_read))? latency_load_value :
    (cpu_data_master_latency_counter)? cpu_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {cpu_data_master_requests_descriptor_memory_s1}} & 1;

  //high_res_timer_s1_irq_from_sa from pll_c2_out to pll_c0_out
  high_res_timer_s1_irq_from_sa_clock_crossing_cpu_data_master_module high_res_timer_s1_irq_from_sa_clock_crossing_cpu_data_master
    (
      .clk      (pll_c0_out),
      .data_in  (high_res_timer_s1_irq_from_sa),
      .data_out (pll_c0_out_high_res_timer_s1_irq_from_sa),
      .reset_n  (pll_c0_out_reset_n)
    );

  //jtag_uart_avalon_jtag_slave_irq_from_sa from pll_c2_out to pll_c0_out
  jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_data_master_module jtag_uart_avalon_jtag_slave_irq_from_sa_clock_crossing_cpu_data_master
    (
      .clk      (pll_c0_out),
      .data_in  (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .data_out (pll_c0_out_jtag_uart_avalon_jtag_slave_irq_from_sa),
      .reset_n  (pll_c0_out_reset_n)
    );

  //sys_clk_timer_s1_irq_from_sa from pll_c2_out to pll_c0_out
  sys_clk_timer_s1_irq_from_sa_clock_crossing_cpu_data_master_module sys_clk_timer_s1_irq_from_sa_clock_crossing_cpu_data_master
    (
      .clk      (pll_c0_out),
      .data_in  (sys_clk_timer_s1_irq_from_sa),
      .data_out (pll_c0_out_sys_clk_timer_s1_irq_from_sa),
      .reset_n  (pll_c0_out_reset_n)
    );


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_address_last_time <= 0;
      else 
        cpu_data_master_address_last_time <= cpu_data_master_address;
    end


  //cpu/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_data_master_waitrequest & (cpu_data_master_read | cpu_data_master_write);
    end


  //cpu_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_address != cpu_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_byteenable_last_time <= 0;
      else 
        cpu_data_master_byteenable_last_time <= cpu_data_master_byteenable;
    end


  //cpu_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_byteenable != cpu_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_last_time <= 0;
      else 
        cpu_data_master_read_last_time <= cpu_data_master_read;
    end


  //cpu_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_read != cpu_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_write_last_time <= 0;
      else 
        cpu_data_master_write_last_time <= cpu_data_master_write;
    end


  //cpu_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_write != cpu_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_writedata_last_time <= 0;
      else 
        cpu_data_master_writedata_last_time <= cpu_data_master_writedata;
    end


  //cpu_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_writedata != cpu_data_master_writedata_last_time) & cpu_data_master_write)
        begin
          $write("%0d ns: cpu_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_instruction_master_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_ddr_clock_bridge_s1_readdata_from_sa,
                                            cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
                                            cpu_instruction_master_address,
                                            cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1,
                                            cpu_instruction_master_granted_cpu_jtag_debug_module,
                                            cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1,
                                            cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1,
                                            cpu_instruction_master_qualified_request_cpu_jtag_debug_module,
                                            cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1,
                                            cpu_instruction_master_read,
                                            cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1,
                                            cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                            cpu_instruction_master_read_data_valid_cpu_jtag_debug_module,
                                            cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1,
                                            cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                            cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1,
                                            cpu_instruction_master_requests_cpu_jtag_debug_module,
                                            cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1,
                                            cpu_jtag_debug_module_readdata_from_sa,
                                            d1_cpu_ddr_clock_bridge_s1_end_xfer,
                                            d1_cpu_jtag_debug_module_end_xfer,
                                            d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer,
                                            pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa,
                                            pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa,
                                            reset_n,

                                           // outputs:
                                            cpu_instruction_master_address_to_slave,
                                            cpu_instruction_master_latency_counter,
                                            cpu_instruction_master_readdata,
                                            cpu_instruction_master_readdatavalid,
                                            cpu_instruction_master_waitrequest
                                         )
;

  output  [ 28: 0] cpu_instruction_master_address_to_slave;
  output           cpu_instruction_master_latency_counter;
  output  [ 31: 0] cpu_instruction_master_readdata;
  output           cpu_instruction_master_readdatavalid;
  output           cpu_instruction_master_waitrequest;
  input            clk;
  input   [ 31: 0] cpu_ddr_clock_bridge_s1_readdata_from_sa;
  input            cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  input   [ 28: 0] cpu_instruction_master_address;
  input            cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1;
  input            cpu_instruction_master_granted_cpu_jtag_debug_module;
  input            cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1;
  input            cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1;
  input            cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  input            cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1;
  input            cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  input            cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1;
  input            cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input            cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  input            cpu_instruction_master_requests_cpu_jtag_debug_module;
  input            cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_ddr_clock_bridge_s1_end_xfer;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer;
  input   [ 31: 0] pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa;
  input            pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 28: 0] cpu_instruction_master_address_last_time;
  wire    [ 28: 0] cpu_instruction_master_address_to_slave;
  wire             cpu_instruction_master_is_granted_some_slave;
  reg              cpu_instruction_master_latency_counter;
  reg              cpu_instruction_master_read_but_no_slave_selected;
  reg              cpu_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_run;
  wire             cpu_instruction_master_waitrequest;
  wire             latency_load_value;
  wire             p1_cpu_instruction_master_latency_counter;
  wire             pre_flush_cpu_instruction_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_instruction_master_qualified_request_cpu_jtag_debug_module | ~cpu_instruction_master_requests_cpu_jtag_debug_module) & (cpu_instruction_master_granted_cpu_jtag_debug_module | ~cpu_instruction_master_qualified_request_cpu_jtag_debug_module) & ((~cpu_instruction_master_qualified_request_cpu_jtag_debug_module | ~cpu_instruction_master_read | (1 & ~d1_cpu_jtag_debug_module_end_xfer & cpu_instruction_master_read))) & 1 & (cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 | ~cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1) & (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1 | ~cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1) & ((~cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 | ~(cpu_instruction_master_read) | (1 & ~cpu_ddr_clock_bridge_s1_waitrequest_from_sa & (cpu_instruction_master_read))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_instruction_master_run = r_0 & r_1;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1 | ~cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1) & (cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1 | ~cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1) & ((~cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1 | ~(cpu_instruction_master_read) | (1 & ~pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa & (cpu_instruction_master_read))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_instruction_master_address_to_slave = cpu_instruction_master_address[28 : 0];

  //cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_instruction_master_read_but_no_slave_selected <= cpu_instruction_master_read & cpu_instruction_master_run & ~cpu_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_instruction_master_is_granted_some_slave = cpu_instruction_master_granted_cpu_jtag_debug_module |
    cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1 |
    cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_instruction_master_readdatavalid = cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 |
    cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_instruction_master_readdatavalid = cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_data_valid_cpu_jtag_debug_module |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid;

  //cpu/instruction_master readdata mux, which is an e_mux
  assign cpu_instruction_master_readdata = ({32 {~(cpu_instruction_master_qualified_request_cpu_jtag_debug_module & cpu_instruction_master_read)}} | cpu_jtag_debug_module_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1}} | cpu_ddr_clock_bridge_s1_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1}} | pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_instruction_master_waitrequest = ~cpu_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_latency_counter <= 0;
      else 
        cpu_instruction_master_latency_counter <= p1_cpu_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_instruction_master_latency_counter = ((cpu_instruction_master_run & cpu_instruction_master_read))? latency_load_value :
    (cpu_instruction_master_latency_counter)? cpu_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_address_last_time <= 0;
      else 
        cpu_instruction_master_address_last_time <= cpu_instruction_master_address;
    end


  //cpu/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_instruction_master_waitrequest & (cpu_instruction_master_read);
    end


  //cpu_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_address != cpu_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_last_time <= 0;
      else 
        cpu_instruction_master_read_last_time <= cpu_instruction_master_read;
    end


  //cpu_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_read != cpu_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_cpu_ddr_clock_bridge_s1_module (
                                                                        // inputs:
                                                                         clear_fifo,
                                                                         clk,
                                                                         data_in,
                                                                         read,
                                                                         reset_n,
                                                                         sync_reset,
                                                                         write,

                                                                        // outputs:
                                                                         data_out,
                                                                         empty,
                                                                         fifo_contains_ones_n,
                                                                         full
                                                                      )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  wire             full_48;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_47;
  assign empty = !full_0;
  assign full_48 = 0;
  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    0;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_cpu_ddr_clock_bridge_s1_module (
                                                                               // inputs:
                                                                                clear_fifo,
                                                                                clk,
                                                                                data_in,
                                                                                read,
                                                                                reset_n,
                                                                                sync_reset,
                                                                                write,

                                                                               // outputs:
                                                                                data_out,
                                                                                empty,
                                                                                fifo_contains_ones_n,
                                                                                full
                                                                             )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  wire             full_48;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_47;
  assign empty = !full_0;
  assign full_48 = 0;
  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    0;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_sgdma_tx_m_read_to_cpu_ddr_clock_bridge_s1_module (
                                                                        // inputs:
                                                                         clear_fifo,
                                                                         clk,
                                                                         data_in,
                                                                         read,
                                                                         reset_n,
                                                                         sync_reset,
                                                                         write,

                                                                        // outputs:
                                                                         data_out,
                                                                         empty,
                                                                         fifo_contains_ones_n,
                                                                         full
                                                                      )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  reg              full_33;
  reg              full_34;
  reg              full_35;
  reg              full_36;
  reg              full_37;
  reg              full_38;
  reg              full_39;
  reg              full_4;
  reg              full_40;
  reg              full_41;
  reg              full_42;
  reg              full_43;
  reg              full_44;
  reg              full_45;
  reg              full_46;
  reg              full_47;
  wire             full_48;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p33_full_33;
  wire             p33_stage_33;
  wire             p34_full_34;
  wire             p34_stage_34;
  wire             p35_full_35;
  wire             p35_stage_35;
  wire             p36_full_36;
  wire             p36_stage_36;
  wire             p37_full_37;
  wire             p37_stage_37;
  wire             p38_full_38;
  wire             p38_stage_38;
  wire             p39_full_39;
  wire             p39_stage_39;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p40_full_40;
  wire             p40_stage_40;
  wire             p41_full_41;
  wire             p41_stage_41;
  wire             p42_full_42;
  wire             p42_stage_42;
  wire             p43_full_43;
  wire             p43_stage_43;
  wire             p44_full_44;
  wire             p44_stage_44;
  wire             p45_full_45;
  wire             p45_stage_45;
  wire             p46_full_46;
  wire             p46_stage_46;
  wire             p47_full_47;
  wire             p47_stage_47;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_33;
  reg              stage_34;
  reg              stage_35;
  reg              stage_36;
  reg              stage_37;
  reg              stage_38;
  reg              stage_39;
  reg              stage_4;
  reg              stage_40;
  reg              stage_41;
  reg              stage_42;
  reg              stage_43;
  reg              stage_44;
  reg              stage_45;
  reg              stage_46;
  reg              stage_47;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_47;
  assign empty = !full_0;
  assign full_48 = 0;
  //data_47, which is an e_mux
  assign p47_stage_47 = ((full_48 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_47 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_47))
          if (sync_reset & full_47 & !((full_48 == 0) & read & write))
              stage_47 <= 0;
          else 
            stage_47 <= p47_stage_47;
    end


  //control_47, which is an e_mux
  assign p47_full_47 = ((read & !write) == 0)? full_46 :
    0;

  //control_reg_47, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_47 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_47 <= 0;
          else 
            full_47 <= p47_full_47;
    end


  //data_46, which is an e_mux
  assign p46_stage_46 = ((full_47 & ~clear_fifo) == 0)? data_in :
    stage_47;

  //data_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_46 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_46))
          if (sync_reset & full_46 & !((full_47 == 0) & read & write))
              stage_46 <= 0;
          else 
            stage_46 <= p46_stage_46;
    end


  //control_46, which is an e_mux
  assign p46_full_46 = ((read & !write) == 0)? full_45 :
    full_47;

  //control_reg_46, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_46 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_46 <= 0;
          else 
            full_46 <= p46_full_46;
    end


  //data_45, which is an e_mux
  assign p45_stage_45 = ((full_46 & ~clear_fifo) == 0)? data_in :
    stage_46;

  //data_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_45 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_45))
          if (sync_reset & full_45 & !((full_46 == 0) & read & write))
              stage_45 <= 0;
          else 
            stage_45 <= p45_stage_45;
    end


  //control_45, which is an e_mux
  assign p45_full_45 = ((read & !write) == 0)? full_44 :
    full_46;

  //control_reg_45, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_45 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_45 <= 0;
          else 
            full_45 <= p45_full_45;
    end


  //data_44, which is an e_mux
  assign p44_stage_44 = ((full_45 & ~clear_fifo) == 0)? data_in :
    stage_45;

  //data_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_44 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_44))
          if (sync_reset & full_44 & !((full_45 == 0) & read & write))
              stage_44 <= 0;
          else 
            stage_44 <= p44_stage_44;
    end


  //control_44, which is an e_mux
  assign p44_full_44 = ((read & !write) == 0)? full_43 :
    full_45;

  //control_reg_44, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_44 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_44 <= 0;
          else 
            full_44 <= p44_full_44;
    end


  //data_43, which is an e_mux
  assign p43_stage_43 = ((full_44 & ~clear_fifo) == 0)? data_in :
    stage_44;

  //data_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_43 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_43))
          if (sync_reset & full_43 & !((full_44 == 0) & read & write))
              stage_43 <= 0;
          else 
            stage_43 <= p43_stage_43;
    end


  //control_43, which is an e_mux
  assign p43_full_43 = ((read & !write) == 0)? full_42 :
    full_44;

  //control_reg_43, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_43 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_43 <= 0;
          else 
            full_43 <= p43_full_43;
    end


  //data_42, which is an e_mux
  assign p42_stage_42 = ((full_43 & ~clear_fifo) == 0)? data_in :
    stage_43;

  //data_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_42 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_42))
          if (sync_reset & full_42 & !((full_43 == 0) & read & write))
              stage_42 <= 0;
          else 
            stage_42 <= p42_stage_42;
    end


  //control_42, which is an e_mux
  assign p42_full_42 = ((read & !write) == 0)? full_41 :
    full_43;

  //control_reg_42, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_42 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_42 <= 0;
          else 
            full_42 <= p42_full_42;
    end


  //data_41, which is an e_mux
  assign p41_stage_41 = ((full_42 & ~clear_fifo) == 0)? data_in :
    stage_42;

  //data_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_41 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_41))
          if (sync_reset & full_41 & !((full_42 == 0) & read & write))
              stage_41 <= 0;
          else 
            stage_41 <= p41_stage_41;
    end


  //control_41, which is an e_mux
  assign p41_full_41 = ((read & !write) == 0)? full_40 :
    full_42;

  //control_reg_41, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_41 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_41 <= 0;
          else 
            full_41 <= p41_full_41;
    end


  //data_40, which is an e_mux
  assign p40_stage_40 = ((full_41 & ~clear_fifo) == 0)? data_in :
    stage_41;

  //data_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_40 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_40))
          if (sync_reset & full_40 & !((full_41 == 0) & read & write))
              stage_40 <= 0;
          else 
            stage_40 <= p40_stage_40;
    end


  //control_40, which is an e_mux
  assign p40_full_40 = ((read & !write) == 0)? full_39 :
    full_41;

  //control_reg_40, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_40 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_40 <= 0;
          else 
            full_40 <= p40_full_40;
    end


  //data_39, which is an e_mux
  assign p39_stage_39 = ((full_40 & ~clear_fifo) == 0)? data_in :
    stage_40;

  //data_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_39 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_39))
          if (sync_reset & full_39 & !((full_40 == 0) & read & write))
              stage_39 <= 0;
          else 
            stage_39 <= p39_stage_39;
    end


  //control_39, which is an e_mux
  assign p39_full_39 = ((read & !write) == 0)? full_38 :
    full_40;

  //control_reg_39, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_39 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_39 <= 0;
          else 
            full_39 <= p39_full_39;
    end


  //data_38, which is an e_mux
  assign p38_stage_38 = ((full_39 & ~clear_fifo) == 0)? data_in :
    stage_39;

  //data_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_38 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_38))
          if (sync_reset & full_38 & !((full_39 == 0) & read & write))
              stage_38 <= 0;
          else 
            stage_38 <= p38_stage_38;
    end


  //control_38, which is an e_mux
  assign p38_full_38 = ((read & !write) == 0)? full_37 :
    full_39;

  //control_reg_38, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_38 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_38 <= 0;
          else 
            full_38 <= p38_full_38;
    end


  //data_37, which is an e_mux
  assign p37_stage_37 = ((full_38 & ~clear_fifo) == 0)? data_in :
    stage_38;

  //data_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_37 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_37))
          if (sync_reset & full_37 & !((full_38 == 0) & read & write))
              stage_37 <= 0;
          else 
            stage_37 <= p37_stage_37;
    end


  //control_37, which is an e_mux
  assign p37_full_37 = ((read & !write) == 0)? full_36 :
    full_38;

  //control_reg_37, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_37 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_37 <= 0;
          else 
            full_37 <= p37_full_37;
    end


  //data_36, which is an e_mux
  assign p36_stage_36 = ((full_37 & ~clear_fifo) == 0)? data_in :
    stage_37;

  //data_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_36 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_36))
          if (sync_reset & full_36 & !((full_37 == 0) & read & write))
              stage_36 <= 0;
          else 
            stage_36 <= p36_stage_36;
    end


  //control_36, which is an e_mux
  assign p36_full_36 = ((read & !write) == 0)? full_35 :
    full_37;

  //control_reg_36, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_36 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_36 <= 0;
          else 
            full_36 <= p36_full_36;
    end


  //data_35, which is an e_mux
  assign p35_stage_35 = ((full_36 & ~clear_fifo) == 0)? data_in :
    stage_36;

  //data_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_35 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_35))
          if (sync_reset & full_35 & !((full_36 == 0) & read & write))
              stage_35 <= 0;
          else 
            stage_35 <= p35_stage_35;
    end


  //control_35, which is an e_mux
  assign p35_full_35 = ((read & !write) == 0)? full_34 :
    full_36;

  //control_reg_35, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_35 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_35 <= 0;
          else 
            full_35 <= p35_full_35;
    end


  //data_34, which is an e_mux
  assign p34_stage_34 = ((full_35 & ~clear_fifo) == 0)? data_in :
    stage_35;

  //data_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_34 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_34))
          if (sync_reset & full_34 & !((full_35 == 0) & read & write))
              stage_34 <= 0;
          else 
            stage_34 <= p34_stage_34;
    end


  //control_34, which is an e_mux
  assign p34_full_34 = ((read & !write) == 0)? full_33 :
    full_35;

  //control_reg_34, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_34 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_34 <= 0;
          else 
            full_34 <= p34_full_34;
    end


  //data_33, which is an e_mux
  assign p33_stage_33 = ((full_34 & ~clear_fifo) == 0)? data_in :
    stage_34;

  //data_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_33 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_33))
          if (sync_reset & full_33 & !((full_34 == 0) & read & write))
              stage_33 <= 0;
          else 
            stage_33 <= p33_stage_33;
    end


  //control_33, which is an e_mux
  assign p33_full_33 = ((read & !write) == 0)? full_32 :
    full_34;

  //control_reg_33, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_33 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_33 <= 0;
          else 
            full_33 <= p33_full_33;
    end


  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    stage_33;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    full_33;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_ddr_clock_bridge_s1_arbitrator (
                                            // inputs:
                                             clk,
                                             cpu_data_master_address_to_slave,
                                             cpu_data_master_byteenable,
                                             cpu_data_master_latency_counter,
                                             cpu_data_master_read,
                                             cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                             cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register,
                                             cpu_data_master_write,
                                             cpu_data_master_writedata,
                                             cpu_ddr_clock_bridge_s1_endofpacket,
                                             cpu_ddr_clock_bridge_s1_readdata,
                                             cpu_ddr_clock_bridge_s1_readdatavalid,
                                             cpu_ddr_clock_bridge_s1_waitrequest,
                                             cpu_instruction_master_address_to_slave,
                                             cpu_instruction_master_latency_counter,
                                             cpu_instruction_master_read,
                                             cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                             reset_n,
                                             sgdma_rx_m_write_address_to_slave,
                                             sgdma_rx_m_write_byteenable,
                                             sgdma_rx_m_write_write,
                                             sgdma_rx_m_write_writedata,
                                             sgdma_tx_m_read_address_to_slave,
                                             sgdma_tx_m_read_latency_counter,
                                             sgdma_tx_m_read_read,

                                            // outputs:
                                             cpu_data_master_granted_cpu_ddr_clock_bridge_s1,
                                             cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1,
                                             cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1,
                                             cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                             cpu_data_master_requests_cpu_ddr_clock_bridge_s1,
                                             cpu_ddr_clock_bridge_s1_address,
                                             cpu_ddr_clock_bridge_s1_byteenable,
                                             cpu_ddr_clock_bridge_s1_endofpacket_from_sa,
                                             cpu_ddr_clock_bridge_s1_nativeaddress,
                                             cpu_ddr_clock_bridge_s1_read,
                                             cpu_ddr_clock_bridge_s1_readdata_from_sa,
                                             cpu_ddr_clock_bridge_s1_reset_n,
                                             cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
                                             cpu_ddr_clock_bridge_s1_write,
                                             cpu_ddr_clock_bridge_s1_writedata,
                                             cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1,
                                             cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1,
                                             cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1,
                                             cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                             cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1,
                                             d1_cpu_ddr_clock_bridge_s1_end_xfer,
                                             sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1,
                                             sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1,
                                             sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1,
                                             sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1,
                                             sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1,
                                             sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1,
                                             sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                             sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1
                                          )
;

  output           cpu_data_master_granted_cpu_ddr_clock_bridge_s1;
  output           cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1;
  output           cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1;
  output           cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  output           cpu_data_master_requests_cpu_ddr_clock_bridge_s1;
  output  [ 23: 0] cpu_ddr_clock_bridge_s1_address;
  output  [  3: 0] cpu_ddr_clock_bridge_s1_byteenable;
  output           cpu_ddr_clock_bridge_s1_endofpacket_from_sa;
  output  [ 23: 0] cpu_ddr_clock_bridge_s1_nativeaddress;
  output           cpu_ddr_clock_bridge_s1_read;
  output  [ 31: 0] cpu_ddr_clock_bridge_s1_readdata_from_sa;
  output           cpu_ddr_clock_bridge_s1_reset_n;
  output           cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  output           cpu_ddr_clock_bridge_s1_write;
  output  [ 31: 0] cpu_ddr_clock_bridge_s1_writedata;
  output           cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1;
  output           cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1;
  output           cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1;
  output           cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  output           cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  output           d1_cpu_ddr_clock_bridge_s1_end_xfer;
  output           sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1;
  output           sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1;
  output           sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1;
  output           sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1;
  output           sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1;
  output           sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1;
  output           sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  output           sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            cpu_ddr_clock_bridge_s1_endofpacket;
  input   [ 31: 0] cpu_ddr_clock_bridge_s1_readdata;
  input            cpu_ddr_clock_bridge_s1_readdatavalid;
  input            cpu_ddr_clock_bridge_s1_waitrequest;
  input   [ 28: 0] cpu_instruction_master_address_to_slave;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_m_write_address_to_slave;
  input   [  3: 0] sgdma_rx_m_write_byteenable;
  input            sgdma_rx_m_write_write;
  input   [ 31: 0] sgdma_rx_m_write_writedata;
  input   [ 31: 0] sgdma_tx_m_read_address_to_slave;
  input            sgdma_tx_m_read_latency_counter;
  input            sgdma_tx_m_read_read;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_cpu_ddr_clock_bridge_s1;
  wire             cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1;
  wire             cpu_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  wire             cpu_data_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1;
  wire             cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1;
  wire             cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  wire             cpu_data_master_requests_cpu_ddr_clock_bridge_s1;
  wire             cpu_data_master_saved_grant_cpu_ddr_clock_bridge_s1;
  wire    [ 23: 0] cpu_ddr_clock_bridge_s1_address;
  wire             cpu_ddr_clock_bridge_s1_allgrants;
  wire             cpu_ddr_clock_bridge_s1_allow_new_arb_cycle;
  wire             cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant;
  wire             cpu_ddr_clock_bridge_s1_any_continuerequest;
  reg     [  3: 0] cpu_ddr_clock_bridge_s1_arb_addend;
  wire             cpu_ddr_clock_bridge_s1_arb_counter_enable;
  reg     [  3: 0] cpu_ddr_clock_bridge_s1_arb_share_counter;
  wire    [  3: 0] cpu_ddr_clock_bridge_s1_arb_share_counter_next_value;
  wire    [  3: 0] cpu_ddr_clock_bridge_s1_arb_share_set_values;
  wire    [  3: 0] cpu_ddr_clock_bridge_s1_arb_winner;
  wire             cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal;
  wire             cpu_ddr_clock_bridge_s1_beginbursttransfer_internal;
  wire             cpu_ddr_clock_bridge_s1_begins_xfer;
  wire    [  3: 0] cpu_ddr_clock_bridge_s1_byteenable;
  wire    [  7: 0] cpu_ddr_clock_bridge_s1_chosen_master_double_vector;
  wire    [  3: 0] cpu_ddr_clock_bridge_s1_chosen_master_rot_left;
  wire             cpu_ddr_clock_bridge_s1_end_xfer;
  wire             cpu_ddr_clock_bridge_s1_endofpacket_from_sa;
  wire             cpu_ddr_clock_bridge_s1_firsttransfer;
  wire    [  3: 0] cpu_ddr_clock_bridge_s1_grant_vector;
  wire             cpu_ddr_clock_bridge_s1_in_a_read_cycle;
  wire             cpu_ddr_clock_bridge_s1_in_a_write_cycle;
  wire    [  3: 0] cpu_ddr_clock_bridge_s1_master_qreq_vector;
  wire             cpu_ddr_clock_bridge_s1_move_on_to_next_transaction;
  wire    [ 23: 0] cpu_ddr_clock_bridge_s1_nativeaddress;
  wire             cpu_ddr_clock_bridge_s1_non_bursting_master_requests;
  wire             cpu_ddr_clock_bridge_s1_read;
  wire    [ 31: 0] cpu_ddr_clock_bridge_s1_readdata_from_sa;
  wire             cpu_ddr_clock_bridge_s1_readdatavalid_from_sa;
  reg              cpu_ddr_clock_bridge_s1_reg_firsttransfer;
  wire             cpu_ddr_clock_bridge_s1_reset_n;
  reg     [  3: 0] cpu_ddr_clock_bridge_s1_saved_chosen_master_vector;
  reg              cpu_ddr_clock_bridge_s1_slavearbiterlockenable;
  wire             cpu_ddr_clock_bridge_s1_slavearbiterlockenable2;
  wire             cpu_ddr_clock_bridge_s1_unreg_firsttransfer;
  wire             cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  wire             cpu_ddr_clock_bridge_s1_waits_for_read;
  wire             cpu_ddr_clock_bridge_s1_waits_for_write;
  wire             cpu_ddr_clock_bridge_s1_write;
  wire    [ 31: 0] cpu_ddr_clock_bridge_s1_writedata;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1;
  wire             cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1;
  wire             cpu_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  wire             cpu_instruction_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1;
  wire             cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1;
  wire             cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  wire             cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  wire             cpu_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1;
  reg              d1_cpu_ddr_clock_bridge_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_cpu_ddr_clock_bridge_s1;
  reg              last_cycle_cpu_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1;
  reg              last_cycle_sgdma_rx_m_write_granted_slave_cpu_ddr_clock_bridge_s1;
  reg              last_cycle_sgdma_tx_m_read_granted_slave_cpu_ddr_clock_bridge_s1;
  wire             sgdma_rx_m_write_arbiterlock;
  wire             sgdma_rx_m_write_arbiterlock2;
  wire             sgdma_rx_m_write_continuerequest;
  wire             sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1;
  wire             sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1;
  wire             sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1;
  wire             sgdma_rx_m_write_saved_grant_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_arbiterlock;
  wire             sgdma_tx_m_read_arbiterlock2;
  wire             sgdma_tx_m_read_continuerequest;
  wire             sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  wire             sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_saved_grant_cpu_ddr_clock_bridge_s1;
  wire    [ 28: 0] shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_data_master;
  wire    [ 28: 0] shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_instruction_master;
  wire    [ 31: 0] shifted_address_to_cpu_ddr_clock_bridge_s1_from_sgdma_rx_m_write;
  wire    [ 31: 0] shifted_address_to_cpu_ddr_clock_bridge_s1_from_sgdma_tx_m_read;
  wire             wait_for_cpu_ddr_clock_bridge_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_ddr_clock_bridge_s1_end_xfer;
    end


  assign cpu_ddr_clock_bridge_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1 | cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 | sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1 | sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1));
  //assign cpu_ddr_clock_bridge_s1_readdatavalid_from_sa = cpu_ddr_clock_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_readdatavalid_from_sa = cpu_ddr_clock_bridge_s1_readdatavalid;

  //assign cpu_ddr_clock_bridge_s1_readdata_from_sa = cpu_ddr_clock_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_readdata_from_sa = cpu_ddr_clock_bridge_s1_readdata;

  assign cpu_data_master_requests_cpu_ddr_clock_bridge_s1 = ({cpu_data_master_address_to_slave[28 : 26] , 26'b0} == 29'h1c000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign cpu_ddr_clock_bridge_s1_waitrequest_from_sa = cpu_ddr_clock_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_waitrequest_from_sa = cpu_ddr_clock_bridge_s1_waitrequest;

  //cpu_ddr_clock_bridge_s1_arb_share_counter set values, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_arb_share_set_values = (cpu_data_master_granted_cpu_ddr_clock_bridge_s1)? 8 :
    (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1)? 8 :
    (cpu_data_master_granted_cpu_ddr_clock_bridge_s1)? 8 :
    (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1)? 8 :
    (cpu_data_master_granted_cpu_ddr_clock_bridge_s1)? 8 :
    (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1)? 8 :
    (cpu_data_master_granted_cpu_ddr_clock_bridge_s1)? 8 :
    (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1)? 8 :
    1;

  //cpu_ddr_clock_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_non_bursting_master_requests = cpu_data_master_requests_cpu_ddr_clock_bridge_s1 |
    cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1 |
    sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1 |
    sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1 |
    cpu_data_master_requests_cpu_ddr_clock_bridge_s1 |
    cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1 |
    sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1 |
    sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1 |
    cpu_data_master_requests_cpu_ddr_clock_bridge_s1 |
    cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1 |
    sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1 |
    sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1 |
    cpu_data_master_requests_cpu_ddr_clock_bridge_s1 |
    cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1 |
    sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1 |
    sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1;

  //cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant = 0;

  //cpu_ddr_clock_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_arb_share_counter_next_value = cpu_ddr_clock_bridge_s1_firsttransfer ? (cpu_ddr_clock_bridge_s1_arb_share_set_values - 1) : |cpu_ddr_clock_bridge_s1_arb_share_counter ? (cpu_ddr_clock_bridge_s1_arb_share_counter - 1) : 0;

  //cpu_ddr_clock_bridge_s1_allgrants all slave grants, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_allgrants = (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector) |
    (|cpu_ddr_clock_bridge_s1_grant_vector);

  //cpu_ddr_clock_bridge_s1_end_xfer assignment, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_end_xfer = ~(cpu_ddr_clock_bridge_s1_waits_for_read | cpu_ddr_clock_bridge_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 = cpu_ddr_clock_bridge_s1_end_xfer & (~cpu_ddr_clock_bridge_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_ddr_clock_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 & cpu_ddr_clock_bridge_s1_allgrants) | (end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 & ~cpu_ddr_clock_bridge_s1_non_bursting_master_requests);

  //cpu_ddr_clock_bridge_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_ddr_clock_bridge_s1_arb_share_counter <= 0;
      else if (cpu_ddr_clock_bridge_s1_arb_counter_enable)
          cpu_ddr_clock_bridge_s1_arb_share_counter <= cpu_ddr_clock_bridge_s1_arb_share_counter_next_value;
    end


  //cpu_ddr_clock_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_ddr_clock_bridge_s1_slavearbiterlockenable <= 0;
      else if ((|cpu_ddr_clock_bridge_s1_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1) | (end_xfer_arb_share_counter_term_cpu_ddr_clock_bridge_s1 & ~cpu_ddr_clock_bridge_s1_non_bursting_master_requests))
          cpu_ddr_clock_bridge_s1_slavearbiterlockenable <= |cpu_ddr_clock_bridge_s1_arb_share_counter_next_value;
    end


  //cpu/data_master cpu_ddr_clock_bridge/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = cpu_ddr_clock_bridge_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 = |cpu_ddr_clock_bridge_s1_arb_share_counter_next_value;

  //cpu/data_master cpu_ddr_clock_bridge/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master cpu_ddr_clock_bridge/s1 arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = cpu_ddr_clock_bridge_s1_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master cpu_ddr_clock_bridge/s1 arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted cpu_ddr_clock_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 <= cpu_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1 ? 1 : (cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal | ~cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1) ? 0 : last_cycle_cpu_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = (last_cycle_cpu_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 & cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1) |
    (last_cycle_cpu_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 & cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1) |
    (last_cycle_cpu_instruction_master_granted_slave_cpu_ddr_clock_bridge_s1 & cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1);

  //cpu_ddr_clock_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_any_continuerequest = cpu_instruction_master_continuerequest |
    sgdma_rx_m_write_continuerequest |
    sgdma_tx_m_read_continuerequest |
    cpu_data_master_continuerequest |
    sgdma_rx_m_write_continuerequest |
    sgdma_tx_m_read_continuerequest |
    cpu_data_master_continuerequest |
    cpu_instruction_master_continuerequest |
    sgdma_tx_m_read_continuerequest |
    cpu_data_master_continuerequest |
    cpu_instruction_master_continuerequest |
    sgdma_rx_m_write_continuerequest;

  //sgdma_rx/m_write cpu_ddr_clock_bridge/s1 arbiterlock, which is an e_assign
  assign sgdma_rx_m_write_arbiterlock = cpu_ddr_clock_bridge_s1_slavearbiterlockenable & sgdma_rx_m_write_continuerequest;

  //sgdma_rx/m_write cpu_ddr_clock_bridge/s1 arbiterlock2, which is an e_assign
  assign sgdma_rx_m_write_arbiterlock2 = cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 & sgdma_rx_m_write_continuerequest;

  //sgdma_rx/m_write granted cpu_ddr_clock_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_rx_m_write_granted_slave_cpu_ddr_clock_bridge_s1 <= 0;
      else 
        last_cycle_sgdma_rx_m_write_granted_slave_cpu_ddr_clock_bridge_s1 <= sgdma_rx_m_write_saved_grant_cpu_ddr_clock_bridge_s1 ? 1 : (cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal | ~sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1) ? 0 : last_cycle_sgdma_rx_m_write_granted_slave_cpu_ddr_clock_bridge_s1;
    end


  //sgdma_rx_m_write_continuerequest continued request, which is an e_mux
  assign sgdma_rx_m_write_continuerequest = (last_cycle_sgdma_rx_m_write_granted_slave_cpu_ddr_clock_bridge_s1 & sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1) |
    (last_cycle_sgdma_rx_m_write_granted_slave_cpu_ddr_clock_bridge_s1 & sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1) |
    (last_cycle_sgdma_rx_m_write_granted_slave_cpu_ddr_clock_bridge_s1 & sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1);

  //sgdma_tx/m_read cpu_ddr_clock_bridge/s1 arbiterlock, which is an e_assign
  assign sgdma_tx_m_read_arbiterlock = cpu_ddr_clock_bridge_s1_slavearbiterlockenable & sgdma_tx_m_read_continuerequest;

  //sgdma_tx/m_read cpu_ddr_clock_bridge/s1 arbiterlock2, which is an e_assign
  assign sgdma_tx_m_read_arbiterlock2 = cpu_ddr_clock_bridge_s1_slavearbiterlockenable2 & sgdma_tx_m_read_continuerequest;

  //sgdma_tx/m_read granted cpu_ddr_clock_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_tx_m_read_granted_slave_cpu_ddr_clock_bridge_s1 <= 0;
      else 
        last_cycle_sgdma_tx_m_read_granted_slave_cpu_ddr_clock_bridge_s1 <= sgdma_tx_m_read_saved_grant_cpu_ddr_clock_bridge_s1 ? 1 : (cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal | ~sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1) ? 0 : last_cycle_sgdma_tx_m_read_granted_slave_cpu_ddr_clock_bridge_s1;
    end


  //sgdma_tx_m_read_continuerequest continued request, which is an e_mux
  assign sgdma_tx_m_read_continuerequest = (last_cycle_sgdma_tx_m_read_granted_slave_cpu_ddr_clock_bridge_s1 & sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1) |
    (last_cycle_sgdma_tx_m_read_granted_slave_cpu_ddr_clock_bridge_s1 & sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1) |
    (last_cycle_sgdma_tx_m_read_granted_slave_cpu_ddr_clock_bridge_s1 & sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1);

  assign cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1 = cpu_data_master_requests_cpu_ddr_clock_bridge_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register))) | cpu_instruction_master_arbiterlock | sgdma_rx_m_write_arbiterlock | sgdma_tx_m_read_arbiterlock);
  //unique name for cpu_ddr_clock_bridge_s1_move_on_to_next_transaction, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_move_on_to_next_transaction = cpu_ddr_clock_bridge_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_cpu_ddr_clock_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_cpu_ddr_clock_bridge_s1_module rdv_fifo_for_cpu_data_master_to_cpu_ddr_clock_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_cpu_ddr_clock_bridge_s1),
      .data_out             (cpu_data_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1),
      .full                 (),
      .read                 (cpu_ddr_clock_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~cpu_ddr_clock_bridge_s1_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register = ~cpu_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  //local readdatavalid cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1 = (cpu_ddr_clock_bridge_s1_readdatavalid_from_sa & cpu_data_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1) & ~ cpu_data_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;

  //cpu_ddr_clock_bridge_s1_writedata mux, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_writedata = (cpu_data_master_granted_cpu_ddr_clock_bridge_s1)? cpu_data_master_writedata :
    sgdma_rx_m_write_writedata;

  //assign cpu_ddr_clock_bridge_s1_endofpacket_from_sa = cpu_ddr_clock_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_endofpacket_from_sa = cpu_ddr_clock_bridge_s1_endofpacket;

  assign cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1 = (({cpu_instruction_master_address_to_slave[28 : 26] , 26'b0} == 29'h1c000000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted cpu_ddr_clock_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_cpu_ddr_clock_bridge_s1 <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_cpu_ddr_clock_bridge_s1 <= cpu_data_master_saved_grant_cpu_ddr_clock_bridge_s1 ? 1 : (cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal | ~cpu_data_master_requests_cpu_ddr_clock_bridge_s1) ? 0 : last_cycle_cpu_data_master_granted_slave_cpu_ddr_clock_bridge_s1;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = (last_cycle_cpu_data_master_granted_slave_cpu_ddr_clock_bridge_s1 & cpu_data_master_requests_cpu_ddr_clock_bridge_s1) |
    (last_cycle_cpu_data_master_granted_slave_cpu_ddr_clock_bridge_s1 & cpu_data_master_requests_cpu_ddr_clock_bridge_s1) |
    (last_cycle_cpu_data_master_granted_slave_cpu_ddr_clock_bridge_s1 & cpu_data_master_requests_cpu_ddr_clock_bridge_s1);

  assign cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1 = cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1 & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register))) | cpu_data_master_arbiterlock | sgdma_rx_m_write_arbiterlock | sgdma_tx_m_read_arbiterlock);
  //rdv_fifo_for_cpu_instruction_master_to_cpu_ddr_clock_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_cpu_ddr_clock_bridge_s1_module rdv_fifo_for_cpu_instruction_master_to_cpu_ddr_clock_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1),
      .full                 (),
      .read                 (cpu_ddr_clock_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~cpu_ddr_clock_bridge_s1_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register = ~cpu_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  //local readdatavalid cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1, which is an e_mux
  assign cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1 = (cpu_ddr_clock_bridge_s1_readdatavalid_from_sa & cpu_instruction_master_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1) & ~ cpu_instruction_master_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;

  assign sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1 = (({sgdma_rx_m_write_address_to_slave[31 : 26] , 26'b0} == 32'h1c000000) & (sgdma_rx_m_write_write)) & sgdma_rx_m_write_write;
  assign sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1 = sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1 & ~(cpu_data_master_arbiterlock | cpu_instruction_master_arbiterlock | sgdma_tx_m_read_arbiterlock);
  assign sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1 = (({sgdma_tx_m_read_address_to_slave[31 : 26] , 26'b0} == 32'h1c000000) & (sgdma_tx_m_read_read)) & sgdma_tx_m_read_read;
  assign sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1 = sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1 & ~((sgdma_tx_m_read_read & ((sgdma_tx_m_read_latency_counter != 0) | (1 < sgdma_tx_m_read_latency_counter))) | cpu_data_master_arbiterlock | cpu_instruction_master_arbiterlock | sgdma_rx_m_write_arbiterlock);
  //rdv_fifo_for_sgdma_tx_m_read_to_cpu_ddr_clock_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_sgdma_tx_m_read_to_cpu_ddr_clock_bridge_s1_module rdv_fifo_for_sgdma_tx_m_read_to_cpu_ddr_clock_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1),
      .data_out             (sgdma_tx_m_read_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (sgdma_tx_m_read_rdv_fifo_empty_cpu_ddr_clock_bridge_s1),
      .full                 (),
      .read                 (cpu_ddr_clock_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~cpu_ddr_clock_bridge_s1_waits_for_read)
    );

  assign sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register = ~sgdma_tx_m_read_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;
  //local readdatavalid sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1, which is an e_mux
  assign sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1 = (cpu_ddr_clock_bridge_s1_readdatavalid_from_sa & sgdma_tx_m_read_rdv_fifo_output_from_cpu_ddr_clock_bridge_s1) & ~ sgdma_tx_m_read_rdv_fifo_empty_cpu_ddr_clock_bridge_s1;

  //allow new arb cycle for cpu_ddr_clock_bridge/s1, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock & ~sgdma_rx_m_write_arbiterlock & ~sgdma_tx_m_read_arbiterlock;

  //sgdma_tx/m_read assignment into master qualified-requests vector for cpu_ddr_clock_bridge/s1, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_master_qreq_vector[0] = sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1;

  //sgdma_tx/m_read grant cpu_ddr_clock_bridge/s1, which is an e_assign
  assign sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1 = cpu_ddr_clock_bridge_s1_grant_vector[0];

  //sgdma_tx/m_read saved-grant cpu_ddr_clock_bridge/s1, which is an e_assign
  assign sgdma_tx_m_read_saved_grant_cpu_ddr_clock_bridge_s1 = cpu_ddr_clock_bridge_s1_arb_winner[0] && sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1;

  //sgdma_rx/m_write assignment into master qualified-requests vector for cpu_ddr_clock_bridge/s1, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_master_qreq_vector[1] = sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1;

  //sgdma_rx/m_write grant cpu_ddr_clock_bridge/s1, which is an e_assign
  assign sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1 = cpu_ddr_clock_bridge_s1_grant_vector[1];

  //sgdma_rx/m_write saved-grant cpu_ddr_clock_bridge/s1, which is an e_assign
  assign sgdma_rx_m_write_saved_grant_cpu_ddr_clock_bridge_s1 = cpu_ddr_clock_bridge_s1_arb_winner[1] && sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1;

  //cpu/instruction_master assignment into master qualified-requests vector for cpu_ddr_clock_bridge/s1, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_master_qreq_vector[2] = cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1;

  //cpu/instruction_master grant cpu_ddr_clock_bridge/s1, which is an e_assign
  assign cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1 = cpu_ddr_clock_bridge_s1_grant_vector[2];

  //cpu/instruction_master saved-grant cpu_ddr_clock_bridge/s1, which is an e_assign
  assign cpu_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1 = cpu_ddr_clock_bridge_s1_arb_winner[2] && cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1;

  //cpu/data_master assignment into master qualified-requests vector for cpu_ddr_clock_bridge/s1, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_master_qreq_vector[3] = cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1;

  //cpu/data_master grant cpu_ddr_clock_bridge/s1, which is an e_assign
  assign cpu_data_master_granted_cpu_ddr_clock_bridge_s1 = cpu_ddr_clock_bridge_s1_grant_vector[3];

  //cpu/data_master saved-grant cpu_ddr_clock_bridge/s1, which is an e_assign
  assign cpu_data_master_saved_grant_cpu_ddr_clock_bridge_s1 = cpu_ddr_clock_bridge_s1_arb_winner[3] && cpu_data_master_requests_cpu_ddr_clock_bridge_s1;

  //cpu_ddr_clock_bridge/s1 chosen-master double-vector, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_chosen_master_double_vector = {cpu_ddr_clock_bridge_s1_master_qreq_vector, cpu_ddr_clock_bridge_s1_master_qreq_vector} & ({~cpu_ddr_clock_bridge_s1_master_qreq_vector, ~cpu_ddr_clock_bridge_s1_master_qreq_vector} + cpu_ddr_clock_bridge_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_ddr_clock_bridge_s1_arb_winner = (cpu_ddr_clock_bridge_s1_allow_new_arb_cycle & | cpu_ddr_clock_bridge_s1_grant_vector) ? cpu_ddr_clock_bridge_s1_grant_vector : cpu_ddr_clock_bridge_s1_saved_chosen_master_vector;

  //saved cpu_ddr_clock_bridge_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_ddr_clock_bridge_s1_saved_chosen_master_vector <= 0;
      else if (cpu_ddr_clock_bridge_s1_allow_new_arb_cycle)
          cpu_ddr_clock_bridge_s1_saved_chosen_master_vector <= |cpu_ddr_clock_bridge_s1_grant_vector ? cpu_ddr_clock_bridge_s1_grant_vector : cpu_ddr_clock_bridge_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_ddr_clock_bridge_s1_grant_vector = {(cpu_ddr_clock_bridge_s1_chosen_master_double_vector[3] | cpu_ddr_clock_bridge_s1_chosen_master_double_vector[7]),
    (cpu_ddr_clock_bridge_s1_chosen_master_double_vector[2] | cpu_ddr_clock_bridge_s1_chosen_master_double_vector[6]),
    (cpu_ddr_clock_bridge_s1_chosen_master_double_vector[1] | cpu_ddr_clock_bridge_s1_chosen_master_double_vector[5]),
    (cpu_ddr_clock_bridge_s1_chosen_master_double_vector[0] | cpu_ddr_clock_bridge_s1_chosen_master_double_vector[4])};

  //cpu_ddr_clock_bridge/s1 chosen master rotated left, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_chosen_master_rot_left = (cpu_ddr_clock_bridge_s1_arb_winner << 1) ? (cpu_ddr_clock_bridge_s1_arb_winner << 1) : 1;

  //cpu_ddr_clock_bridge/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_ddr_clock_bridge_s1_arb_addend <= 1;
      else if (|cpu_ddr_clock_bridge_s1_grant_vector)
          cpu_ddr_clock_bridge_s1_arb_addend <= cpu_ddr_clock_bridge_s1_end_xfer? cpu_ddr_clock_bridge_s1_chosen_master_rot_left : cpu_ddr_clock_bridge_s1_grant_vector;
    end


  //cpu_ddr_clock_bridge_s1_reset_n assignment, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_reset_n = reset_n;

  //cpu_ddr_clock_bridge_s1_firsttransfer first transaction, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_firsttransfer = cpu_ddr_clock_bridge_s1_begins_xfer ? cpu_ddr_clock_bridge_s1_unreg_firsttransfer : cpu_ddr_clock_bridge_s1_reg_firsttransfer;

  //cpu_ddr_clock_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_unreg_firsttransfer = ~(cpu_ddr_clock_bridge_s1_slavearbiterlockenable & cpu_ddr_clock_bridge_s1_any_continuerequest);

  //cpu_ddr_clock_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_ddr_clock_bridge_s1_reg_firsttransfer <= 1'b1;
      else if (cpu_ddr_clock_bridge_s1_begins_xfer)
          cpu_ddr_clock_bridge_s1_reg_firsttransfer <= cpu_ddr_clock_bridge_s1_unreg_firsttransfer;
    end


  //cpu_ddr_clock_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_beginbursttransfer_internal = cpu_ddr_clock_bridge_s1_begins_xfer;

  //cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_arbitration_holdoff_internal = cpu_ddr_clock_bridge_s1_begins_xfer & cpu_ddr_clock_bridge_s1_firsttransfer;

  //cpu_ddr_clock_bridge_s1_read assignment, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_read = (cpu_data_master_granted_cpu_ddr_clock_bridge_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1 & cpu_instruction_master_read) | (sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1 & sgdma_tx_m_read_read);

  //cpu_ddr_clock_bridge_s1_write assignment, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_write = (cpu_data_master_granted_cpu_ddr_clock_bridge_s1 & cpu_data_master_write) | (sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1 & sgdma_rx_m_write_write);

  assign shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //cpu_ddr_clock_bridge_s1_address mux, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_address = (cpu_data_master_granted_cpu_ddr_clock_bridge_s1)? (shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_data_master >> 2) :
    (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1)? (shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_instruction_master >> 2) :
    (sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1)? (shifted_address_to_cpu_ddr_clock_bridge_s1_from_sgdma_rx_m_write >> 2) :
    (shifted_address_to_cpu_ddr_clock_bridge_s1_from_sgdma_tx_m_read >> 2);

  assign shifted_address_to_cpu_ddr_clock_bridge_s1_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  assign shifted_address_to_cpu_ddr_clock_bridge_s1_from_sgdma_rx_m_write = sgdma_rx_m_write_address_to_slave;
  assign shifted_address_to_cpu_ddr_clock_bridge_s1_from_sgdma_tx_m_read = sgdma_tx_m_read_address_to_slave;
  //slaveid cpu_ddr_clock_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_nativeaddress = (cpu_data_master_granted_cpu_ddr_clock_bridge_s1)? (cpu_data_master_address_to_slave >> 2) :
    (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1)? (cpu_instruction_master_address_to_slave >> 2) :
    (sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1)? (sgdma_rx_m_write_address_to_slave >> 2) :
    (sgdma_tx_m_read_address_to_slave >> 2);

  //d1_cpu_ddr_clock_bridge_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_ddr_clock_bridge_s1_end_xfer <= 1;
      else 
        d1_cpu_ddr_clock_bridge_s1_end_xfer <= cpu_ddr_clock_bridge_s1_end_xfer;
    end


  //cpu_ddr_clock_bridge_s1_waits_for_read in a cycle, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_waits_for_read = cpu_ddr_clock_bridge_s1_in_a_read_cycle & cpu_ddr_clock_bridge_s1_waitrequest_from_sa;

  //cpu_ddr_clock_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_in_a_read_cycle = (cpu_data_master_granted_cpu_ddr_clock_bridge_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1 & cpu_instruction_master_read) | (sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1 & sgdma_tx_m_read_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_ddr_clock_bridge_s1_in_a_read_cycle;

  //cpu_ddr_clock_bridge_s1_waits_for_write in a cycle, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_waits_for_write = cpu_ddr_clock_bridge_s1_in_a_write_cycle & cpu_ddr_clock_bridge_s1_waitrequest_from_sa;

  //cpu_ddr_clock_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  assign cpu_ddr_clock_bridge_s1_in_a_write_cycle = (cpu_data_master_granted_cpu_ddr_clock_bridge_s1 & cpu_data_master_write) | (sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1 & sgdma_rx_m_write_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_ddr_clock_bridge_s1_in_a_write_cycle;

  assign wait_for_cpu_ddr_clock_bridge_s1_counter = 0;
  //cpu_ddr_clock_bridge_s1_byteenable byte enable port mux, which is an e_mux
  assign cpu_ddr_clock_bridge_s1_byteenable = (cpu_data_master_granted_cpu_ddr_clock_bridge_s1)? cpu_data_master_byteenable :
    (sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1)? sgdma_rx_m_write_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_ddr_clock_bridge/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_cpu_ddr_clock_bridge_s1 + cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1 + sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1 + sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_cpu_ddr_clock_bridge_s1 + cpu_instruction_master_saved_grant_cpu_ddr_clock_bridge_s1 + sgdma_rx_m_write_saved_grant_cpu_ddr_clock_bridge_s1 + sgdma_tx_m_read_saved_grant_cpu_ddr_clock_bridge_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_ddr_clock_bridge_m1_arbitrator (
                                            // inputs:
                                             clk,
                                             cpu_ddr_clock_bridge_m1_address,
                                             cpu_ddr_clock_bridge_m1_byteenable,
                                             cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1,
                                             cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1,
                                             cpu_ddr_clock_bridge_m1_read,
                                             cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1,
                                             cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register,
                                             cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1,
                                             cpu_ddr_clock_bridge_m1_write,
                                             cpu_ddr_clock_bridge_m1_writedata,
                                             d1_ddr2_sdram_s1_end_xfer,
                                             ddr2_sdram_s1_readdata_from_sa,
                                             ddr2_sdram_s1_waitrequest_n_from_sa,
                                             reset_n,

                                            // outputs:
                                             cpu_ddr_clock_bridge_m1_address_to_slave,
                                             cpu_ddr_clock_bridge_m1_latency_counter,
                                             cpu_ddr_clock_bridge_m1_readdata,
                                             cpu_ddr_clock_bridge_m1_readdatavalid,
                                             cpu_ddr_clock_bridge_m1_reset_n,
                                             cpu_ddr_clock_bridge_m1_waitrequest
                                          )
;

  output  [ 25: 0] cpu_ddr_clock_bridge_m1_address_to_slave;
  output           cpu_ddr_clock_bridge_m1_latency_counter;
  output  [ 31: 0] cpu_ddr_clock_bridge_m1_readdata;
  output           cpu_ddr_clock_bridge_m1_readdatavalid;
  output           cpu_ddr_clock_bridge_m1_reset_n;
  output           cpu_ddr_clock_bridge_m1_waitrequest;
  input            clk;
  input   [ 25: 0] cpu_ddr_clock_bridge_m1_address;
  input   [  3: 0] cpu_ddr_clock_bridge_m1_byteenable;
  input            cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1;
  input            cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1;
  input            cpu_ddr_clock_bridge_m1_read;
  input            cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1;
  input            cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register;
  input            cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1;
  input            cpu_ddr_clock_bridge_m1_write;
  input   [ 31: 0] cpu_ddr_clock_bridge_m1_writedata;
  input            d1_ddr2_sdram_s1_end_xfer;
  input   [ 31: 0] ddr2_sdram_s1_readdata_from_sa;
  input            ddr2_sdram_s1_waitrequest_n_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 25: 0] cpu_ddr_clock_bridge_m1_address_last_time;
  wire    [ 25: 0] cpu_ddr_clock_bridge_m1_address_to_slave;
  reg     [  3: 0] cpu_ddr_clock_bridge_m1_byteenable_last_time;
  wire             cpu_ddr_clock_bridge_m1_latency_counter;
  reg              cpu_ddr_clock_bridge_m1_read_last_time;
  wire    [ 31: 0] cpu_ddr_clock_bridge_m1_readdata;
  wire             cpu_ddr_clock_bridge_m1_readdatavalid;
  wire             cpu_ddr_clock_bridge_m1_reset_n;
  wire             cpu_ddr_clock_bridge_m1_run;
  wire             cpu_ddr_clock_bridge_m1_waitrequest;
  reg              cpu_ddr_clock_bridge_m1_write_last_time;
  reg     [ 31: 0] cpu_ddr_clock_bridge_m1_writedata_last_time;
  wire             pre_flush_cpu_ddr_clock_bridge_m1_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1 | ~cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1) & ((~cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1 | ~(cpu_ddr_clock_bridge_m1_read | cpu_ddr_clock_bridge_m1_write) | (1 & ddr2_sdram_s1_waitrequest_n_from_sa & (cpu_ddr_clock_bridge_m1_read | cpu_ddr_clock_bridge_m1_write)))) & ((~cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1 | ~(cpu_ddr_clock_bridge_m1_read | cpu_ddr_clock_bridge_m1_write) | (1 & ddr2_sdram_s1_waitrequest_n_from_sa & (cpu_ddr_clock_bridge_m1_read | cpu_ddr_clock_bridge_m1_write))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_ddr_clock_bridge_m1_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_ddr_clock_bridge_m1_address_to_slave = cpu_ddr_clock_bridge_m1_address[25 : 0];

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_ddr_clock_bridge_m1_readdatavalid = cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_ddr_clock_bridge_m1_readdatavalid = 0 |
    pre_flush_cpu_ddr_clock_bridge_m1_readdatavalid;

  //cpu_ddr_clock_bridge/m1 readdata mux, which is an e_mux
  assign cpu_ddr_clock_bridge_m1_readdata = ddr2_sdram_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign cpu_ddr_clock_bridge_m1_waitrequest = ~cpu_ddr_clock_bridge_m1_run;

  //latent max counter, which is an e_assign
  assign cpu_ddr_clock_bridge_m1_latency_counter = 0;

  //cpu_ddr_clock_bridge_m1_reset_n assignment, which is an e_assign
  assign cpu_ddr_clock_bridge_m1_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_ddr_clock_bridge_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_ddr_clock_bridge_m1_address_last_time <= 0;
      else 
        cpu_ddr_clock_bridge_m1_address_last_time <= cpu_ddr_clock_bridge_m1_address;
    end


  //cpu_ddr_clock_bridge/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_ddr_clock_bridge_m1_waitrequest & (cpu_ddr_clock_bridge_m1_read | cpu_ddr_clock_bridge_m1_write);
    end


  //cpu_ddr_clock_bridge_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_ddr_clock_bridge_m1_address != cpu_ddr_clock_bridge_m1_address_last_time))
        begin
          $write("%0d ns: cpu_ddr_clock_bridge_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_ddr_clock_bridge_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_ddr_clock_bridge_m1_byteenable_last_time <= 0;
      else 
        cpu_ddr_clock_bridge_m1_byteenable_last_time <= cpu_ddr_clock_bridge_m1_byteenable;
    end


  //cpu_ddr_clock_bridge_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_ddr_clock_bridge_m1_byteenable != cpu_ddr_clock_bridge_m1_byteenable_last_time))
        begin
          $write("%0d ns: cpu_ddr_clock_bridge_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_ddr_clock_bridge_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_ddr_clock_bridge_m1_read_last_time <= 0;
      else 
        cpu_ddr_clock_bridge_m1_read_last_time <= cpu_ddr_clock_bridge_m1_read;
    end


  //cpu_ddr_clock_bridge_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_ddr_clock_bridge_m1_read != cpu_ddr_clock_bridge_m1_read_last_time))
        begin
          $write("%0d ns: cpu_ddr_clock_bridge_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_ddr_clock_bridge_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_ddr_clock_bridge_m1_write_last_time <= 0;
      else 
        cpu_ddr_clock_bridge_m1_write_last_time <= cpu_ddr_clock_bridge_m1_write;
    end


  //cpu_ddr_clock_bridge_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_ddr_clock_bridge_m1_write != cpu_ddr_clock_bridge_m1_write_last_time))
        begin
          $write("%0d ns: cpu_ddr_clock_bridge_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_ddr_clock_bridge_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_ddr_clock_bridge_m1_writedata_last_time <= 0;
      else 
        cpu_ddr_clock_bridge_m1_writedata_last_time <= cpu_ddr_clock_bridge_m1_writedata;
    end


  //cpu_ddr_clock_bridge_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_ddr_clock_bridge_m1_writedata != cpu_ddr_clock_bridge_m1_writedata_last_time) & cpu_ddr_clock_bridge_m1_write)
        begin
          $write("%0d ns: cpu_ddr_clock_bridge_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_ddr_clock_bridge_bridge_arbitrator 
;



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arbitrator (
                                                                     // inputs:
                                                                      clk,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest,
                                                                      reset_n,
                                                                      slow_peripheral_bridge_m1_address_to_slave,
                                                                      slow_peripheral_bridge_m1_byteenable,
                                                                      slow_peripheral_bridge_m1_latency_counter,
                                                                      slow_peripheral_bridge_m1_nativeaddress,
                                                                      slow_peripheral_bridge_m1_read,
                                                                      slow_peripheral_bridge_m1_write,
                                                                      slow_peripheral_bridge_m1_writedata,

                                                                     // outputs:
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_address,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_byteenable,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_nativeaddress,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_read,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reset_n,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_write,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_0_in_writedata,
                                                                      d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer,
                                                                      slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in,
                                                                      slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in,
                                                                      slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in,
                                                                      slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in
                                                                   )
;

  output  [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_address;
  output  [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_byteenable;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa;
  output  [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_nativeaddress;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_in_read;
  output  [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reset_n;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_in_write;
  output  [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_writedata;
  output           d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer;
  output           slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  output           slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  output           slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  output           slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  input            clk;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  input   [  3: 0] slow_peripheral_bridge_m1_byteenable;
  input            slow_peripheral_bridge_m1_latency_counter;
  input   [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] slow_peripheral_bridge_m1_writedata;

  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_address;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_allgrants;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_allow_new_arb_cycle;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_any_bursting_master_saved_grant;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_any_continuerequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_counter_enable;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter_next_value;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_set_values;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_beginbursttransfer_internal;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_begins_xfer;
  wire    [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_byteenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_firsttransfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_grant_vector;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_in_a_read_cycle;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_in_a_write_cycle;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_master_qreq_vector;
  wire    [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_nativeaddress;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_non_bursting_master_requests;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_read;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reg_firsttransfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reset_n;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_0_in_slavearbiterlockenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_slavearbiterlockenable2;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_unreg_firsttransfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waits_for_read;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waits_for_write;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_write;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_writedata;
  reg              d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             slow_peripheral_bridge_m1_arbiterlock;
  wire             slow_peripheral_bridge_m1_arbiterlock2;
  wire             slow_peripheral_bridge_m1_continuerequest;
  wire             slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  wire             slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  wire             slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  wire             slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  wire             slow_peripheral_bridge_m1_saved_grant_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  wire             wait_for_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer;
    end


  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_begins_xfer = ~d1_reasons_to_wait & ((slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in));
  //assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata;

  assign slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in = ({slow_peripheral_bridge_m1_address_to_slave[7 : 5] , 5'b0} == 8'h40) & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write);
  //assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter set values, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_set_values = 1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_non_bursting_master_requests = slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_any_bursting_master_saved_grant = 0;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter_next_value = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_firsttransfer ? (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_set_values - 1) : |cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter ? (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter - 1) : 0;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_allgrants all slave grants, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_allgrants = |cycloneIII_3c120_niosII_standard_sopc_clock_0_in_grant_vector;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer = ~(cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waits_for_read | cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waits_for_write);

  //end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_0_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_0_in = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer & (~cycloneIII_3c120_niosII_standard_sopc_clock_0_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_counter_enable = (end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_0_in & cycloneIII_3c120_niosII_standard_sopc_clock_0_in_allgrants) | (end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_0_in & ~cycloneIII_3c120_niosII_standard_sopc_clock_0_in_non_bursting_master_requests);

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter <= 0;
      else if (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_counter_enable)
          cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter <= cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter_next_value;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_0_in_slavearbiterlockenable <= 0;
      else if ((|cycloneIII_3c120_niosII_standard_sopc_clock_0_in_master_qreq_vector & end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_0_in) | (end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_0_in & ~cycloneIII_3c120_niosII_standard_sopc_clock_0_in_non_bursting_master_requests))
          cycloneIII_3c120_niosII_standard_sopc_clock_0_in_slavearbiterlockenable <= |cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge/m1 cycloneIII_3c120_niosII_standard_sopc_clock_0/in arbiterlock, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_slavearbiterlockenable & slow_peripheral_bridge_m1_continuerequest;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_slavearbiterlockenable2 = |cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arb_share_counter_next_value;

  //slow_peripheral_bridge/m1 cycloneIII_3c120_niosII_standard_sopc_clock_0/in arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock2 = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_slavearbiterlockenable2 & slow_peripheral_bridge_m1_continuerequest;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_any_continuerequest = 1;

  //slow_peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  assign slow_peripheral_bridge_m1_continuerequest = 1;

  assign slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in = slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in & ~((slow_peripheral_bridge_m1_read & ((slow_peripheral_bridge_m1_latency_counter != 0))));
  //local readdatavalid slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in & slow_peripheral_bridge_m1_read & ~cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waits_for_read;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_writedata mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_writedata = slow_peripheral_bridge_m1_writedata;

  //assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket;

  //master is always granted when requested
  assign slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in = slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;

  //slow_peripheral_bridge/m1 saved-grant cycloneIII_3c120_niosII_standard_sopc_clock_0/in, which is an e_assign
  assign slow_peripheral_bridge_m1_saved_grant_cycloneIII_3c120_niosII_standard_sopc_clock_0_in = slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;

  //allow new arb cycle for cycloneIII_3c120_niosII_standard_sopc_clock_0/in, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_master_qreq_vector = 1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reset_n assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reset_n = reset_n;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_firsttransfer first transaction, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_firsttransfer = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_begins_xfer ? cycloneIII_3c120_niosII_standard_sopc_clock_0_in_unreg_firsttransfer : cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reg_firsttransfer;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_unreg_firsttransfer = ~(cycloneIII_3c120_niosII_standard_sopc_clock_0_in_slavearbiterlockenable & cycloneIII_3c120_niosII_standard_sopc_clock_0_in_any_continuerequest);

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reg_firsttransfer <= 1'b1;
      else if (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_begins_xfer)
          cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reg_firsttransfer <= cycloneIII_3c120_niosII_standard_sopc_clock_0_in_unreg_firsttransfer;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_beginbursttransfer_internal = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_begins_xfer;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_read assignment, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_read = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in & slow_peripheral_bridge_m1_read;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_write assignment, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_write = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in & slow_peripheral_bridge_m1_write;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_address mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_address = slow_peripheral_bridge_m1_address_to_slave;

  //slaveid cycloneIII_3c120_niosII_standard_sopc_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_nativeaddress = slow_peripheral_bridge_m1_nativeaddress;

  //d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer <= 1;
      else 
        d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer <= cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waits_for_read in a cycle, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waits_for_read = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_in_a_read_cycle & cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_in_a_read_cycle = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in & slow_peripheral_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_in_a_read_cycle;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waits_for_write in a cycle, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waits_for_write = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_in_a_write_cycle & cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_in_a_write_cycle = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in & slow_peripheral_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_0_in_in_a_write_cycle;

  assign wait_for_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_counter = 0;
  //cycloneIII_3c120_niosII_standard_sopc_clock_0_in_byteenable byte enable port mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_in_byteenable = (slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in)? slow_peripheral_bridge_m1_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cycloneIII_3c120_niosII_standard_sopc_clock_0/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_clock_0_out_arbitrator (
                                                                      // inputs:
                                                                       clk,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_data_valid_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata,
                                                                       d1_pll_s1_end_xfer,
                                                                       pll_s1_readdata_from_sa,
                                                                       reset_n,

                                                                      // outputs:
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_readdata,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_reset_n,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_0_out_waitrequest
                                                                    )
;

  output  [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave;
  output  [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_readdata;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_out_reset_n;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_out_waitrequest;
  input            clk;
  input   [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address;
  input   [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_data_valid_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata;
  input            d1_pll_s1_end_xfer;
  input   [ 15: 0] pll_s1_readdata_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_last_time;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave;
  reg     [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable_last_time;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_last_time;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_readdata;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_reset_n;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_run;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_waitrequest;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write_last_time;
  reg     [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata_last_time;
  wire             r_1;
  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & ((~cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1 | ~cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read | (1 & ~d1_pll_s1_end_xfer & cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read))) & ((~cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1 | ~cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write | (1 & cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write)));

  //cascaded wait assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_run = r_1;

  //optimize select-logic by passing only those address bits which matter.
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0/out readdata mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_readdata = pll_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_waitrequest = ~cycloneIII_3c120_niosII_standard_sopc_clock_0_out_run;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_reset_n assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_0_out_waitrequest & (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read | cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write);
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address != cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable != cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read != cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write != cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata != cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata_last_time) & cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write)
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arbitrator (
                                                                     // inputs:
                                                                      clk,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest,
                                                                      reset_n,
                                                                      slow_peripheral_bridge_m1_address_to_slave,
                                                                      slow_peripheral_bridge_m1_byteenable,
                                                                      slow_peripheral_bridge_m1_latency_counter,
                                                                      slow_peripheral_bridge_m1_nativeaddress,
                                                                      slow_peripheral_bridge_m1_read,
                                                                      slow_peripheral_bridge_m1_write,
                                                                      slow_peripheral_bridge_m1_writedata,

                                                                     // outputs:
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_address,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_byteenable,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_nativeaddress,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_read,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reset_n,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_write,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_1_in_writedata,
                                                                      d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer,
                                                                      slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in,
                                                                      slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in,
                                                                      slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in,
                                                                      slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in
                                                                   )
;

  output  [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_address;
  output  [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_byteenable;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa;
  output  [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_nativeaddress;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_in_read;
  output  [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reset_n;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_in_write;
  output  [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_writedata;
  output           d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer;
  output           slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  output           slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  output           slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  output           slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  input            clk;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  input   [  3: 0] slow_peripheral_bridge_m1_byteenable;
  input            slow_peripheral_bridge_m1_latency_counter;
  input   [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] slow_peripheral_bridge_m1_writedata;

  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_address;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_allgrants;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_allow_new_arb_cycle;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_any_bursting_master_saved_grant;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_any_continuerequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_counter_enable;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter_next_value;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_set_values;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_beginbursttransfer_internal;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_begins_xfer;
  wire    [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_byteenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_firsttransfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_grant_vector;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_in_a_read_cycle;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_in_a_write_cycle;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_master_qreq_vector;
  wire    [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_nativeaddress;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_non_bursting_master_requests;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_read;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reg_firsttransfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reset_n;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_1_in_slavearbiterlockenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_slavearbiterlockenable2;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_unreg_firsttransfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waits_for_read;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waits_for_write;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_write;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_writedata;
  reg              d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             slow_peripheral_bridge_m1_arbiterlock;
  wire             slow_peripheral_bridge_m1_arbiterlock2;
  wire             slow_peripheral_bridge_m1_continuerequest;
  wire             slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  wire             slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  wire             slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  wire             slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  wire             slow_peripheral_bridge_m1_saved_grant_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  wire             wait_for_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer;
    end


  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_begins_xfer = ~d1_reasons_to_wait & ((slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in));
  //assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata;

  assign slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in = ({slow_peripheral_bridge_m1_address_to_slave[7 : 5] , 5'b0} == 8'h80) & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write);
  //assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter set values, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_set_values = 1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_non_bursting_master_requests mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_non_bursting_master_requests = slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_any_bursting_master_saved_grant = 0;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter_next_value assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter_next_value = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_firsttransfer ? (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_set_values - 1) : |cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter ? (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter - 1) : 0;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_allgrants all slave grants, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_allgrants = |cycloneIII_3c120_niosII_standard_sopc_clock_1_in_grant_vector;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer = ~(cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waits_for_read | cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waits_for_write);

  //end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_1_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_1_in = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer & (~cycloneIII_3c120_niosII_standard_sopc_clock_1_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_counter_enable = (end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_1_in & cycloneIII_3c120_niosII_standard_sopc_clock_1_in_allgrants) | (end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_1_in & ~cycloneIII_3c120_niosII_standard_sopc_clock_1_in_non_bursting_master_requests);

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter <= 0;
      else if (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_counter_enable)
          cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter <= cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter_next_value;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_1_in_slavearbiterlockenable <= 0;
      else if ((|cycloneIII_3c120_niosII_standard_sopc_clock_1_in_master_qreq_vector & end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_1_in) | (end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_1_in & ~cycloneIII_3c120_niosII_standard_sopc_clock_1_in_non_bursting_master_requests))
          cycloneIII_3c120_niosII_standard_sopc_clock_1_in_slavearbiterlockenable <= |cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge/m1 cycloneIII_3c120_niosII_standard_sopc_clock_1/in arbiterlock, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_slavearbiterlockenable & slow_peripheral_bridge_m1_continuerequest;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_slavearbiterlockenable2 = |cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arb_share_counter_next_value;

  //slow_peripheral_bridge/m1 cycloneIII_3c120_niosII_standard_sopc_clock_1/in arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock2 = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_slavearbiterlockenable2 & slow_peripheral_bridge_m1_continuerequest;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_any_continuerequest = 1;

  //slow_peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  assign slow_peripheral_bridge_m1_continuerequest = 1;

  assign slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in = slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in & ~((slow_peripheral_bridge_m1_read & ((slow_peripheral_bridge_m1_latency_counter != 0))));
  //local readdatavalid slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in & slow_peripheral_bridge_m1_read & ~cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waits_for_read;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_writedata mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_writedata = slow_peripheral_bridge_m1_writedata;

  //assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket;

  //master is always granted when requested
  assign slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in = slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;

  //slow_peripheral_bridge/m1 saved-grant cycloneIII_3c120_niosII_standard_sopc_clock_1/in, which is an e_assign
  assign slow_peripheral_bridge_m1_saved_grant_cycloneIII_3c120_niosII_standard_sopc_clock_1_in = slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;

  //allow new arb cycle for cycloneIII_3c120_niosII_standard_sopc_clock_1/in, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_master_qreq_vector = 1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reset_n assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reset_n = reset_n;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_firsttransfer first transaction, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_firsttransfer = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_begins_xfer ? cycloneIII_3c120_niosII_standard_sopc_clock_1_in_unreg_firsttransfer : cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reg_firsttransfer;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_unreg_firsttransfer first transaction, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_unreg_firsttransfer = ~(cycloneIII_3c120_niosII_standard_sopc_clock_1_in_slavearbiterlockenable & cycloneIII_3c120_niosII_standard_sopc_clock_1_in_any_continuerequest);

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reg_firsttransfer <= 1'b1;
      else if (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_begins_xfer)
          cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reg_firsttransfer <= cycloneIII_3c120_niosII_standard_sopc_clock_1_in_unreg_firsttransfer;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_beginbursttransfer_internal = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_begins_xfer;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_read assignment, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_read = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in & slow_peripheral_bridge_m1_read;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_write assignment, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_write = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in & slow_peripheral_bridge_m1_write;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_address mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_address = slow_peripheral_bridge_m1_address_to_slave;

  //slaveid cycloneIII_3c120_niosII_standard_sopc_clock_1_in_nativeaddress nativeaddress mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_nativeaddress = slow_peripheral_bridge_m1_nativeaddress;

  //d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer <= 1;
      else 
        d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer <= cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waits_for_read in a cycle, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waits_for_read = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_in_a_read_cycle & cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_in_a_read_cycle assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_in_a_read_cycle = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in & slow_peripheral_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_in_a_read_cycle;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waits_for_write in a cycle, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waits_for_write = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_in_a_write_cycle & cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_in_a_write_cycle assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_in_a_write_cycle = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in & slow_peripheral_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_1_in_in_a_write_cycle;

  assign wait_for_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_counter = 0;
  //cycloneIII_3c120_niosII_standard_sopc_clock_1_in_byteenable byte enable port mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_in_byteenable = (slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in)? slow_peripheral_bridge_m1_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cycloneIII_3c120_niosII_standard_sopc_clock_1/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_clock_1_out_arbitrator (
                                                                      // inputs:
                                                                       clk,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_data_valid_tse_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata,
                                                                       d1_tse_pll_s1_end_xfer,
                                                                       reset_n,
                                                                       tse_pll_s1_readdata_from_sa,

                                                                      // outputs:
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_readdata,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_reset_n,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_1_out_waitrequest
                                                                    )
;

  output  [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave;
  output  [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_readdata;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_out_reset_n;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_out_waitrequest;
  input            clk;
  input   [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address;
  input   [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_data_valid_tse_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata;
  input            d1_tse_pll_s1_end_xfer;
  input            reset_n;
  input   [ 15: 0] tse_pll_s1_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_last_time;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave;
  reg     [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable_last_time;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_last_time;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_readdata;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_reset_n;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_run;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_waitrequest;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write_last_time;
  reg     [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata_last_time;
  wire             r_2;
  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & ((~cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1 | ~cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read | (1 & ~d1_tse_pll_s1_end_xfer & cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read))) & ((~cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1 | ~cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write | (1 & cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write)));

  //cascaded wait assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_run = r_2;

  //optimize select-logic by passing only those address bits which matter.
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1/out readdata mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_readdata = tse_pll_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_waitrequest = ~cycloneIII_3c120_niosII_standard_sopc_clock_1_out_run;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_reset_n assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_1_out_waitrequest & (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read | cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write);
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address != cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable != cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read != cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write != cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata != cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata_last_time) & cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write)
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arbitrator (
                                                                     // inputs:
                                                                      clk,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest,
                                                                      reset_n,
                                                                      slow_peripheral_bridge_m1_address_to_slave,
                                                                      slow_peripheral_bridge_m1_byteenable,
                                                                      slow_peripheral_bridge_m1_latency_counter,
                                                                      slow_peripheral_bridge_m1_nativeaddress,
                                                                      slow_peripheral_bridge_m1_read,
                                                                      slow_peripheral_bridge_m1_write,
                                                                      slow_peripheral_bridge_m1_writedata,

                                                                     // outputs:
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_address,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_byteenable,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_nativeaddress,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_read,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reset_n,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_write,
                                                                      cycloneIII_3c120_niosII_standard_sopc_clock_2_in_writedata,
                                                                      d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer,
                                                                      slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in,
                                                                      slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in,
                                                                      slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in,
                                                                      slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in
                                                                   )
;

  output  [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_address;
  output  [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_byteenable;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa;
  output  [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_nativeaddress;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_in_read;
  output  [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reset_n;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_in_write;
  output  [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_writedata;
  output           d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer;
  output           slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  output           slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  output           slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  output           slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  input            clk;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  input   [  3: 0] slow_peripheral_bridge_m1_byteenable;
  input            slow_peripheral_bridge_m1_latency_counter;
  input   [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] slow_peripheral_bridge_m1_writedata;

  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_address;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_allgrants;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_allow_new_arb_cycle;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_any_bursting_master_saved_grant;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_any_continuerequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_counter_enable;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter_next_value;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_set_values;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_beginbursttransfer_internal;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_begins_xfer;
  wire    [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_byteenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_firsttransfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_grant_vector;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_in_a_read_cycle;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_in_a_write_cycle;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_master_qreq_vector;
  wire    [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_nativeaddress;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_non_bursting_master_requests;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_read;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reg_firsttransfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reset_n;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_2_in_slavearbiterlockenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_slavearbiterlockenable2;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_unreg_firsttransfer;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waits_for_read;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waits_for_write;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_write;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_writedata;
  reg              d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             slow_peripheral_bridge_m1_arbiterlock;
  wire             slow_peripheral_bridge_m1_arbiterlock2;
  wire             slow_peripheral_bridge_m1_continuerequest;
  wire             slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  wire             slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  wire             slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  wire             slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  wire             slow_peripheral_bridge_m1_saved_grant_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  wire             wait_for_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer;
    end


  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_begins_xfer = ~d1_reasons_to_wait & ((slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in));
  //assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata;

  assign slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in = ({slow_peripheral_bridge_m1_address_to_slave[7 : 5] , 5'b0} == 8'h60) & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write);
  //assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter set values, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_set_values = 1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_non_bursting_master_requests mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_non_bursting_master_requests = slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_any_bursting_master_saved_grant = 0;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter_next_value assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter_next_value = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_firsttransfer ? (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_set_values - 1) : |cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter ? (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter - 1) : 0;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_allgrants all slave grants, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_allgrants = |cycloneIII_3c120_niosII_standard_sopc_clock_2_in_grant_vector;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer = ~(cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waits_for_read | cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waits_for_write);

  //end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_2_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_2_in = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer & (~cycloneIII_3c120_niosII_standard_sopc_clock_2_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_counter_enable = (end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_2_in & cycloneIII_3c120_niosII_standard_sopc_clock_2_in_allgrants) | (end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_2_in & ~cycloneIII_3c120_niosII_standard_sopc_clock_2_in_non_bursting_master_requests);

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter <= 0;
      else if (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_counter_enable)
          cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter <= cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter_next_value;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_2_in_slavearbiterlockenable <= 0;
      else if ((|cycloneIII_3c120_niosII_standard_sopc_clock_2_in_master_qreq_vector & end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_2_in) | (end_xfer_arb_share_counter_term_cycloneIII_3c120_niosII_standard_sopc_clock_2_in & ~cycloneIII_3c120_niosII_standard_sopc_clock_2_in_non_bursting_master_requests))
          cycloneIII_3c120_niosII_standard_sopc_clock_2_in_slavearbiterlockenable <= |cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge/m1 cycloneIII_3c120_niosII_standard_sopc_clock_2/in arbiterlock, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_slavearbiterlockenable & slow_peripheral_bridge_m1_continuerequest;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_slavearbiterlockenable2 = |cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arb_share_counter_next_value;

  //slow_peripheral_bridge/m1 cycloneIII_3c120_niosII_standard_sopc_clock_2/in arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock2 = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_slavearbiterlockenable2 & slow_peripheral_bridge_m1_continuerequest;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_any_continuerequest = 1;

  //slow_peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  assign slow_peripheral_bridge_m1_continuerequest = 1;

  assign slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in = slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in & ~((slow_peripheral_bridge_m1_read & ((slow_peripheral_bridge_m1_latency_counter != 0))));
  //local readdatavalid slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in & slow_peripheral_bridge_m1_read & ~cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waits_for_read;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_writedata mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_writedata = slow_peripheral_bridge_m1_writedata;

  //assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket;

  //master is always granted when requested
  assign slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in = slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;

  //slow_peripheral_bridge/m1 saved-grant cycloneIII_3c120_niosII_standard_sopc_clock_2/in, which is an e_assign
  assign slow_peripheral_bridge_m1_saved_grant_cycloneIII_3c120_niosII_standard_sopc_clock_2_in = slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;

  //allow new arb cycle for cycloneIII_3c120_niosII_standard_sopc_clock_2/in, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_master_qreq_vector = 1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reset_n assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reset_n = reset_n;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_firsttransfer first transaction, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_firsttransfer = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_begins_xfer ? cycloneIII_3c120_niosII_standard_sopc_clock_2_in_unreg_firsttransfer : cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reg_firsttransfer;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_unreg_firsttransfer first transaction, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_unreg_firsttransfer = ~(cycloneIII_3c120_niosII_standard_sopc_clock_2_in_slavearbiterlockenable & cycloneIII_3c120_niosII_standard_sopc_clock_2_in_any_continuerequest);

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reg_firsttransfer <= 1'b1;
      else if (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_begins_xfer)
          cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reg_firsttransfer <= cycloneIII_3c120_niosII_standard_sopc_clock_2_in_unreg_firsttransfer;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_beginbursttransfer_internal = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_begins_xfer;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_read assignment, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_read = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in & slow_peripheral_bridge_m1_read;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_write assignment, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_write = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in & slow_peripheral_bridge_m1_write;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_address mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_address = slow_peripheral_bridge_m1_address_to_slave;

  //slaveid cycloneIII_3c120_niosII_standard_sopc_clock_2_in_nativeaddress nativeaddress mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_nativeaddress = slow_peripheral_bridge_m1_nativeaddress;

  //d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer <= 1;
      else 
        d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer <= cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waits_for_read in a cycle, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waits_for_read = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_in_a_read_cycle & cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_in_a_read_cycle assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_in_a_read_cycle = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in & slow_peripheral_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_in_a_read_cycle;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waits_for_write in a cycle, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waits_for_write = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_in_a_write_cycle & cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_in_a_write_cycle assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_in_a_write_cycle = slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in & slow_peripheral_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_2_in_in_a_write_cycle;

  assign wait_for_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_counter = 0;
  //cycloneIII_3c120_niosII_standard_sopc_clock_2_in_byteenable byte enable port mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_in_byteenable = (slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in)? slow_peripheral_bridge_m1_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cycloneIII_3c120_niosII_standard_sopc_clock_2/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_clock_2_out_arbitrator (
                                                                      // inputs:
                                                                       clk,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_data_valid_tse_tx_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata,
                                                                       d1_tse_tx_pll_s1_end_xfer,
                                                                       reset_n,
                                                                       tse_tx_pll_s1_readdata_from_sa,

                                                                      // outputs:
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_readdata,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_reset_n,
                                                                       cycloneIII_3c120_niosII_standard_sopc_clock_2_out_waitrequest
                                                                    )
;

  output  [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave;
  output  [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_readdata;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_out_reset_n;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_out_waitrequest;
  input            clk;
  input   [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address;
  input   [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_data_valid_tse_tx_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata;
  input            d1_tse_tx_pll_s1_end_xfer;
  input            reset_n;
  input   [ 15: 0] tse_tx_pll_s1_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_last_time;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave;
  reg     [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable_last_time;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_last_time;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_readdata;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_reset_n;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_run;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_waitrequest;
  reg              cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write_last_time;
  reg     [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata_last_time;
  wire             r_2;
  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & ((~cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1 | ~cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read | (1 & ~d1_tse_tx_pll_s1_end_xfer & cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read))) & ((~cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1 | ~cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write | (1 & cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write)));

  //cascaded wait assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_run = r_2;

  //optimize select-logic by passing only those address bits which matter.
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2/out readdata mux, which is an e_mux
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_readdata = tse_tx_pll_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_waitrequest = ~cycloneIII_3c120_niosII_standard_sopc_clock_2_out_run;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_reset_n assignment, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_2_out_waitrequest & (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read | cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write);
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address != cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable != cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read != cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write != cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write_last_time))
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata_last_time <= 0;
      else 
        cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata_last_time <= cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata != cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata_last_time) & cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write)
        begin
          $write("%0d ns: cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr2_sdram_s1_module (
                                                                      // inputs:
                                                                       clear_fifo,
                                                                       clk,
                                                                       data_in,
                                                                       read,
                                                                       reset_n,
                                                                       sync_reset,
                                                                       write,

                                                                      // outputs:
                                                                       data_out,
                                                                       empty,
                                                                       fifo_contains_ones_n,
                                                                       full
                                                                    )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  wire             full_32;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_31;
  assign empty = !full_0;
  assign full_32 = 0;
  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    0;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ddr2_sdram_s1_arbitrator (
                                  // inputs:
                                   clk,
                                   cpu_ddr_clock_bridge_m1_address_to_slave,
                                   cpu_ddr_clock_bridge_m1_byteenable,
                                   cpu_ddr_clock_bridge_m1_latency_counter,
                                   cpu_ddr_clock_bridge_m1_read,
                                   cpu_ddr_clock_bridge_m1_write,
                                   cpu_ddr_clock_bridge_m1_writedata,
                                   ddr2_sdram_s1_readdata,
                                   ddr2_sdram_s1_readdatavalid,
                                   ddr2_sdram_s1_resetrequest_n,
                                   ddr2_sdram_s1_waitrequest_n,
                                   reset_n,

                                  // outputs:
                                   cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1,
                                   cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1,
                                   cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1,
                                   cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register,
                                   cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1,
                                   d1_ddr2_sdram_s1_end_xfer,
                                   ddr2_sdram_s1_address,
                                   ddr2_sdram_s1_beginbursttransfer,
                                   ddr2_sdram_s1_burstcount,
                                   ddr2_sdram_s1_byteenable,
                                   ddr2_sdram_s1_read,
                                   ddr2_sdram_s1_readdata_from_sa,
                                   ddr2_sdram_s1_resetrequest_n_from_sa,
                                   ddr2_sdram_s1_waitrequest_n_from_sa,
                                   ddr2_sdram_s1_write,
                                   ddr2_sdram_s1_writedata
                                )
;

  output           cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1;
  output           cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1;
  output           cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1;
  output           cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register;
  output           cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1;
  output           d1_ddr2_sdram_s1_end_xfer;
  output  [ 23: 0] ddr2_sdram_s1_address;
  output           ddr2_sdram_s1_beginbursttransfer;
  output  [  2: 0] ddr2_sdram_s1_burstcount;
  output  [  3: 0] ddr2_sdram_s1_byteenable;
  output           ddr2_sdram_s1_read;
  output  [ 31: 0] ddr2_sdram_s1_readdata_from_sa;
  output           ddr2_sdram_s1_resetrequest_n_from_sa;
  output           ddr2_sdram_s1_waitrequest_n_from_sa;
  output           ddr2_sdram_s1_write;
  output  [ 31: 0] ddr2_sdram_s1_writedata;
  input            clk;
  input   [ 25: 0] cpu_ddr_clock_bridge_m1_address_to_slave;
  input   [  3: 0] cpu_ddr_clock_bridge_m1_byteenable;
  input            cpu_ddr_clock_bridge_m1_latency_counter;
  input            cpu_ddr_clock_bridge_m1_read;
  input            cpu_ddr_clock_bridge_m1_write;
  input   [ 31: 0] cpu_ddr_clock_bridge_m1_writedata;
  input   [ 31: 0] ddr2_sdram_s1_readdata;
  input            ddr2_sdram_s1_readdatavalid;
  input            ddr2_sdram_s1_resetrequest_n;
  input            ddr2_sdram_s1_waitrequest_n;
  input            reset_n;

  wire             cpu_ddr_clock_bridge_m1_arbiterlock;
  wire             cpu_ddr_clock_bridge_m1_arbiterlock2;
  wire             cpu_ddr_clock_bridge_m1_continuerequest;
  wire             cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1;
  wire             cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1;
  wire             cpu_ddr_clock_bridge_m1_rdv_fifo_empty_ddr2_sdram_s1;
  wire             cpu_ddr_clock_bridge_m1_rdv_fifo_output_from_ddr2_sdram_s1;
  wire             cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1;
  wire             cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register;
  wire             cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1;
  wire             cpu_ddr_clock_bridge_m1_saved_grant_ddr2_sdram_s1;
  reg              d1_ddr2_sdram_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [ 23: 0] ddr2_sdram_s1_address;
  wire             ddr2_sdram_s1_allgrants;
  wire             ddr2_sdram_s1_allow_new_arb_cycle;
  wire             ddr2_sdram_s1_any_bursting_master_saved_grant;
  wire             ddr2_sdram_s1_any_continuerequest;
  wire             ddr2_sdram_s1_arb_counter_enable;
  reg              ddr2_sdram_s1_arb_share_counter;
  wire             ddr2_sdram_s1_arb_share_counter_next_value;
  wire             ddr2_sdram_s1_arb_share_set_values;
  reg     [  1: 0] ddr2_sdram_s1_bbt_burstcounter;
  wire             ddr2_sdram_s1_beginbursttransfer;
  wire             ddr2_sdram_s1_beginbursttransfer_internal;
  wire             ddr2_sdram_s1_begins_xfer;
  wire    [  2: 0] ddr2_sdram_s1_burstcount;
  wire    [  3: 0] ddr2_sdram_s1_byteenable;
  wire             ddr2_sdram_s1_end_xfer;
  wire             ddr2_sdram_s1_firsttransfer;
  wire             ddr2_sdram_s1_grant_vector;
  wire             ddr2_sdram_s1_in_a_read_cycle;
  wire             ddr2_sdram_s1_in_a_write_cycle;
  wire             ddr2_sdram_s1_master_qreq_vector;
  wire             ddr2_sdram_s1_move_on_to_next_transaction;
  wire    [  1: 0] ddr2_sdram_s1_next_bbt_burstcount;
  wire             ddr2_sdram_s1_non_bursting_master_requests;
  wire             ddr2_sdram_s1_read;
  wire    [ 31: 0] ddr2_sdram_s1_readdata_from_sa;
  wire             ddr2_sdram_s1_readdatavalid_from_sa;
  reg              ddr2_sdram_s1_reg_firsttransfer;
  wire             ddr2_sdram_s1_resetrequest_n_from_sa;
  reg              ddr2_sdram_s1_slavearbiterlockenable;
  wire             ddr2_sdram_s1_slavearbiterlockenable2;
  wire             ddr2_sdram_s1_unreg_firsttransfer;
  wire             ddr2_sdram_s1_waitrequest_n_from_sa;
  wire             ddr2_sdram_s1_waits_for_read;
  wire             ddr2_sdram_s1_waits_for_write;
  wire             ddr2_sdram_s1_write;
  wire    [ 31: 0] ddr2_sdram_s1_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_ddr2_sdram_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 25: 0] shifted_address_to_ddr2_sdram_s1_from_cpu_ddr_clock_bridge_m1;
  wire             wait_for_ddr2_sdram_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~ddr2_sdram_s1_end_xfer;
    end


  assign ddr2_sdram_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1));
  //assign ddr2_sdram_s1_readdata_from_sa = ddr2_sdram_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr2_sdram_s1_readdata_from_sa = ddr2_sdram_s1_readdata;

  assign cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1 = (1) & (cpu_ddr_clock_bridge_m1_read | cpu_ddr_clock_bridge_m1_write);
  //assign ddr2_sdram_s1_waitrequest_n_from_sa = ddr2_sdram_s1_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr2_sdram_s1_waitrequest_n_from_sa = ddr2_sdram_s1_waitrequest_n;

  //assign ddr2_sdram_s1_readdatavalid_from_sa = ddr2_sdram_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr2_sdram_s1_readdatavalid_from_sa = ddr2_sdram_s1_readdatavalid;

  //ddr2_sdram_s1_arb_share_counter set values, which is an e_mux
  assign ddr2_sdram_s1_arb_share_set_values = 1;

  //ddr2_sdram_s1_non_bursting_master_requests mux, which is an e_mux
  assign ddr2_sdram_s1_non_bursting_master_requests = cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1;

  //ddr2_sdram_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign ddr2_sdram_s1_any_bursting_master_saved_grant = 0;

  //ddr2_sdram_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign ddr2_sdram_s1_arb_share_counter_next_value = ddr2_sdram_s1_firsttransfer ? (ddr2_sdram_s1_arb_share_set_values - 1) : |ddr2_sdram_s1_arb_share_counter ? (ddr2_sdram_s1_arb_share_counter - 1) : 0;

  //ddr2_sdram_s1_allgrants all slave grants, which is an e_mux
  assign ddr2_sdram_s1_allgrants = |ddr2_sdram_s1_grant_vector;

  //ddr2_sdram_s1_end_xfer assignment, which is an e_assign
  assign ddr2_sdram_s1_end_xfer = ~(ddr2_sdram_s1_waits_for_read | ddr2_sdram_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_ddr2_sdram_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_ddr2_sdram_s1 = ddr2_sdram_s1_end_xfer & (~ddr2_sdram_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //ddr2_sdram_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign ddr2_sdram_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_ddr2_sdram_s1 & ddr2_sdram_s1_allgrants) | (end_xfer_arb_share_counter_term_ddr2_sdram_s1 & ~ddr2_sdram_s1_non_bursting_master_requests);

  //ddr2_sdram_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_sdram_s1_arb_share_counter <= 0;
      else if (ddr2_sdram_s1_arb_counter_enable)
          ddr2_sdram_s1_arb_share_counter <= ddr2_sdram_s1_arb_share_counter_next_value;
    end


  //ddr2_sdram_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_sdram_s1_slavearbiterlockenable <= 0;
      else if ((|ddr2_sdram_s1_master_qreq_vector & end_xfer_arb_share_counter_term_ddr2_sdram_s1) | (end_xfer_arb_share_counter_term_ddr2_sdram_s1 & ~ddr2_sdram_s1_non_bursting_master_requests))
          ddr2_sdram_s1_slavearbiterlockenable <= |ddr2_sdram_s1_arb_share_counter_next_value;
    end


  //cpu_ddr_clock_bridge/m1 ddr2_sdram/s1 arbiterlock, which is an e_assign
  assign cpu_ddr_clock_bridge_m1_arbiterlock = ddr2_sdram_s1_slavearbiterlockenable & cpu_ddr_clock_bridge_m1_continuerequest;

  //ddr2_sdram_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign ddr2_sdram_s1_slavearbiterlockenable2 = |ddr2_sdram_s1_arb_share_counter_next_value;

  //cpu_ddr_clock_bridge/m1 ddr2_sdram/s1 arbiterlock2, which is an e_assign
  assign cpu_ddr_clock_bridge_m1_arbiterlock2 = ddr2_sdram_s1_slavearbiterlockenable2 & cpu_ddr_clock_bridge_m1_continuerequest;

  //ddr2_sdram_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign ddr2_sdram_s1_any_continuerequest = 1;

  //cpu_ddr_clock_bridge_m1_continuerequest continued request, which is an e_assign
  assign cpu_ddr_clock_bridge_m1_continuerequest = 1;

  assign cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1 = cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1 & ~((cpu_ddr_clock_bridge_m1_read & ((cpu_ddr_clock_bridge_m1_latency_counter != 0) | (1 < cpu_ddr_clock_bridge_m1_latency_counter))));
  //unique name for ddr2_sdram_s1_move_on_to_next_transaction, which is an e_assign
  assign ddr2_sdram_s1_move_on_to_next_transaction = ddr2_sdram_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr2_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr2_sdram_s1_module rdv_fifo_for_cpu_ddr_clock_bridge_m1_to_ddr2_sdram_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1),
      .data_out             (cpu_ddr_clock_bridge_m1_rdv_fifo_output_from_ddr2_sdram_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_ddr_clock_bridge_m1_rdv_fifo_empty_ddr2_sdram_s1),
      .full                 (),
      .read                 (ddr2_sdram_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr2_sdram_s1_waits_for_read)
    );

  assign cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register = ~cpu_ddr_clock_bridge_m1_rdv_fifo_empty_ddr2_sdram_s1;
  //local readdatavalid cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1, which is an e_mux
  assign cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1 = ddr2_sdram_s1_readdatavalid_from_sa;

  //ddr2_sdram_s1_writedata mux, which is an e_mux
  assign ddr2_sdram_s1_writedata = cpu_ddr_clock_bridge_m1_writedata;

  //master is always granted when requested
  assign cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1 = cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1;

  //cpu_ddr_clock_bridge/m1 saved-grant ddr2_sdram/s1, which is an e_assign
  assign cpu_ddr_clock_bridge_m1_saved_grant_ddr2_sdram_s1 = cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1;

  //allow new arb cycle for ddr2_sdram/s1, which is an e_assign
  assign ddr2_sdram_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign ddr2_sdram_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign ddr2_sdram_s1_master_qreq_vector = 1;

  //assign ddr2_sdram_s1_resetrequest_n_from_sa = ddr2_sdram_s1_resetrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr2_sdram_s1_resetrequest_n_from_sa = ddr2_sdram_s1_resetrequest_n;

  //ddr2_sdram_s1_firsttransfer first transaction, which is an e_assign
  assign ddr2_sdram_s1_firsttransfer = ddr2_sdram_s1_begins_xfer ? ddr2_sdram_s1_unreg_firsttransfer : ddr2_sdram_s1_reg_firsttransfer;

  //ddr2_sdram_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign ddr2_sdram_s1_unreg_firsttransfer = ~(ddr2_sdram_s1_slavearbiterlockenable & ddr2_sdram_s1_any_continuerequest);

  //ddr2_sdram_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_sdram_s1_reg_firsttransfer <= 1'b1;
      else if (ddr2_sdram_s1_begins_xfer)
          ddr2_sdram_s1_reg_firsttransfer <= ddr2_sdram_s1_unreg_firsttransfer;
    end


  //ddr2_sdram_s1_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign ddr2_sdram_s1_next_bbt_burstcount = ((((ddr2_sdram_s1_write) && (ddr2_sdram_s1_bbt_burstcounter == 0))))? (ddr2_sdram_s1_burstcount - 1) :
    ((((ddr2_sdram_s1_read) && (ddr2_sdram_s1_bbt_burstcounter == 0))))? 0 :
    (ddr2_sdram_s1_bbt_burstcounter - 1);

  //ddr2_sdram_s1_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr2_sdram_s1_bbt_burstcounter <= 0;
      else if (ddr2_sdram_s1_begins_xfer)
          ddr2_sdram_s1_bbt_burstcounter <= ddr2_sdram_s1_next_bbt_burstcount;
    end


  //ddr2_sdram_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign ddr2_sdram_s1_beginbursttransfer_internal = ddr2_sdram_s1_begins_xfer & (ddr2_sdram_s1_bbt_burstcounter == 0);

  //ddr2_sdram/s1 begin burst transfer to slave, which is an e_assign
  assign ddr2_sdram_s1_beginbursttransfer = ddr2_sdram_s1_beginbursttransfer_internal;

  //ddr2_sdram_s1_read assignment, which is an e_mux
  assign ddr2_sdram_s1_read = cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1 & cpu_ddr_clock_bridge_m1_read;

  //ddr2_sdram_s1_write assignment, which is an e_mux
  assign ddr2_sdram_s1_write = cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1 & cpu_ddr_clock_bridge_m1_write;

  assign shifted_address_to_ddr2_sdram_s1_from_cpu_ddr_clock_bridge_m1 = cpu_ddr_clock_bridge_m1_address_to_slave;
  //ddr2_sdram_s1_address mux, which is an e_mux
  assign ddr2_sdram_s1_address = shifted_address_to_ddr2_sdram_s1_from_cpu_ddr_clock_bridge_m1 >> 2;

  //d1_ddr2_sdram_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_ddr2_sdram_s1_end_xfer <= 1;
      else 
        d1_ddr2_sdram_s1_end_xfer <= ddr2_sdram_s1_end_xfer;
    end


  //ddr2_sdram_s1_waits_for_read in a cycle, which is an e_mux
  assign ddr2_sdram_s1_waits_for_read = ddr2_sdram_s1_in_a_read_cycle & ~ddr2_sdram_s1_waitrequest_n_from_sa;

  //ddr2_sdram_s1_in_a_read_cycle assignment, which is an e_assign
  assign ddr2_sdram_s1_in_a_read_cycle = cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1 & cpu_ddr_clock_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ddr2_sdram_s1_in_a_read_cycle;

  //ddr2_sdram_s1_waits_for_write in a cycle, which is an e_mux
  assign ddr2_sdram_s1_waits_for_write = ddr2_sdram_s1_in_a_write_cycle & ~ddr2_sdram_s1_waitrequest_n_from_sa;

  //ddr2_sdram_s1_in_a_write_cycle assignment, which is an e_assign
  assign ddr2_sdram_s1_in_a_write_cycle = cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1 & cpu_ddr_clock_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ddr2_sdram_s1_in_a_write_cycle;

  assign wait_for_ddr2_sdram_s1_counter = 0;
  //ddr2_sdram_s1_byteenable byte enable port mux, which is an e_mux
  assign ddr2_sdram_s1_byteenable = (cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1)? cpu_ddr_clock_bridge_m1_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign ddr2_sdram_s1_burstcount = 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //ddr2_sdram/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_reset_clk_125_domain_synch_module (
                                                                                 // inputs:
                                                                                  clk,
                                                                                  data_in,
                                                                                  reset_n,

                                                                                 // outputs:
                                                                                  data_out
                                                                               )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module descriptor_memory_s1_arbitrator (
                                         // inputs:
                                          clk,
                                          cpu_data_master_address_to_slave,
                                          cpu_data_master_byteenable,
                                          cpu_data_master_latency_counter,
                                          cpu_data_master_read,
                                          cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                          cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                          cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register,
                                          cpu_data_master_write,
                                          cpu_data_master_writedata,
                                          descriptor_memory_s1_readdata,
                                          reset_n,
                                          sgdma_rx_descriptor_read_address_to_slave,
                                          sgdma_rx_descriptor_read_latency_counter,
                                          sgdma_rx_descriptor_read_read,
                                          sgdma_rx_descriptor_write_address_to_slave,
                                          sgdma_rx_descriptor_write_write,
                                          sgdma_rx_descriptor_write_writedata,
                                          sgdma_tx_descriptor_read_address_to_slave,
                                          sgdma_tx_descriptor_read_latency_counter,
                                          sgdma_tx_descriptor_read_read,
                                          sgdma_tx_descriptor_write_address_to_slave,
                                          sgdma_tx_descriptor_write_write,
                                          sgdma_tx_descriptor_write_writedata,

                                         // outputs:
                                          cpu_data_master_granted_descriptor_memory_s1,
                                          cpu_data_master_qualified_request_descriptor_memory_s1,
                                          cpu_data_master_read_data_valid_descriptor_memory_s1,
                                          cpu_data_master_requests_descriptor_memory_s1,
                                          d1_descriptor_memory_s1_end_xfer,
                                          descriptor_memory_s1_address,
                                          descriptor_memory_s1_byteenable,
                                          descriptor_memory_s1_chipselect,
                                          descriptor_memory_s1_clken,
                                          descriptor_memory_s1_readdata_from_sa,
                                          descriptor_memory_s1_reset,
                                          descriptor_memory_s1_write,
                                          descriptor_memory_s1_writedata,
                                          sgdma_rx_descriptor_read_granted_descriptor_memory_s1,
                                          sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1,
                                          sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1,
                                          sgdma_rx_descriptor_read_requests_descriptor_memory_s1,
                                          sgdma_rx_descriptor_write_granted_descriptor_memory_s1,
                                          sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1,
                                          sgdma_rx_descriptor_write_requests_descriptor_memory_s1,
                                          sgdma_tx_descriptor_read_granted_descriptor_memory_s1,
                                          sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1,
                                          sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1,
                                          sgdma_tx_descriptor_read_requests_descriptor_memory_s1,
                                          sgdma_tx_descriptor_write_granted_descriptor_memory_s1,
                                          sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1,
                                          sgdma_tx_descriptor_write_requests_descriptor_memory_s1
                                       )
;

  output           cpu_data_master_granted_descriptor_memory_s1;
  output           cpu_data_master_qualified_request_descriptor_memory_s1;
  output           cpu_data_master_read_data_valid_descriptor_memory_s1;
  output           cpu_data_master_requests_descriptor_memory_s1;
  output           d1_descriptor_memory_s1_end_xfer;
  output  [  9: 0] descriptor_memory_s1_address;
  output  [  3: 0] descriptor_memory_s1_byteenable;
  output           descriptor_memory_s1_chipselect;
  output           descriptor_memory_s1_clken;
  output  [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  output           descriptor_memory_s1_reset;
  output           descriptor_memory_s1_write;
  output  [ 31: 0] descriptor_memory_s1_writedata;
  output           sgdma_rx_descriptor_read_granted_descriptor_memory_s1;
  output           sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;
  output           sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;
  output           sgdma_rx_descriptor_read_requests_descriptor_memory_s1;
  output           sgdma_rx_descriptor_write_granted_descriptor_memory_s1;
  output           sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;
  output           sgdma_rx_descriptor_write_requests_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_granted_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;
  output           sgdma_tx_descriptor_read_requests_descriptor_memory_s1;
  output           sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  output           sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;
  output           sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 31: 0] descriptor_memory_s1_readdata;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  input            sgdma_rx_descriptor_read_latency_counter;
  input            sgdma_rx_descriptor_read_read;
  input   [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  input            sgdma_rx_descriptor_write_write;
  input   [ 31: 0] sgdma_rx_descriptor_write_writedata;
  input   [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  input            sgdma_tx_descriptor_read_latency_counter;
  input            sgdma_tx_descriptor_read_read;
  input   [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  input            sgdma_tx_descriptor_write_write;
  input   [ 31: 0] sgdma_tx_descriptor_write_writedata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_descriptor_memory_s1;
  wire             cpu_data_master_qualified_request_descriptor_memory_s1;
  wire             cpu_data_master_read_data_valid_descriptor_memory_s1;
  reg              cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register;
  wire             cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in;
  wire             cpu_data_master_requests_descriptor_memory_s1;
  wire             cpu_data_master_saved_grant_descriptor_memory_s1;
  reg              d1_descriptor_memory_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [  9: 0] descriptor_memory_s1_address;
  wire             descriptor_memory_s1_allgrants;
  wire             descriptor_memory_s1_allow_new_arb_cycle;
  wire             descriptor_memory_s1_any_bursting_master_saved_grant;
  wire             descriptor_memory_s1_any_continuerequest;
  reg     [  4: 0] descriptor_memory_s1_arb_addend;
  wire             descriptor_memory_s1_arb_counter_enable;
  reg     [  3: 0] descriptor_memory_s1_arb_share_counter;
  wire    [  3: 0] descriptor_memory_s1_arb_share_counter_next_value;
  wire    [  3: 0] descriptor_memory_s1_arb_share_set_values;
  wire    [  4: 0] descriptor_memory_s1_arb_winner;
  wire             descriptor_memory_s1_arbitration_holdoff_internal;
  wire             descriptor_memory_s1_beginbursttransfer_internal;
  wire             descriptor_memory_s1_begins_xfer;
  wire    [  3: 0] descriptor_memory_s1_byteenable;
  wire             descriptor_memory_s1_chipselect;
  wire    [  9: 0] descriptor_memory_s1_chosen_master_double_vector;
  wire    [  4: 0] descriptor_memory_s1_chosen_master_rot_left;
  wire             descriptor_memory_s1_clken;
  wire             descriptor_memory_s1_end_xfer;
  wire             descriptor_memory_s1_firsttransfer;
  wire    [  4: 0] descriptor_memory_s1_grant_vector;
  wire             descriptor_memory_s1_in_a_read_cycle;
  wire             descriptor_memory_s1_in_a_write_cycle;
  wire    [  4: 0] descriptor_memory_s1_master_qreq_vector;
  wire             descriptor_memory_s1_non_bursting_master_requests;
  wire    [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  reg              descriptor_memory_s1_reg_firsttransfer;
  wire             descriptor_memory_s1_reset;
  reg     [  4: 0] descriptor_memory_s1_saved_chosen_master_vector;
  reg              descriptor_memory_s1_slavearbiterlockenable;
  wire             descriptor_memory_s1_slavearbiterlockenable2;
  wire             descriptor_memory_s1_unreg_firsttransfer;
  wire             descriptor_memory_s1_waits_for_read;
  wire             descriptor_memory_s1_waits_for_write;
  wire             descriptor_memory_s1_write;
  wire    [ 31: 0] descriptor_memory_s1_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_descriptor_memory_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1;
  reg              last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1;
  reg              last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1;
  reg              last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1;
  reg              last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1;
  wire             p1_cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register;
  wire             p1_sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
  wire             p1_sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
  wire             sgdma_rx_descriptor_read_arbiterlock;
  wire             sgdma_rx_descriptor_read_arbiterlock2;
  wire             sgdma_rx_descriptor_read_continuerequest;
  wire             sgdma_rx_descriptor_read_granted_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;
  reg              sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
  wire             sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in;
  wire             sgdma_rx_descriptor_read_requests_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_arbiterlock;
  wire             sgdma_rx_descriptor_write_arbiterlock2;
  wire             sgdma_rx_descriptor_write_continuerequest;
  wire             sgdma_rx_descriptor_write_granted_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_requests_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_arbiterlock;
  wire             sgdma_tx_descriptor_read_arbiterlock2;
  wire             sgdma_tx_descriptor_read_continuerequest;
  wire             sgdma_tx_descriptor_read_granted_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;
  reg              sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
  wire             sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in;
  wire             sgdma_tx_descriptor_read_requests_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_arbiterlock;
  wire             sgdma_tx_descriptor_write_arbiterlock2;
  wire             sgdma_tx_descriptor_write_continuerequest;
  wire             sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1;
  wire    [ 28: 0] shifted_address_to_descriptor_memory_s1_from_cpu_data_master;
  wire    [ 31: 0] shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read;
  wire    [ 31: 0] shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write;
  wire    [ 31: 0] shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read;
  wire    [ 31: 0] shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write;
  wire             wait_for_descriptor_memory_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~descriptor_memory_s1_end_xfer;
    end


  assign descriptor_memory_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_descriptor_memory_s1 | sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 | sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 | sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 | sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1));
  //assign descriptor_memory_s1_readdata_from_sa = descriptor_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign descriptor_memory_s1_readdata_from_sa = descriptor_memory_s1_readdata;

  assign cpu_data_master_requests_descriptor_memory_s1 = ({cpu_data_master_address_to_slave[28 : 12] , 12'b0} == 29'h1000000) & (cpu_data_master_read | cpu_data_master_write);
  //descriptor_memory_s1_arb_share_counter set values, which is an e_mux
  assign descriptor_memory_s1_arb_share_set_values = (sgdma_rx_descriptor_read_granted_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_read_granted_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_write_granted_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_read_granted_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_read_granted_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_write_granted_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_read_granted_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_read_granted_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_write_granted_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_read_granted_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_read_granted_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_write_granted_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_read_granted_descriptor_memory_s1)? 8 :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_read_granted_descriptor_memory_s1)? 8 :
    (sgdma_tx_descriptor_write_granted_descriptor_memory_s1)? 8 :
    1;

  //descriptor_memory_s1_non_bursting_master_requests mux, which is an e_mux
  assign descriptor_memory_s1_non_bursting_master_requests = cpu_data_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1 |
    cpu_data_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1 |
    cpu_data_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1 |
    cpu_data_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1 |
    cpu_data_master_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_rx_descriptor_write_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_read_requests_descriptor_memory_s1 |
    sgdma_tx_descriptor_write_requests_descriptor_memory_s1;

  //descriptor_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign descriptor_memory_s1_any_bursting_master_saved_grant = 0;

  //descriptor_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign descriptor_memory_s1_arb_share_counter_next_value = descriptor_memory_s1_firsttransfer ? (descriptor_memory_s1_arb_share_set_values - 1) : |descriptor_memory_s1_arb_share_counter ? (descriptor_memory_s1_arb_share_counter - 1) : 0;

  //descriptor_memory_s1_allgrants all slave grants, which is an e_mux
  assign descriptor_memory_s1_allgrants = (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector) |
    (|descriptor_memory_s1_grant_vector);

  //descriptor_memory_s1_end_xfer assignment, which is an e_assign
  assign descriptor_memory_s1_end_xfer = ~(descriptor_memory_s1_waits_for_read | descriptor_memory_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_descriptor_memory_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_descriptor_memory_s1 = descriptor_memory_s1_end_xfer & (~descriptor_memory_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //descriptor_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign descriptor_memory_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_descriptor_memory_s1 & descriptor_memory_s1_allgrants) | (end_xfer_arb_share_counter_term_descriptor_memory_s1 & ~descriptor_memory_s1_non_bursting_master_requests);

  //descriptor_memory_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_arb_share_counter <= 0;
      else if (descriptor_memory_s1_arb_counter_enable)
          descriptor_memory_s1_arb_share_counter <= descriptor_memory_s1_arb_share_counter_next_value;
    end


  //descriptor_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_slavearbiterlockenable <= 0;
      else if ((|descriptor_memory_s1_master_qreq_vector & end_xfer_arb_share_counter_term_descriptor_memory_s1) | (end_xfer_arb_share_counter_term_descriptor_memory_s1 & ~descriptor_memory_s1_non_bursting_master_requests))
          descriptor_memory_s1_slavearbiterlockenable <= |descriptor_memory_s1_arb_share_counter_next_value;
    end


  //cpu/data_master descriptor_memory/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //descriptor_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign descriptor_memory_s1_slavearbiterlockenable2 = |descriptor_memory_s1_arb_share_counter_next_value;

  //cpu/data_master descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //sgdma_rx/descriptor_read descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_rx_descriptor_read_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & sgdma_rx_descriptor_read_continuerequest;

  //sgdma_rx/descriptor_read descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_rx_descriptor_read_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & sgdma_rx_descriptor_read_continuerequest;

  //sgdma_rx/descriptor_read granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 <= sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_rx_descriptor_read_requests_descriptor_memory_s1) ? 0 : last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1;
    end


  //sgdma_rx_descriptor_read_continuerequest continued request, which is an e_mux
  assign sgdma_rx_descriptor_read_continuerequest = (last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_read_requests_descriptor_memory_s1);

  //descriptor_memory_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign descriptor_memory_s1_any_continuerequest = sgdma_rx_descriptor_read_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    cpu_data_master_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    cpu_data_master_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_read_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    cpu_data_master_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_write_continuerequest |
    cpu_data_master_continuerequest |
    sgdma_rx_descriptor_read_continuerequest |
    sgdma_rx_descriptor_write_continuerequest |
    sgdma_tx_descriptor_read_continuerequest;

  //sgdma_rx/descriptor_write descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_rx_descriptor_write_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & sgdma_rx_descriptor_write_continuerequest;

  //sgdma_rx/descriptor_write descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_rx_descriptor_write_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & sgdma_rx_descriptor_write_continuerequest;

  //sgdma_rx/descriptor_write granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 <= sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_rx_descriptor_write_requests_descriptor_memory_s1) ? 0 : last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1;
    end


  //sgdma_rx_descriptor_write_continuerequest continued request, which is an e_mux
  assign sgdma_rx_descriptor_write_continuerequest = (last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_rx_descriptor_write_requests_descriptor_memory_s1);

  //sgdma_tx/descriptor_read descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_tx_descriptor_read_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & sgdma_tx_descriptor_read_continuerequest;

  //sgdma_tx/descriptor_read descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_tx_descriptor_read_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & sgdma_tx_descriptor_read_continuerequest;

  //sgdma_tx/descriptor_read granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 <= sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_tx_descriptor_read_requests_descriptor_memory_s1) ? 0 : last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1;
    end


  //sgdma_tx_descriptor_read_continuerequest continued request, which is an e_mux
  assign sgdma_tx_descriptor_read_continuerequest = (last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_read_requests_descriptor_memory_s1);

  //sgdma_tx/descriptor_write descriptor_memory/s1 arbiterlock, which is an e_assign
  assign sgdma_tx_descriptor_write_arbiterlock = descriptor_memory_s1_slavearbiterlockenable & sgdma_tx_descriptor_write_continuerequest;

  //sgdma_tx/descriptor_write descriptor_memory/s1 arbiterlock2, which is an e_assign
  assign sgdma_tx_descriptor_write_arbiterlock2 = descriptor_memory_s1_slavearbiterlockenable2 & sgdma_tx_descriptor_write_continuerequest;

  //sgdma_tx/descriptor_write granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 <= sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~sgdma_tx_descriptor_write_requests_descriptor_memory_s1) ? 0 : last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1;
    end


  //sgdma_tx_descriptor_write_continuerequest continued request, which is an e_mux
  assign sgdma_tx_descriptor_write_continuerequest = (last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_descriptor_memory_s1) |
    (last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 & sgdma_tx_descriptor_write_requests_descriptor_memory_s1);

  assign cpu_data_master_qualified_request_descriptor_memory_s1 = cpu_data_master_requests_descriptor_memory_s1 & ~((cpu_data_master_read & ((1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register))) | sgdma_rx_descriptor_read_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_read_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  //cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in = cpu_data_master_granted_descriptor_memory_s1 & cpu_data_master_read & ~descriptor_memory_s1_waits_for_read;

  //shift register p1 cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register = {cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register, cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in};

  //cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register <= 0;
      else 
        cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register <= p1_cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register;
    end


  //local readdatavalid cpu_data_master_read_data_valid_descriptor_memory_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_descriptor_memory_s1 = cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register;

  //descriptor_memory_s1_writedata mux, which is an e_mux
  assign descriptor_memory_s1_writedata = (cpu_data_master_granted_descriptor_memory_s1)? cpu_data_master_writedata :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? sgdma_rx_descriptor_write_writedata :
    sgdma_tx_descriptor_write_writedata;

  //mux descriptor_memory_s1_clken, which is an e_mux
  assign descriptor_memory_s1_clken = 1'b1;

  assign sgdma_rx_descriptor_read_requests_descriptor_memory_s1 = (({sgdma_rx_descriptor_read_address_to_slave[31 : 12] , 12'b0} == 32'h1000000) & (sgdma_rx_descriptor_read_read)) & sgdma_rx_descriptor_read_read;
  //cpu/data_master granted descriptor_memory/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 <= cpu_data_master_saved_grant_descriptor_memory_s1 ? 1 : (descriptor_memory_s1_arbitration_holdoff_internal | ~cpu_data_master_requests_descriptor_memory_s1) ? 0 : last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = (last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 & cpu_data_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 & cpu_data_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 & cpu_data_master_requests_descriptor_memory_s1) |
    (last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 & cpu_data_master_requests_descriptor_memory_s1);

  assign sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 = sgdma_rx_descriptor_read_requests_descriptor_memory_s1 & ~(cpu_data_master_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_read_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  //sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in = sgdma_rx_descriptor_read_granted_descriptor_memory_s1 & sgdma_rx_descriptor_read_read & ~descriptor_memory_s1_waits_for_read;

  //shift register p1 sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register = {sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register, sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in};

  //sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= 0;
      else 
        sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= p1_sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
    end


  //local readdatavalid sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1, which is an e_mux
  assign sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1 = sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;

  assign sgdma_rx_descriptor_write_requests_descriptor_memory_s1 = (({sgdma_rx_descriptor_write_address_to_slave[31 : 12] , 12'b0} == 32'h1000000) & (sgdma_rx_descriptor_write_write)) & sgdma_rx_descriptor_write_write;
  assign sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 = sgdma_rx_descriptor_write_requests_descriptor_memory_s1 & ~(cpu_data_master_arbiterlock | sgdma_rx_descriptor_read_arbiterlock | sgdma_tx_descriptor_read_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  assign sgdma_tx_descriptor_read_requests_descriptor_memory_s1 = (({sgdma_tx_descriptor_read_address_to_slave[31 : 12] , 12'b0} == 32'h1000000) & (sgdma_tx_descriptor_read_read)) & sgdma_tx_descriptor_read_read;
  assign sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 = sgdma_tx_descriptor_read_requests_descriptor_memory_s1 & ~(cpu_data_master_arbiterlock | sgdma_rx_descriptor_read_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_write_arbiterlock);
  //sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in = sgdma_tx_descriptor_read_granted_descriptor_memory_s1 & sgdma_tx_descriptor_read_read & ~descriptor_memory_s1_waits_for_read;

  //shift register p1 sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register = {sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register, sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in};

  //sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= 0;
      else 
        sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= p1_sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
    end


  //local readdatavalid sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1, which is an e_mux
  assign sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1 = sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;

  assign sgdma_tx_descriptor_write_requests_descriptor_memory_s1 = (({sgdma_tx_descriptor_write_address_to_slave[31 : 12] , 12'b0} == 32'h1000000) & (sgdma_tx_descriptor_write_write)) & sgdma_tx_descriptor_write_write;
  assign sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 = sgdma_tx_descriptor_write_requests_descriptor_memory_s1 & ~(cpu_data_master_arbiterlock | sgdma_rx_descriptor_read_arbiterlock | sgdma_rx_descriptor_write_arbiterlock | sgdma_tx_descriptor_read_arbiterlock);
  //allow new arb cycle for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~sgdma_rx_descriptor_read_arbiterlock & ~sgdma_rx_descriptor_write_arbiterlock & ~sgdma_tx_descriptor_read_arbiterlock & ~sgdma_tx_descriptor_write_arbiterlock;

  //sgdma_tx/descriptor_write assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[0] = sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;

  //sgdma_tx/descriptor_write grant descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_write_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[0];

  //sgdma_tx/descriptor_write saved-grant descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[0] && sgdma_tx_descriptor_write_requests_descriptor_memory_s1;

  //sgdma_tx/descriptor_read assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[1] = sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;

  //sgdma_tx/descriptor_read grant descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_read_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[1];

  //sgdma_tx/descriptor_read saved-grant descriptor_memory/s1, which is an e_assign
  assign sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[1] && sgdma_tx_descriptor_read_requests_descriptor_memory_s1;

  //sgdma_rx/descriptor_write assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[2] = sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;

  //sgdma_rx/descriptor_write grant descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_write_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[2];

  //sgdma_rx/descriptor_write saved-grant descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[2] && sgdma_rx_descriptor_write_requests_descriptor_memory_s1;

  //sgdma_rx/descriptor_read assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[3] = sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;

  //sgdma_rx/descriptor_read grant descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_read_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[3];

  //sgdma_rx/descriptor_read saved-grant descriptor_memory/s1, which is an e_assign
  assign sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[3] && sgdma_rx_descriptor_read_requests_descriptor_memory_s1;

  //cpu/data_master assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  assign descriptor_memory_s1_master_qreq_vector[4] = cpu_data_master_qualified_request_descriptor_memory_s1;

  //cpu/data_master grant descriptor_memory/s1, which is an e_assign
  assign cpu_data_master_granted_descriptor_memory_s1 = descriptor_memory_s1_grant_vector[4];

  //cpu/data_master saved-grant descriptor_memory/s1, which is an e_assign
  assign cpu_data_master_saved_grant_descriptor_memory_s1 = descriptor_memory_s1_arb_winner[4] && cpu_data_master_requests_descriptor_memory_s1;

  //descriptor_memory/s1 chosen-master double-vector, which is an e_assign
  assign descriptor_memory_s1_chosen_master_double_vector = {descriptor_memory_s1_master_qreq_vector, descriptor_memory_s1_master_qreq_vector} & ({~descriptor_memory_s1_master_qreq_vector, ~descriptor_memory_s1_master_qreq_vector} + descriptor_memory_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign descriptor_memory_s1_arb_winner = (descriptor_memory_s1_allow_new_arb_cycle & | descriptor_memory_s1_grant_vector) ? descriptor_memory_s1_grant_vector : descriptor_memory_s1_saved_chosen_master_vector;

  //saved descriptor_memory_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_saved_chosen_master_vector <= 0;
      else if (descriptor_memory_s1_allow_new_arb_cycle)
          descriptor_memory_s1_saved_chosen_master_vector <= |descriptor_memory_s1_grant_vector ? descriptor_memory_s1_grant_vector : descriptor_memory_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign descriptor_memory_s1_grant_vector = {(descriptor_memory_s1_chosen_master_double_vector[4] | descriptor_memory_s1_chosen_master_double_vector[9]),
    (descriptor_memory_s1_chosen_master_double_vector[3] | descriptor_memory_s1_chosen_master_double_vector[8]),
    (descriptor_memory_s1_chosen_master_double_vector[2] | descriptor_memory_s1_chosen_master_double_vector[7]),
    (descriptor_memory_s1_chosen_master_double_vector[1] | descriptor_memory_s1_chosen_master_double_vector[6]),
    (descriptor_memory_s1_chosen_master_double_vector[0] | descriptor_memory_s1_chosen_master_double_vector[5])};

  //descriptor_memory/s1 chosen master rotated left, which is an e_assign
  assign descriptor_memory_s1_chosen_master_rot_left = (descriptor_memory_s1_arb_winner << 1) ? (descriptor_memory_s1_arb_winner << 1) : 1;

  //descriptor_memory/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_arb_addend <= 1;
      else if (|descriptor_memory_s1_grant_vector)
          descriptor_memory_s1_arb_addend <= descriptor_memory_s1_end_xfer? descriptor_memory_s1_chosen_master_rot_left : descriptor_memory_s1_grant_vector;
    end


  //~descriptor_memory_s1_reset assignment, which is an e_assign
  assign descriptor_memory_s1_reset = ~reset_n;

  assign descriptor_memory_s1_chipselect = cpu_data_master_granted_descriptor_memory_s1 | sgdma_rx_descriptor_read_granted_descriptor_memory_s1 | sgdma_rx_descriptor_write_granted_descriptor_memory_s1 | sgdma_tx_descriptor_read_granted_descriptor_memory_s1 | sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  //descriptor_memory_s1_firsttransfer first transaction, which is an e_assign
  assign descriptor_memory_s1_firsttransfer = descriptor_memory_s1_begins_xfer ? descriptor_memory_s1_unreg_firsttransfer : descriptor_memory_s1_reg_firsttransfer;

  //descriptor_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign descriptor_memory_s1_unreg_firsttransfer = ~(descriptor_memory_s1_slavearbiterlockenable & descriptor_memory_s1_any_continuerequest);

  //descriptor_memory_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          descriptor_memory_s1_reg_firsttransfer <= 1'b1;
      else if (descriptor_memory_s1_begins_xfer)
          descriptor_memory_s1_reg_firsttransfer <= descriptor_memory_s1_unreg_firsttransfer;
    end


  //descriptor_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign descriptor_memory_s1_beginbursttransfer_internal = descriptor_memory_s1_begins_xfer;

  //descriptor_memory_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign descriptor_memory_s1_arbitration_holdoff_internal = descriptor_memory_s1_begins_xfer & descriptor_memory_s1_firsttransfer;

  //descriptor_memory_s1_write assignment, which is an e_mux
  assign descriptor_memory_s1_write = (cpu_data_master_granted_descriptor_memory_s1 & cpu_data_master_write) | (sgdma_rx_descriptor_write_granted_descriptor_memory_s1 & sgdma_rx_descriptor_write_write) | (sgdma_tx_descriptor_write_granted_descriptor_memory_s1 & sgdma_tx_descriptor_write_write);

  assign shifted_address_to_descriptor_memory_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //descriptor_memory_s1_address mux, which is an e_mux
  assign descriptor_memory_s1_address = (cpu_data_master_granted_descriptor_memory_s1)? (shifted_address_to_descriptor_memory_s1_from_cpu_data_master >> 2) :
    (sgdma_rx_descriptor_read_granted_descriptor_memory_s1)? (shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read >> 2) :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? (shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write >> 2) :
    (sgdma_tx_descriptor_read_granted_descriptor_memory_s1)? (shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read >> 2) :
    (shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write >> 2);

  assign shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read = sgdma_rx_descriptor_read_address_to_slave;
  assign shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write = sgdma_rx_descriptor_write_address_to_slave;
  assign shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read = sgdma_tx_descriptor_read_address_to_slave;
  assign shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write = sgdma_tx_descriptor_write_address_to_slave;
  //d1_descriptor_memory_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_descriptor_memory_s1_end_xfer <= 1;
      else 
        d1_descriptor_memory_s1_end_xfer <= descriptor_memory_s1_end_xfer;
    end


  //descriptor_memory_s1_waits_for_read in a cycle, which is an e_mux
  assign descriptor_memory_s1_waits_for_read = descriptor_memory_s1_in_a_read_cycle & 0;

  //descriptor_memory_s1_in_a_read_cycle assignment, which is an e_assign
  assign descriptor_memory_s1_in_a_read_cycle = (cpu_data_master_granted_descriptor_memory_s1 & cpu_data_master_read) | (sgdma_rx_descriptor_read_granted_descriptor_memory_s1 & sgdma_rx_descriptor_read_read) | (sgdma_tx_descriptor_read_granted_descriptor_memory_s1 & sgdma_tx_descriptor_read_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = descriptor_memory_s1_in_a_read_cycle;

  //descriptor_memory_s1_waits_for_write in a cycle, which is an e_mux
  assign descriptor_memory_s1_waits_for_write = descriptor_memory_s1_in_a_write_cycle & 0;

  //descriptor_memory_s1_in_a_write_cycle assignment, which is an e_assign
  assign descriptor_memory_s1_in_a_write_cycle = (cpu_data_master_granted_descriptor_memory_s1 & cpu_data_master_write) | (sgdma_rx_descriptor_write_granted_descriptor_memory_s1 & sgdma_rx_descriptor_write_write) | (sgdma_tx_descriptor_write_granted_descriptor_memory_s1 & sgdma_tx_descriptor_write_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = descriptor_memory_s1_in_a_write_cycle;

  assign wait_for_descriptor_memory_s1_counter = 0;
  //descriptor_memory_s1_byteenable byte enable port mux, which is an e_mux
  assign descriptor_memory_s1_byteenable = (cpu_data_master_granted_descriptor_memory_s1)? cpu_data_master_byteenable :
    (sgdma_rx_descriptor_write_granted_descriptor_memory_s1)? {4 {1'b1}} :
    (sgdma_tx_descriptor_write_granted_descriptor_memory_s1)? {4 {1'b1}} :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //descriptor_memory/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_descriptor_memory_s1 + sgdma_rx_descriptor_read_granted_descriptor_memory_s1 + sgdma_rx_descriptor_write_granted_descriptor_memory_s1 + sgdma_tx_descriptor_read_granted_descriptor_memory_s1 + sgdma_tx_descriptor_write_granted_descriptor_memory_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_descriptor_memory_s1 + sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1 + sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1 + sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1 + sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module flash_tristate_bridge_avalon_slave_arbitrator (
                                                       // inputs:
                                                        clk,
                                                        pipeline_bridge_before_tristate_bridge_m1_address_to_slave,
                                                        pipeline_bridge_before_tristate_bridge_m1_burstcount,
                                                        pipeline_bridge_before_tristate_bridge_m1_byteenable,
                                                        pipeline_bridge_before_tristate_bridge_m1_chipselect,
                                                        pipeline_bridge_before_tristate_bridge_m1_dbs_address,
                                                        pipeline_bridge_before_tristate_bridge_m1_dbs_write_16,
                                                        pipeline_bridge_before_tristate_bridge_m1_latency_counter,
                                                        pipeline_bridge_before_tristate_bridge_m1_read,
                                                        pipeline_bridge_before_tristate_bridge_m1_write,
                                                        pipeline_bridge_before_tristate_bridge_m1_writedata,
                                                        reset_n,

                                                       // outputs:
                                                        cs_n_to_the_max2,
                                                        d1_flash_tristate_bridge_avalon_slave_end_xfer,
                                                        ext_flash_s1_wait_counter_eq_0,
                                                        flash_tristate_bridge_address,
                                                        flash_tristate_bridge_data,
                                                        incoming_flash_tristate_bridge_data,
                                                        incoming_flash_tristate_bridge_data_with_Xs_converted_to_0,
                                                        max2_s1_wait_counter_eq_0,
                                                        oe_n_to_the_max2,
                                                        pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1,
                                                        pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1,
                                                        pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1,
                                                        pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1,
                                                        pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1,
                                                        pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1,
                                                        pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1,
                                                        pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1,
                                                        pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1,
                                                        read_n_to_the_ext_flash,
                                                        select_n_to_the_ext_flash,
                                                        we_n_to_the_max2,
                                                        write_n_to_the_ext_flash
                                                     )
;

  output           cs_n_to_the_max2;
  output           d1_flash_tristate_bridge_avalon_slave_end_xfer;
  output           ext_flash_s1_wait_counter_eq_0;
  output  [ 25: 0] flash_tristate_bridge_address;
  inout   [ 31: 0] flash_tristate_bridge_data;
  output  [ 31: 0] incoming_flash_tristate_bridge_data;
  output  [ 15: 0] incoming_flash_tristate_bridge_data_with_Xs_converted_to_0;
  output           max2_s1_wait_counter_eq_0;
  output           oe_n_to_the_max2;
  output  [  1: 0] pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1;
  output           pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1;
  output           pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1;
  output           pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1;
  output           pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1;
  output           pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1;
  output           pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1;
  output           pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1;
  output           pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1;
  output           read_n_to_the_ext_flash;
  output           select_n_to_the_ext_flash;
  output           we_n_to_the_max2;
  output           write_n_to_the_ext_flash;
  input            clk;
  input   [ 26: 0] pipeline_bridge_before_tristate_bridge_m1_address_to_slave;
  input            pipeline_bridge_before_tristate_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_before_tristate_bridge_m1_byteenable;
  input            pipeline_bridge_before_tristate_bridge_m1_chipselect;
  input   [  1: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_address;
  input   [ 15: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_write_16;
  input   [  1: 0] pipeline_bridge_before_tristate_bridge_m1_latency_counter;
  input            pipeline_bridge_before_tristate_bridge_m1_read;
  input            pipeline_bridge_before_tristate_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_before_tristate_bridge_m1_writedata;
  input            reset_n;

  reg              cs_n_to_the_max2 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_flash_tristate_bridge_avalon_slave_end_xfer;
  reg              d1_in_a_write_cycle /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_ENABLE_REGISTER=ON"  */;
  reg     [ 31: 0] d1_outgoing_flash_tristate_bridge_data /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave;
  wire    [  3: 0] ext_flash_s1_counter_load_value;
  wire             ext_flash_s1_in_a_read_cycle;
  wire             ext_flash_s1_in_a_write_cycle;
  reg     [  3: 0] ext_flash_s1_wait_counter;
  wire             ext_flash_s1_wait_counter_eq_0;
  wire             ext_flash_s1_waits_for_read;
  wire             ext_flash_s1_waits_for_write;
  wire             ext_flash_s1_with_write_latency;
  reg     [ 25: 0] flash_tristate_bridge_address /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             flash_tristate_bridge_avalon_slave_allgrants;
  wire             flash_tristate_bridge_avalon_slave_allow_new_arb_cycle;
  wire             flash_tristate_bridge_avalon_slave_any_bursting_master_saved_grant;
  wire             flash_tristate_bridge_avalon_slave_any_continuerequest;
  wire             flash_tristate_bridge_avalon_slave_arb_counter_enable;
  reg     [  1: 0] flash_tristate_bridge_avalon_slave_arb_share_counter;
  wire    [  1: 0] flash_tristate_bridge_avalon_slave_arb_share_counter_next_value;
  wire    [  1: 0] flash_tristate_bridge_avalon_slave_arb_share_set_values;
  wire             flash_tristate_bridge_avalon_slave_beginbursttransfer_internal;
  wire             flash_tristate_bridge_avalon_slave_begins_xfer;
  wire             flash_tristate_bridge_avalon_slave_end_xfer;
  wire             flash_tristate_bridge_avalon_slave_firsttransfer;
  wire             flash_tristate_bridge_avalon_slave_grant_vector;
  wire             flash_tristate_bridge_avalon_slave_master_qreq_vector;
  wire             flash_tristate_bridge_avalon_slave_non_bursting_master_requests;
  wire             flash_tristate_bridge_avalon_slave_read_pending;
  reg              flash_tristate_bridge_avalon_slave_reg_firsttransfer;
  reg              flash_tristate_bridge_avalon_slave_slavearbiterlockenable;
  wire             flash_tristate_bridge_avalon_slave_slavearbiterlockenable2;
  wire             flash_tristate_bridge_avalon_slave_unreg_firsttransfer;
  wire             flash_tristate_bridge_avalon_slave_write_pending;
  wire    [ 31: 0] flash_tristate_bridge_data;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg     [ 31: 0] incoming_flash_tristate_bridge_data /* synthesis ALTERA_ATTRIBUTE = "FAST_INPUT_REGISTER=ON"  */;
  wire             incoming_flash_tristate_bridge_data_bit_0_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_10_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_11_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_12_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_13_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_14_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_15_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_1_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_2_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_3_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_4_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_5_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_6_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_7_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_8_is_x;
  wire             incoming_flash_tristate_bridge_data_bit_9_is_x;
  wire    [ 15: 0] incoming_flash_tristate_bridge_data_with_Xs_converted_to_0;
  wire    [  3: 0] max2_s1_counter_load_value;
  wire             max2_s1_in_a_read_cycle;
  wire             max2_s1_in_a_write_cycle;
  reg     [  3: 0] max2_s1_wait_counter;
  wire             max2_s1_wait_counter_eq_0;
  wire             max2_s1_waits_for_read;
  wire             max2_s1_waits_for_write;
  wire             max2_s1_with_write_latency;
  reg              oe_n_to_the_max2 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire    [ 31: 0] outgoing_flash_tristate_bridge_data;
  wire             p1_cs_n_to_the_max2;
  wire    [ 25: 0] p1_flash_tristate_bridge_address;
  wire             p1_oe_n_to_the_max2;
  wire    [  1: 0] p1_pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register;
  wire    [  1: 0] p1_pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register;
  wire             p1_read_n_to_the_ext_flash;
  wire             p1_select_n_to_the_ext_flash;
  wire             p1_we_n_to_the_max2;
  wire             p1_write_n_to_the_ext_flash;
  wire             pipeline_bridge_before_tristate_bridge_m1_arbiterlock;
  wire             pipeline_bridge_before_tristate_bridge_m1_arbiterlock2;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1_segment_0;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1_segment_1;
  wire             pipeline_bridge_before_tristate_bridge_m1_continuerequest;
  wire             pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1;
  reg     [  1: 0] pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register;
  wire             pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register_in;
  wire             pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1;
  reg     [  1: 0] pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register;
  wire             pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register_in;
  wire             pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_saved_grant_ext_flash_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_saved_grant_max2_s1;
  reg              read_n_to_the_ext_flash /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              select_n_to_the_ext_flash /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             time_to_write;
  wire             wait_for_ext_flash_s1_counter;
  wire             wait_for_max2_s1_counter;
  reg              we_n_to_the_max2 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              write_n_to_the_ext_flash /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~flash_tristate_bridge_avalon_slave_end_xfer;
    end


  assign flash_tristate_bridge_avalon_slave_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1 | pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1));
  assign pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1 = ({pipeline_bridge_before_tristate_bridge_m1_address_to_slave[26 : 5] , 5'b0} == 27'h14000000) & pipeline_bridge_before_tristate_bridge_m1_chipselect;
  //~cs_n_to_the_max2 of type chipselect to ~p1_cs_n_to_the_max2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cs_n_to_the_max2 <= ~0;
      else 
        cs_n_to_the_max2 <= p1_cs_n_to_the_max2;
    end


  //~select_n_to_the_ext_flash of type chipselect to ~p1_select_n_to_the_ext_flash, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          select_n_to_the_ext_flash <= ~0;
      else 
        select_n_to_the_ext_flash <= p1_select_n_to_the_ext_flash;
    end


  assign flash_tristate_bridge_avalon_slave_write_pending = 0;
  //flash_tristate_bridge/avalon_slave read pending calc, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_read_pending = 0;

  //flash_tristate_bridge_avalon_slave_arb_share_counter set values, which is an e_mux
  assign flash_tristate_bridge_avalon_slave_arb_share_set_values = (pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1)? 2 :
    1;

  //flash_tristate_bridge_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  assign flash_tristate_bridge_avalon_slave_non_bursting_master_requests = pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1 |
    pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1;

  //flash_tristate_bridge_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign flash_tristate_bridge_avalon_slave_any_bursting_master_saved_grant = 0;

  //flash_tristate_bridge_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_arb_share_counter_next_value = flash_tristate_bridge_avalon_slave_firsttransfer ? (flash_tristate_bridge_avalon_slave_arb_share_set_values - 1) : |flash_tristate_bridge_avalon_slave_arb_share_counter ? (flash_tristate_bridge_avalon_slave_arb_share_counter - 1) : 0;

  //flash_tristate_bridge_avalon_slave_allgrants all slave grants, which is an e_mux
  assign flash_tristate_bridge_avalon_slave_allgrants = (|flash_tristate_bridge_avalon_slave_grant_vector) |
    (|flash_tristate_bridge_avalon_slave_grant_vector);

  //flash_tristate_bridge_avalon_slave_end_xfer assignment, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_end_xfer = ~(max2_s1_waits_for_read | max2_s1_waits_for_write | ext_flash_s1_waits_for_read | ext_flash_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave = flash_tristate_bridge_avalon_slave_end_xfer & (~flash_tristate_bridge_avalon_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //flash_tristate_bridge_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave & flash_tristate_bridge_avalon_slave_allgrants) | (end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave & ~flash_tristate_bridge_avalon_slave_non_bursting_master_requests);

  //flash_tristate_bridge_avalon_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_avalon_slave_arb_share_counter <= 0;
      else if (flash_tristate_bridge_avalon_slave_arb_counter_enable)
          flash_tristate_bridge_avalon_slave_arb_share_counter <= flash_tristate_bridge_avalon_slave_arb_share_counter_next_value;
    end


  //flash_tristate_bridge_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_avalon_slave_slavearbiterlockenable <= 0;
      else if ((|flash_tristate_bridge_avalon_slave_master_qreq_vector & end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave) | (end_xfer_arb_share_counter_term_flash_tristate_bridge_avalon_slave & ~flash_tristate_bridge_avalon_slave_non_bursting_master_requests))
          flash_tristate_bridge_avalon_slave_slavearbiterlockenable <= |flash_tristate_bridge_avalon_slave_arb_share_counter_next_value;
    end


  //pipeline_bridge_before_tristate_bridge/m1 flash_tristate_bridge/avalon_slave arbiterlock, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_m1_arbiterlock = flash_tristate_bridge_avalon_slave_slavearbiterlockenable & pipeline_bridge_before_tristate_bridge_m1_continuerequest;

  //flash_tristate_bridge_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_slavearbiterlockenable2 = |flash_tristate_bridge_avalon_slave_arb_share_counter_next_value;

  //pipeline_bridge_before_tristate_bridge/m1 flash_tristate_bridge/avalon_slave arbiterlock2, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_m1_arbiterlock2 = flash_tristate_bridge_avalon_slave_slavearbiterlockenable2 & pipeline_bridge_before_tristate_bridge_m1_continuerequest;

  //flash_tristate_bridge_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_any_continuerequest = 1;

  //pipeline_bridge_before_tristate_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1 = pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1 & ~(((pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect) & (flash_tristate_bridge_avalon_slave_write_pending | (flash_tristate_bridge_avalon_slave_read_pending) | (2 < pipeline_bridge_before_tristate_bridge_m1_latency_counter))) | ((flash_tristate_bridge_avalon_slave_read_pending) & (pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect)));
  //pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register_in = pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1 & (pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect) & ~max2_s1_waits_for_read;

  //shift register p1 pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register = {pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register, pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register_in};

  //pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register <= p1_pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register;
    end


  //local readdatavalid pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1 = pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1_shift_register[1];

  //flash_tristate_bridge_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          incoming_flash_tristate_bridge_data <= 0;
      else 
        incoming_flash_tristate_bridge_data <= flash_tristate_bridge_data;
    end


  //max2_s1_with_write_latency assignment, which is an e_assign
  assign max2_s1_with_write_latency = in_a_write_cycle & (pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1);

  //time to write the data, which is an e_mux
  assign time_to_write = (max2_s1_with_write_latency)? 1 :
    (ext_flash_s1_with_write_latency)? 1 :
    0;

  //d1_outgoing_flash_tristate_bridge_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_outgoing_flash_tristate_bridge_data <= 0;
      else 
        d1_outgoing_flash_tristate_bridge_data <= outgoing_flash_tristate_bridge_data;
    end


  //write cycle delayed by 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_in_a_write_cycle <= 0;
      else 
        d1_in_a_write_cycle <= time_to_write;
    end


  //d1_outgoing_flash_tristate_bridge_data tristate driver, which is an e_assign
  assign flash_tristate_bridge_data = (d1_in_a_write_cycle)? d1_outgoing_flash_tristate_bridge_data:{32{1'bz}};

  //outgoing_flash_tristate_bridge_data mux, which is an e_mux
  assign outgoing_flash_tristate_bridge_data = (pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1)? pipeline_bridge_before_tristate_bridge_m1_writedata :
    pipeline_bridge_before_tristate_bridge_m1_dbs_write_16;

  assign pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1 = ({pipeline_bridge_before_tristate_bridge_m1_address_to_slave[26] , 26'b0} == 27'h10000000) & pipeline_bridge_before_tristate_bridge_m1_chipselect;
  assign pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1 = pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1 & ~(((pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect) & (flash_tristate_bridge_avalon_slave_write_pending | (flash_tristate_bridge_avalon_slave_read_pending) | (2 < pipeline_bridge_before_tristate_bridge_m1_latency_counter))) | ((flash_tristate_bridge_avalon_slave_read_pending | !pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1) & (pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect)));
  //pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register_in = pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1 & (pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect) & ~ext_flash_s1_waits_for_read;

  //shift register p1 pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register = {pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register, pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register_in};

  //pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register <= p1_pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register;
    end


  //local readdatavalid pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1 = pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1_shift_register[1];

  //ext_flash_s1_with_write_latency assignment, which is an e_assign
  assign ext_flash_s1_with_write_latency = in_a_write_cycle & (pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1);

  //master is always granted when requested
  assign pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1 = pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1;

  //pipeline_bridge_before_tristate_bridge/m1 saved-grant max2/s1, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_m1_saved_grant_max2_s1 = pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1;

  //allow new arb cycle for flash_tristate_bridge/avalon_slave, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign flash_tristate_bridge_avalon_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign flash_tristate_bridge_avalon_slave_master_qreq_vector = 1;

  //master is always granted when requested
  assign pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1 = pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1;

  //pipeline_bridge_before_tristate_bridge/m1 saved-grant ext_flash/s1, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_m1_saved_grant_ext_flash_s1 = pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1;

  assign p1_cs_n_to_the_max2 = ~pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1;
  //flash_tristate_bridge_avalon_slave_firsttransfer first transaction, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_firsttransfer = flash_tristate_bridge_avalon_slave_begins_xfer ? flash_tristate_bridge_avalon_slave_unreg_firsttransfer : flash_tristate_bridge_avalon_slave_reg_firsttransfer;

  //flash_tristate_bridge_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_unreg_firsttransfer = ~(flash_tristate_bridge_avalon_slave_slavearbiterlockenable & flash_tristate_bridge_avalon_slave_any_continuerequest);

  //flash_tristate_bridge_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_avalon_slave_reg_firsttransfer <= 1'b1;
      else if (flash_tristate_bridge_avalon_slave_begins_xfer)
          flash_tristate_bridge_avalon_slave_reg_firsttransfer <= flash_tristate_bridge_avalon_slave_unreg_firsttransfer;
    end


  //flash_tristate_bridge_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign flash_tristate_bridge_avalon_slave_beginbursttransfer_internal = flash_tristate_bridge_avalon_slave_begins_xfer;

  //~oe_n_to_the_max2 of type read to ~p1_oe_n_to_the_max2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          oe_n_to_the_max2 <= ~0;
      else 
        oe_n_to_the_max2 <= p1_oe_n_to_the_max2;
    end


  //~p1_oe_n_to_the_max2 assignment, which is an e_mux
  assign p1_oe_n_to_the_max2 = ~(pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1 & (pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect));

  //~we_n_to_the_max2 of type write to ~p1_we_n_to_the_max2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          we_n_to_the_max2 <= ~0;
      else 
        we_n_to_the_max2 <= p1_we_n_to_the_max2;
    end


  //~p1_we_n_to_the_max2 assignment, which is an e_mux
  assign p1_we_n_to_the_max2 = ~(pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1 & (pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect));

  //flash_tristate_bridge_address of type address to p1_flash_tristate_bridge_address, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          flash_tristate_bridge_address <= 0;
      else 
        flash_tristate_bridge_address <= p1_flash_tristate_bridge_address;
    end


  //p1_flash_tristate_bridge_address mux, which is an e_mux
  assign p1_flash_tristate_bridge_address = (pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1)? pipeline_bridge_before_tristate_bridge_m1_address_to_slave :
    ({pipeline_bridge_before_tristate_bridge_m1_address_to_slave >> 2,
    pipeline_bridge_before_tristate_bridge_m1_dbs_address[1],
    {1 {1'b0}}});

  //d1_flash_tristate_bridge_avalon_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_flash_tristate_bridge_avalon_slave_end_xfer <= 1;
      else 
        d1_flash_tristate_bridge_avalon_slave_end_xfer <= flash_tristate_bridge_avalon_slave_end_xfer;
    end


  //max2_s1_waits_for_read in a cycle, which is an e_mux
  assign max2_s1_waits_for_read = max2_s1_in_a_read_cycle & wait_for_max2_s1_counter;

  //max2_s1_in_a_read_cycle assignment, which is an e_assign
  assign max2_s1_in_a_read_cycle = pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1 & (pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = max2_s1_in_a_read_cycle |
    ext_flash_s1_in_a_read_cycle;

  //max2_s1_waits_for_write in a cycle, which is an e_mux
  assign max2_s1_waits_for_write = max2_s1_in_a_write_cycle & wait_for_max2_s1_counter;

  //max2_s1_in_a_write_cycle assignment, which is an e_assign
  assign max2_s1_in_a_write_cycle = pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1 & (pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = max2_s1_in_a_write_cycle |
    ext_flash_s1_in_a_write_cycle;

  assign max2_s1_wait_counter_eq_0 = max2_s1_wait_counter == 0;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          max2_s1_wait_counter <= 0;
      else 
        max2_s1_wait_counter <= max2_s1_counter_load_value;
    end


  assign max2_s1_counter_load_value = ((max2_s1_in_a_write_cycle & flash_tristate_bridge_avalon_slave_begins_xfer))? 8 :
    ((max2_s1_in_a_read_cycle & flash_tristate_bridge_avalon_slave_begins_xfer))? 8 :
    (~max2_s1_wait_counter_eq_0)? max2_s1_wait_counter - 1 :
    0;

  assign wait_for_max2_s1_counter = flash_tristate_bridge_avalon_slave_begins_xfer | ~max2_s1_wait_counter_eq_0;
  assign p1_select_n_to_the_ext_flash = ~pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1;
  //~read_n_to_the_ext_flash of type read to ~p1_read_n_to_the_ext_flash, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          read_n_to_the_ext_flash <= ~0;
      else 
        read_n_to_the_ext_flash <= p1_read_n_to_the_ext_flash;
    end


  //~p1_read_n_to_the_ext_flash assignment, which is an e_mux
  assign p1_read_n_to_the_ext_flash = ~(((pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1 & (pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect)))& ~flash_tristate_bridge_avalon_slave_begins_xfer & (ext_flash_s1_wait_counter < 4));

  //~write_n_to_the_ext_flash of type write to ~p1_write_n_to_the_ext_flash, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_n_to_the_ext_flash <= ~0;
      else 
        write_n_to_the_ext_flash <= p1_write_n_to_the_ext_flash;
    end


  //~p1_write_n_to_the_ext_flash assignment, which is an e_mux
  assign p1_write_n_to_the_ext_flash = ~(((pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1 & (pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect))) & ~flash_tristate_bridge_avalon_slave_begins_xfer & (ext_flash_s1_wait_counter >= 2) & (ext_flash_s1_wait_counter < 6));

  //ext_flash_s1_waits_for_read in a cycle, which is an e_mux
  assign ext_flash_s1_waits_for_read = ext_flash_s1_in_a_read_cycle & wait_for_ext_flash_s1_counter;

  //ext_flash_s1_in_a_read_cycle assignment, which is an e_assign
  assign ext_flash_s1_in_a_read_cycle = pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1 & (pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect);

  //ext_flash_s1_waits_for_write in a cycle, which is an e_mux
  assign ext_flash_s1_waits_for_write = ext_flash_s1_in_a_write_cycle & wait_for_ext_flash_s1_counter;

  //ext_flash_s1_in_a_write_cycle assignment, which is an e_assign
  assign ext_flash_s1_in_a_write_cycle = pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1 & (pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect);

  assign ext_flash_s1_wait_counter_eq_0 = ext_flash_s1_wait_counter == 0;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_flash_s1_wait_counter <= 0;
      else 
        ext_flash_s1_wait_counter <= ext_flash_s1_counter_load_value;
    end


  assign ext_flash_s1_counter_load_value = ((ext_flash_s1_in_a_read_cycle & flash_tristate_bridge_avalon_slave_begins_xfer))? 10 :
    ((ext_flash_s1_in_a_write_cycle & flash_tristate_bridge_avalon_slave_begins_xfer))? 12 :
    (~ext_flash_s1_wait_counter_eq_0)? ext_flash_s1_wait_counter - 1 :
    0;

  assign wait_for_ext_flash_s1_counter = flash_tristate_bridge_avalon_slave_begins_xfer | ~ext_flash_s1_wait_counter_eq_0;
  assign {pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1_segment_1,
pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1_segment_0} = pipeline_bridge_before_tristate_bridge_m1_byteenable;
  assign pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1 = ((pipeline_bridge_before_tristate_bridge_m1_dbs_address[1] == 0))? pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1_segment_0 :
    pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //max2/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge_before_tristate_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1 && (pipeline_bridge_before_tristate_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge_before_tristate_bridge/m1 drove 0 on its 'burstcount' port while accessing slave max2/s1", $time);
          $stop;
        end
    end


  //incoming_flash_tristate_bridge_data_bit_0_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_0_is_x = ^(incoming_flash_tristate_bridge_data[0]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[0] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[0] = incoming_flash_tristate_bridge_data_bit_0_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[0];

  //incoming_flash_tristate_bridge_data_bit_1_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_1_is_x = ^(incoming_flash_tristate_bridge_data[1]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[1] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[1] = incoming_flash_tristate_bridge_data_bit_1_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[1];

  //incoming_flash_tristate_bridge_data_bit_2_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_2_is_x = ^(incoming_flash_tristate_bridge_data[2]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[2] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[2] = incoming_flash_tristate_bridge_data_bit_2_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[2];

  //incoming_flash_tristate_bridge_data_bit_3_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_3_is_x = ^(incoming_flash_tristate_bridge_data[3]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[3] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[3] = incoming_flash_tristate_bridge_data_bit_3_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[3];

  //incoming_flash_tristate_bridge_data_bit_4_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_4_is_x = ^(incoming_flash_tristate_bridge_data[4]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[4] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[4] = incoming_flash_tristate_bridge_data_bit_4_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[4];

  //incoming_flash_tristate_bridge_data_bit_5_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_5_is_x = ^(incoming_flash_tristate_bridge_data[5]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[5] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[5] = incoming_flash_tristate_bridge_data_bit_5_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[5];

  //incoming_flash_tristate_bridge_data_bit_6_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_6_is_x = ^(incoming_flash_tristate_bridge_data[6]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[6] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[6] = incoming_flash_tristate_bridge_data_bit_6_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[6];

  //incoming_flash_tristate_bridge_data_bit_7_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_7_is_x = ^(incoming_flash_tristate_bridge_data[7]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[7] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[7] = incoming_flash_tristate_bridge_data_bit_7_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[7];

  //incoming_flash_tristate_bridge_data_bit_8_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_8_is_x = ^(incoming_flash_tristate_bridge_data[8]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[8] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[8] = incoming_flash_tristate_bridge_data_bit_8_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[8];

  //incoming_flash_tristate_bridge_data_bit_9_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_9_is_x = ^(incoming_flash_tristate_bridge_data[9]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[9] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[9] = incoming_flash_tristate_bridge_data_bit_9_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[9];

  //incoming_flash_tristate_bridge_data_bit_10_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_10_is_x = ^(incoming_flash_tristate_bridge_data[10]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[10] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[10] = incoming_flash_tristate_bridge_data_bit_10_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[10];

  //incoming_flash_tristate_bridge_data_bit_11_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_11_is_x = ^(incoming_flash_tristate_bridge_data[11]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[11] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[11] = incoming_flash_tristate_bridge_data_bit_11_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[11];

  //incoming_flash_tristate_bridge_data_bit_12_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_12_is_x = ^(incoming_flash_tristate_bridge_data[12]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[12] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[12] = incoming_flash_tristate_bridge_data_bit_12_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[12];

  //incoming_flash_tristate_bridge_data_bit_13_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_13_is_x = ^(incoming_flash_tristate_bridge_data[13]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[13] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[13] = incoming_flash_tristate_bridge_data_bit_13_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[13];

  //incoming_flash_tristate_bridge_data_bit_14_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_14_is_x = ^(incoming_flash_tristate_bridge_data[14]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[14] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[14] = incoming_flash_tristate_bridge_data_bit_14_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[14];

  //incoming_flash_tristate_bridge_data_bit_15_is_x x check, which is an e_assign_is_x
  assign incoming_flash_tristate_bridge_data_bit_15_is_x = ^(incoming_flash_tristate_bridge_data[15]) === 1'bx;

  //Crush incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[15] Xs to 0, which is an e_assign
  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[15] = incoming_flash_tristate_bridge_data_bit_15_is_x ? 1'b0 : incoming_flash_tristate_bridge_data[15];

  //ext_flash/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1 + pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_before_tristate_bridge_m1_saved_grant_ext_flash_s1 + pipeline_bridge_before_tristate_bridge_m1_saved_grant_max2_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  
//  assign incoming_flash_tristate_bridge_data_with_Xs_converted_to_0 = incoming_flash_tristate_bridge_data;
//
//synthesis read_comments_as_HDL off

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module flash_tristate_bridge_bridge_arbitrator 
;



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module high_res_timer_s1_arbitrator (
                                      // inputs:
                                       clk,
                                       high_res_timer_s1_irq,
                                       high_res_timer_s1_readdata,
                                       reset_n,
                                       slow_peripheral_bridge_m1_address_to_slave,
                                       slow_peripheral_bridge_m1_latency_counter,
                                       slow_peripheral_bridge_m1_nativeaddress,
                                       slow_peripheral_bridge_m1_read,
                                       slow_peripheral_bridge_m1_write,
                                       slow_peripheral_bridge_m1_writedata,

                                      // outputs:
                                       d1_high_res_timer_s1_end_xfer,
                                       high_res_timer_s1_address,
                                       high_res_timer_s1_chipselect,
                                       high_res_timer_s1_irq_from_sa,
                                       high_res_timer_s1_readdata_from_sa,
                                       high_res_timer_s1_reset_n,
                                       high_res_timer_s1_write_n,
                                       high_res_timer_s1_writedata,
                                       slow_peripheral_bridge_m1_granted_high_res_timer_s1,
                                       slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1,
                                       slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1,
                                       slow_peripheral_bridge_m1_requests_high_res_timer_s1
                                    )
;

  output           d1_high_res_timer_s1_end_xfer;
  output  [  2: 0] high_res_timer_s1_address;
  output           high_res_timer_s1_chipselect;
  output           high_res_timer_s1_irq_from_sa;
  output  [ 15: 0] high_res_timer_s1_readdata_from_sa;
  output           high_res_timer_s1_reset_n;
  output           high_res_timer_s1_write_n;
  output  [ 15: 0] high_res_timer_s1_writedata;
  output           slow_peripheral_bridge_m1_granted_high_res_timer_s1;
  output           slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1;
  output           slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1;
  output           slow_peripheral_bridge_m1_requests_high_res_timer_s1;
  input            clk;
  input            high_res_timer_s1_irq;
  input   [ 15: 0] high_res_timer_s1_readdata;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  input            slow_peripheral_bridge_m1_latency_counter;
  input   [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] slow_peripheral_bridge_m1_writedata;

  reg              d1_high_res_timer_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_high_res_timer_s1;
  wire    [  2: 0] high_res_timer_s1_address;
  wire             high_res_timer_s1_allgrants;
  wire             high_res_timer_s1_allow_new_arb_cycle;
  wire             high_res_timer_s1_any_bursting_master_saved_grant;
  wire             high_res_timer_s1_any_continuerequest;
  wire             high_res_timer_s1_arb_counter_enable;
  reg              high_res_timer_s1_arb_share_counter;
  wire             high_res_timer_s1_arb_share_counter_next_value;
  wire             high_res_timer_s1_arb_share_set_values;
  wire             high_res_timer_s1_beginbursttransfer_internal;
  wire             high_res_timer_s1_begins_xfer;
  wire             high_res_timer_s1_chipselect;
  wire             high_res_timer_s1_end_xfer;
  wire             high_res_timer_s1_firsttransfer;
  wire             high_res_timer_s1_grant_vector;
  wire             high_res_timer_s1_in_a_read_cycle;
  wire             high_res_timer_s1_in_a_write_cycle;
  wire             high_res_timer_s1_irq_from_sa;
  wire             high_res_timer_s1_master_qreq_vector;
  wire             high_res_timer_s1_non_bursting_master_requests;
  wire    [ 15: 0] high_res_timer_s1_readdata_from_sa;
  reg              high_res_timer_s1_reg_firsttransfer;
  wire             high_res_timer_s1_reset_n;
  reg              high_res_timer_s1_slavearbiterlockenable;
  wire             high_res_timer_s1_slavearbiterlockenable2;
  wire             high_res_timer_s1_unreg_firsttransfer;
  wire             high_res_timer_s1_waits_for_read;
  wire             high_res_timer_s1_waits_for_write;
  wire             high_res_timer_s1_write_n;
  wire    [ 15: 0] high_res_timer_s1_writedata;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             slow_peripheral_bridge_m1_arbiterlock;
  wire             slow_peripheral_bridge_m1_arbiterlock2;
  wire             slow_peripheral_bridge_m1_continuerequest;
  wire             slow_peripheral_bridge_m1_granted_high_res_timer_s1;
  wire             slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1;
  wire             slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1;
  wire             slow_peripheral_bridge_m1_requests_high_res_timer_s1;
  wire             slow_peripheral_bridge_m1_saved_grant_high_res_timer_s1;
  wire             wait_for_high_res_timer_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~high_res_timer_s1_end_xfer;
    end


  assign high_res_timer_s1_begins_xfer = ~d1_reasons_to_wait & ((slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1));
  //assign high_res_timer_s1_readdata_from_sa = high_res_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign high_res_timer_s1_readdata_from_sa = high_res_timer_s1_readdata;

  assign slow_peripheral_bridge_m1_requests_high_res_timer_s1 = ({slow_peripheral_bridge_m1_address_to_slave[7 : 5] , 5'b0} == 8'h0) & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write);
  //high_res_timer_s1_arb_share_counter set values, which is an e_mux
  assign high_res_timer_s1_arb_share_set_values = 1;

  //high_res_timer_s1_non_bursting_master_requests mux, which is an e_mux
  assign high_res_timer_s1_non_bursting_master_requests = slow_peripheral_bridge_m1_requests_high_res_timer_s1;

  //high_res_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign high_res_timer_s1_any_bursting_master_saved_grant = 0;

  //high_res_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign high_res_timer_s1_arb_share_counter_next_value = high_res_timer_s1_firsttransfer ? (high_res_timer_s1_arb_share_set_values - 1) : |high_res_timer_s1_arb_share_counter ? (high_res_timer_s1_arb_share_counter - 1) : 0;

  //high_res_timer_s1_allgrants all slave grants, which is an e_mux
  assign high_res_timer_s1_allgrants = |high_res_timer_s1_grant_vector;

  //high_res_timer_s1_end_xfer assignment, which is an e_assign
  assign high_res_timer_s1_end_xfer = ~(high_res_timer_s1_waits_for_read | high_res_timer_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_high_res_timer_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_high_res_timer_s1 = high_res_timer_s1_end_xfer & (~high_res_timer_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //high_res_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign high_res_timer_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_high_res_timer_s1 & high_res_timer_s1_allgrants) | (end_xfer_arb_share_counter_term_high_res_timer_s1 & ~high_res_timer_s1_non_bursting_master_requests);

  //high_res_timer_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          high_res_timer_s1_arb_share_counter <= 0;
      else if (high_res_timer_s1_arb_counter_enable)
          high_res_timer_s1_arb_share_counter <= high_res_timer_s1_arb_share_counter_next_value;
    end


  //high_res_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          high_res_timer_s1_slavearbiterlockenable <= 0;
      else if ((|high_res_timer_s1_master_qreq_vector & end_xfer_arb_share_counter_term_high_res_timer_s1) | (end_xfer_arb_share_counter_term_high_res_timer_s1 & ~high_res_timer_s1_non_bursting_master_requests))
          high_res_timer_s1_slavearbiterlockenable <= |high_res_timer_s1_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge/m1 high_res_timer/s1 arbiterlock, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock = high_res_timer_s1_slavearbiterlockenable & slow_peripheral_bridge_m1_continuerequest;

  //high_res_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign high_res_timer_s1_slavearbiterlockenable2 = |high_res_timer_s1_arb_share_counter_next_value;

  //slow_peripheral_bridge/m1 high_res_timer/s1 arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock2 = high_res_timer_s1_slavearbiterlockenable2 & slow_peripheral_bridge_m1_continuerequest;

  //high_res_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign high_res_timer_s1_any_continuerequest = 1;

  //slow_peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  assign slow_peripheral_bridge_m1_continuerequest = 1;

  assign slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1 = slow_peripheral_bridge_m1_requests_high_res_timer_s1 & ~((slow_peripheral_bridge_m1_read & ((slow_peripheral_bridge_m1_latency_counter != 0))));
  //local readdatavalid slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1 = slow_peripheral_bridge_m1_granted_high_res_timer_s1 & slow_peripheral_bridge_m1_read & ~high_res_timer_s1_waits_for_read;

  //high_res_timer_s1_writedata mux, which is an e_mux
  assign high_res_timer_s1_writedata = slow_peripheral_bridge_m1_writedata;

  //master is always granted when requested
  assign slow_peripheral_bridge_m1_granted_high_res_timer_s1 = slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1;

  //slow_peripheral_bridge/m1 saved-grant high_res_timer/s1, which is an e_assign
  assign slow_peripheral_bridge_m1_saved_grant_high_res_timer_s1 = slow_peripheral_bridge_m1_requests_high_res_timer_s1;

  //allow new arb cycle for high_res_timer/s1, which is an e_assign
  assign high_res_timer_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign high_res_timer_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign high_res_timer_s1_master_qreq_vector = 1;

  //high_res_timer_s1_reset_n assignment, which is an e_assign
  assign high_res_timer_s1_reset_n = reset_n;

  assign high_res_timer_s1_chipselect = slow_peripheral_bridge_m1_granted_high_res_timer_s1;
  //high_res_timer_s1_firsttransfer first transaction, which is an e_assign
  assign high_res_timer_s1_firsttransfer = high_res_timer_s1_begins_xfer ? high_res_timer_s1_unreg_firsttransfer : high_res_timer_s1_reg_firsttransfer;

  //high_res_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign high_res_timer_s1_unreg_firsttransfer = ~(high_res_timer_s1_slavearbiterlockenable & high_res_timer_s1_any_continuerequest);

  //high_res_timer_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          high_res_timer_s1_reg_firsttransfer <= 1'b1;
      else if (high_res_timer_s1_begins_xfer)
          high_res_timer_s1_reg_firsttransfer <= high_res_timer_s1_unreg_firsttransfer;
    end


  //high_res_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign high_res_timer_s1_beginbursttransfer_internal = high_res_timer_s1_begins_xfer;

  //~high_res_timer_s1_write_n assignment, which is an e_mux
  assign high_res_timer_s1_write_n = ~(slow_peripheral_bridge_m1_granted_high_res_timer_s1 & slow_peripheral_bridge_m1_write);

  //high_res_timer_s1_address mux, which is an e_mux
  assign high_res_timer_s1_address = slow_peripheral_bridge_m1_nativeaddress;

  //d1_high_res_timer_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_high_res_timer_s1_end_xfer <= 1;
      else 
        d1_high_res_timer_s1_end_xfer <= high_res_timer_s1_end_xfer;
    end


  //high_res_timer_s1_waits_for_read in a cycle, which is an e_mux
  assign high_res_timer_s1_waits_for_read = high_res_timer_s1_in_a_read_cycle & high_res_timer_s1_begins_xfer;

  //high_res_timer_s1_in_a_read_cycle assignment, which is an e_assign
  assign high_res_timer_s1_in_a_read_cycle = slow_peripheral_bridge_m1_granted_high_res_timer_s1 & slow_peripheral_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = high_res_timer_s1_in_a_read_cycle;

  //high_res_timer_s1_waits_for_write in a cycle, which is an e_mux
  assign high_res_timer_s1_waits_for_write = high_res_timer_s1_in_a_write_cycle & 0;

  //high_res_timer_s1_in_a_write_cycle assignment, which is an e_assign
  assign high_res_timer_s1_in_a_write_cycle = slow_peripheral_bridge_m1_granted_high_res_timer_s1 & slow_peripheral_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = high_res_timer_s1_in_a_write_cycle;

  assign wait_for_high_res_timer_s1_counter = 0;
  //assign high_res_timer_s1_irq_from_sa = high_res_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign high_res_timer_s1_irq_from_sa = high_res_timer_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //high_res_timer/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_avalon_jtag_slave_arbitrator (
                                                // inputs:
                                                 clk,
                                                 jtag_uart_avalon_jtag_slave_dataavailable,
                                                 jtag_uart_avalon_jtag_slave_irq,
                                                 jtag_uart_avalon_jtag_slave_readdata,
                                                 jtag_uart_avalon_jtag_slave_readyfordata,
                                                 jtag_uart_avalon_jtag_slave_waitrequest,
                                                 reset_n,
                                                 slow_peripheral_bridge_m1_address_to_slave,
                                                 slow_peripheral_bridge_m1_latency_counter,
                                                 slow_peripheral_bridge_m1_nativeaddress,
                                                 slow_peripheral_bridge_m1_read,
                                                 slow_peripheral_bridge_m1_write,
                                                 slow_peripheral_bridge_m1_writedata,

                                                // outputs:
                                                 d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                                 jtag_uart_avalon_jtag_slave_address,
                                                 jtag_uart_avalon_jtag_slave_chipselect,
                                                 jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
                                                 jtag_uart_avalon_jtag_slave_irq_from_sa,
                                                 jtag_uart_avalon_jtag_slave_read_n,
                                                 jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_reset_n,
                                                 jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                                 jtag_uart_avalon_jtag_slave_write_n,
                                                 jtag_uart_avalon_jtag_slave_writedata,
                                                 slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave,
                                                 slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave,
                                                 slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
                                                 slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave
                                              )
;

  output           d1_jtag_uart_avalon_jtag_slave_end_xfer;
  output           jtag_uart_avalon_jtag_slave_address;
  output           jtag_uart_avalon_jtag_slave_chipselect;
  output           jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_avalon_jtag_slave_reset_n;
  output           jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  output           slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  output           slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  output           slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  output           slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  input            clk;
  input            jtag_uart_avalon_jtag_slave_dataavailable;
  input            jtag_uart_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  input            jtag_uart_avalon_jtag_slave_readyfordata;
  input            jtag_uart_avalon_jtag_slave_waitrequest;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  input            slow_peripheral_bridge_m1_latency_counter;
  input   [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] slow_peripheral_bridge_m1_writedata;

  reg              d1_jtag_uart_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_allgrants;
  wire             jtag_uart_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_avalon_jtag_slave_arb_counter_enable;
  reg              jtag_uart_avalon_jtag_slave_arb_share_counter;
  wire             jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
  wire             jtag_uart_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  reg              jtag_uart_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire             slow_peripheral_bridge_m1_arbiterlock;
  wire             slow_peripheral_bridge_m1_arbiterlock2;
  wire             slow_peripheral_bridge_m1_continuerequest;
  wire             slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  wire             slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  wire             slow_peripheral_bridge_m1_saved_grant_jtag_uart_avalon_jtag_slave;
  wire             wait_for_jtag_uart_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave));
  //assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata;

  assign slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave = ({slow_peripheral_bridge_m1_address_to_slave[7 : 3] , 3'b0} == 8'he0) & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write);
  //assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest;

  //jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_non_bursting_master_requests = slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave;

  //jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_avalon_jtag_slave_firsttransfer ? (jtag_uart_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_avalon_jtag_slave_arb_share_counter ? (jtag_uart_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_allgrants = |jtag_uart_avalon_jtag_slave_grant_vector;

  //jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_end_xfer = ~(jtag_uart_avalon_jtag_slave_waits_for_read | jtag_uart_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave = jtag_uart_avalon_jtag_slave_end_xfer & (~jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & jtag_uart_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge/m1 jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock = jtag_uart_avalon_jtag_slave_slavearbiterlockenable & slow_peripheral_bridge_m1_continuerequest;

  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;

  //slow_peripheral_bridge/m1 jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock2 = jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 & slow_peripheral_bridge_m1_continuerequest;

  //jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_any_continuerequest = 1;

  //slow_peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  assign slow_peripheral_bridge_m1_continuerequest = 1;

  assign slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave = slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave & ~((slow_peripheral_bridge_m1_read & ((slow_peripheral_bridge_m1_latency_counter != 0))));
  //local readdatavalid slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave = slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave & slow_peripheral_bridge_m1_read & ~jtag_uart_avalon_jtag_slave_waits_for_read;

  //jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_writedata = slow_peripheral_bridge_m1_writedata;

  //master is always granted when requested
  assign slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave = slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;

  //slow_peripheral_bridge/m1 saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  assign slow_peripheral_bridge_m1_saved_grant_jtag_uart_avalon_jtag_slave = slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_avalon_jtag_slave_chipselect = slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  //jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_firsttransfer = jtag_uart_avalon_jtag_slave_begins_xfer ? jtag_uart_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_avalon_jtag_slave_begins_xfer)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_read_n = ~(slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave & slow_peripheral_bridge_m1_read);

  //~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_write_n = ~(slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave & slow_peripheral_bridge_m1_write);

  //jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_address = slow_peripheral_bridge_m1_nativeaddress;

  //d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_read = jtag_uart_avalon_jtag_slave_in_a_read_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_read_cycle = slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave & slow_peripheral_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_write = jtag_uart_avalon_jtag_slave_in_a_write_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_write_cycle = slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave & slow_peripheral_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module led_pio_s1_arbitrator (
                               // inputs:
                                clk,
                                led_pio_s1_readdata,
                                reset_n,
                                slow_peripheral_bridge_m1_address_to_slave,
                                slow_peripheral_bridge_m1_latency_counter,
                                slow_peripheral_bridge_m1_nativeaddress,
                                slow_peripheral_bridge_m1_read,
                                slow_peripheral_bridge_m1_write,
                                slow_peripheral_bridge_m1_writedata,

                               // outputs:
                                d1_led_pio_s1_end_xfer,
                                led_pio_s1_address,
                                led_pio_s1_chipselect,
                                led_pio_s1_readdata_from_sa,
                                led_pio_s1_reset_n,
                                led_pio_s1_write_n,
                                led_pio_s1_writedata,
                                slow_peripheral_bridge_m1_granted_led_pio_s1,
                                slow_peripheral_bridge_m1_qualified_request_led_pio_s1,
                                slow_peripheral_bridge_m1_read_data_valid_led_pio_s1,
                                slow_peripheral_bridge_m1_requests_led_pio_s1
                             )
;

  output           d1_led_pio_s1_end_xfer;
  output  [  1: 0] led_pio_s1_address;
  output           led_pio_s1_chipselect;
  output  [ 31: 0] led_pio_s1_readdata_from_sa;
  output           led_pio_s1_reset_n;
  output           led_pio_s1_write_n;
  output  [ 31: 0] led_pio_s1_writedata;
  output           slow_peripheral_bridge_m1_granted_led_pio_s1;
  output           slow_peripheral_bridge_m1_qualified_request_led_pio_s1;
  output           slow_peripheral_bridge_m1_read_data_valid_led_pio_s1;
  output           slow_peripheral_bridge_m1_requests_led_pio_s1;
  input            clk;
  input   [ 31: 0] led_pio_s1_readdata;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  input            slow_peripheral_bridge_m1_latency_counter;
  input   [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] slow_peripheral_bridge_m1_writedata;

  reg              d1_led_pio_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_led_pio_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] led_pio_s1_address;
  wire             led_pio_s1_allgrants;
  wire             led_pio_s1_allow_new_arb_cycle;
  wire             led_pio_s1_any_bursting_master_saved_grant;
  wire             led_pio_s1_any_continuerequest;
  wire             led_pio_s1_arb_counter_enable;
  reg              led_pio_s1_arb_share_counter;
  wire             led_pio_s1_arb_share_counter_next_value;
  wire             led_pio_s1_arb_share_set_values;
  wire             led_pio_s1_beginbursttransfer_internal;
  wire             led_pio_s1_begins_xfer;
  wire             led_pio_s1_chipselect;
  wire             led_pio_s1_end_xfer;
  wire             led_pio_s1_firsttransfer;
  wire             led_pio_s1_grant_vector;
  wire             led_pio_s1_in_a_read_cycle;
  wire             led_pio_s1_in_a_write_cycle;
  wire             led_pio_s1_master_qreq_vector;
  wire             led_pio_s1_non_bursting_master_requests;
  wire    [ 31: 0] led_pio_s1_readdata_from_sa;
  reg              led_pio_s1_reg_firsttransfer;
  wire             led_pio_s1_reset_n;
  reg              led_pio_s1_slavearbiterlockenable;
  wire             led_pio_s1_slavearbiterlockenable2;
  wire             led_pio_s1_unreg_firsttransfer;
  wire             led_pio_s1_waits_for_read;
  wire             led_pio_s1_waits_for_write;
  wire             led_pio_s1_write_n;
  wire    [ 31: 0] led_pio_s1_writedata;
  wire             slow_peripheral_bridge_m1_arbiterlock;
  wire             slow_peripheral_bridge_m1_arbiterlock2;
  wire             slow_peripheral_bridge_m1_continuerequest;
  wire             slow_peripheral_bridge_m1_granted_led_pio_s1;
  wire             slow_peripheral_bridge_m1_qualified_request_led_pio_s1;
  wire             slow_peripheral_bridge_m1_read_data_valid_led_pio_s1;
  wire             slow_peripheral_bridge_m1_requests_led_pio_s1;
  wire             slow_peripheral_bridge_m1_saved_grant_led_pio_s1;
  wire             wait_for_led_pio_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~led_pio_s1_end_xfer;
    end


  assign led_pio_s1_begins_xfer = ~d1_reasons_to_wait & ((slow_peripheral_bridge_m1_qualified_request_led_pio_s1));
  //assign led_pio_s1_readdata_from_sa = led_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign led_pio_s1_readdata_from_sa = led_pio_s1_readdata;

  assign slow_peripheral_bridge_m1_requests_led_pio_s1 = ({slow_peripheral_bridge_m1_address_to_slave[7 : 4] , 4'b0} == 8'hd0) & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write);
  //led_pio_s1_arb_share_counter set values, which is an e_mux
  assign led_pio_s1_arb_share_set_values = 1;

  //led_pio_s1_non_bursting_master_requests mux, which is an e_mux
  assign led_pio_s1_non_bursting_master_requests = slow_peripheral_bridge_m1_requests_led_pio_s1;

  //led_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign led_pio_s1_any_bursting_master_saved_grant = 0;

  //led_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign led_pio_s1_arb_share_counter_next_value = led_pio_s1_firsttransfer ? (led_pio_s1_arb_share_set_values - 1) : |led_pio_s1_arb_share_counter ? (led_pio_s1_arb_share_counter - 1) : 0;

  //led_pio_s1_allgrants all slave grants, which is an e_mux
  assign led_pio_s1_allgrants = |led_pio_s1_grant_vector;

  //led_pio_s1_end_xfer assignment, which is an e_assign
  assign led_pio_s1_end_xfer = ~(led_pio_s1_waits_for_read | led_pio_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_led_pio_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_led_pio_s1 = led_pio_s1_end_xfer & (~led_pio_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //led_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign led_pio_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_led_pio_s1 & led_pio_s1_allgrants) | (end_xfer_arb_share_counter_term_led_pio_s1 & ~led_pio_s1_non_bursting_master_requests);

  //led_pio_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          led_pio_s1_arb_share_counter <= 0;
      else if (led_pio_s1_arb_counter_enable)
          led_pio_s1_arb_share_counter <= led_pio_s1_arb_share_counter_next_value;
    end


  //led_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          led_pio_s1_slavearbiterlockenable <= 0;
      else if ((|led_pio_s1_master_qreq_vector & end_xfer_arb_share_counter_term_led_pio_s1) | (end_xfer_arb_share_counter_term_led_pio_s1 & ~led_pio_s1_non_bursting_master_requests))
          led_pio_s1_slavearbiterlockenable <= |led_pio_s1_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge/m1 led_pio/s1 arbiterlock, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock = led_pio_s1_slavearbiterlockenable & slow_peripheral_bridge_m1_continuerequest;

  //led_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign led_pio_s1_slavearbiterlockenable2 = |led_pio_s1_arb_share_counter_next_value;

  //slow_peripheral_bridge/m1 led_pio/s1 arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock2 = led_pio_s1_slavearbiterlockenable2 & slow_peripheral_bridge_m1_continuerequest;

  //led_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign led_pio_s1_any_continuerequest = 1;

  //slow_peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  assign slow_peripheral_bridge_m1_continuerequest = 1;

  assign slow_peripheral_bridge_m1_qualified_request_led_pio_s1 = slow_peripheral_bridge_m1_requests_led_pio_s1 & ~((slow_peripheral_bridge_m1_read & ((slow_peripheral_bridge_m1_latency_counter != 0))));
  //local readdatavalid slow_peripheral_bridge_m1_read_data_valid_led_pio_s1, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_led_pio_s1 = slow_peripheral_bridge_m1_granted_led_pio_s1 & slow_peripheral_bridge_m1_read & ~led_pio_s1_waits_for_read;

  //led_pio_s1_writedata mux, which is an e_mux
  assign led_pio_s1_writedata = slow_peripheral_bridge_m1_writedata;

  //master is always granted when requested
  assign slow_peripheral_bridge_m1_granted_led_pio_s1 = slow_peripheral_bridge_m1_qualified_request_led_pio_s1;

  //slow_peripheral_bridge/m1 saved-grant led_pio/s1, which is an e_assign
  assign slow_peripheral_bridge_m1_saved_grant_led_pio_s1 = slow_peripheral_bridge_m1_requests_led_pio_s1;

  //allow new arb cycle for led_pio/s1, which is an e_assign
  assign led_pio_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign led_pio_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign led_pio_s1_master_qreq_vector = 1;

  //led_pio_s1_reset_n assignment, which is an e_assign
  assign led_pio_s1_reset_n = reset_n;

  assign led_pio_s1_chipselect = slow_peripheral_bridge_m1_granted_led_pio_s1;
  //led_pio_s1_firsttransfer first transaction, which is an e_assign
  assign led_pio_s1_firsttransfer = led_pio_s1_begins_xfer ? led_pio_s1_unreg_firsttransfer : led_pio_s1_reg_firsttransfer;

  //led_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign led_pio_s1_unreg_firsttransfer = ~(led_pio_s1_slavearbiterlockenable & led_pio_s1_any_continuerequest);

  //led_pio_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          led_pio_s1_reg_firsttransfer <= 1'b1;
      else if (led_pio_s1_begins_xfer)
          led_pio_s1_reg_firsttransfer <= led_pio_s1_unreg_firsttransfer;
    end


  //led_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign led_pio_s1_beginbursttransfer_internal = led_pio_s1_begins_xfer;

  //~led_pio_s1_write_n assignment, which is an e_mux
  assign led_pio_s1_write_n = ~(slow_peripheral_bridge_m1_granted_led_pio_s1 & slow_peripheral_bridge_m1_write);

  //led_pio_s1_address mux, which is an e_mux
  assign led_pio_s1_address = slow_peripheral_bridge_m1_nativeaddress;

  //d1_led_pio_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_led_pio_s1_end_xfer <= 1;
      else 
        d1_led_pio_s1_end_xfer <= led_pio_s1_end_xfer;
    end


  //led_pio_s1_waits_for_read in a cycle, which is an e_mux
  assign led_pio_s1_waits_for_read = led_pio_s1_in_a_read_cycle & led_pio_s1_begins_xfer;

  //led_pio_s1_in_a_read_cycle assignment, which is an e_assign
  assign led_pio_s1_in_a_read_cycle = slow_peripheral_bridge_m1_granted_led_pio_s1 & slow_peripheral_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = led_pio_s1_in_a_read_cycle;

  //led_pio_s1_waits_for_write in a cycle, which is an e_mux
  assign led_pio_s1_waits_for_write = led_pio_s1_in_a_write_cycle & 0;

  //led_pio_s1_in_a_write_cycle assignment, which is an e_assign
  assign led_pio_s1_in_a_write_cycle = slow_peripheral_bridge_m1_granted_led_pio_s1 & slow_peripheral_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = led_pio_s1_in_a_write_cycle;

  assign wait_for_led_pio_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //led_pio/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module performance_counter_control_slave_arbitrator (
                                                      // inputs:
                                                       clk,
                                                       performance_counter_control_slave_readdata,
                                                       reset_n,
                                                       slow_peripheral_bridge_m1_address_to_slave,
                                                       slow_peripheral_bridge_m1_latency_counter,
                                                       slow_peripheral_bridge_m1_nativeaddress,
                                                       slow_peripheral_bridge_m1_read,
                                                       slow_peripheral_bridge_m1_write,
                                                       slow_peripheral_bridge_m1_writedata,

                                                      // outputs:
                                                       d1_performance_counter_control_slave_end_xfer,
                                                       performance_counter_control_slave_address,
                                                       performance_counter_control_slave_begintransfer,
                                                       performance_counter_control_slave_readdata_from_sa,
                                                       performance_counter_control_slave_reset_n,
                                                       performance_counter_control_slave_write,
                                                       performance_counter_control_slave_writedata,
                                                       slow_peripheral_bridge_m1_granted_performance_counter_control_slave,
                                                       slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave,
                                                       slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave,
                                                       slow_peripheral_bridge_m1_requests_performance_counter_control_slave
                                                    )
;

  output           d1_performance_counter_control_slave_end_xfer;
  output  [  2: 0] performance_counter_control_slave_address;
  output           performance_counter_control_slave_begintransfer;
  output  [ 31: 0] performance_counter_control_slave_readdata_from_sa;
  output           performance_counter_control_slave_reset_n;
  output           performance_counter_control_slave_write;
  output  [ 31: 0] performance_counter_control_slave_writedata;
  output           slow_peripheral_bridge_m1_granted_performance_counter_control_slave;
  output           slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave;
  output           slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave;
  output           slow_peripheral_bridge_m1_requests_performance_counter_control_slave;
  input            clk;
  input   [ 31: 0] performance_counter_control_slave_readdata;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  input            slow_peripheral_bridge_m1_latency_counter;
  input   [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] slow_peripheral_bridge_m1_writedata;

  reg              d1_performance_counter_control_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_performance_counter_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p1_slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register;
  wire    [  2: 0] performance_counter_control_slave_address;
  wire             performance_counter_control_slave_allgrants;
  wire             performance_counter_control_slave_allow_new_arb_cycle;
  wire             performance_counter_control_slave_any_bursting_master_saved_grant;
  wire             performance_counter_control_slave_any_continuerequest;
  wire             performance_counter_control_slave_arb_counter_enable;
  reg              performance_counter_control_slave_arb_share_counter;
  wire             performance_counter_control_slave_arb_share_counter_next_value;
  wire             performance_counter_control_slave_arb_share_set_values;
  wire             performance_counter_control_slave_beginbursttransfer_internal;
  wire             performance_counter_control_slave_begins_xfer;
  wire             performance_counter_control_slave_begintransfer;
  wire             performance_counter_control_slave_end_xfer;
  wire             performance_counter_control_slave_firsttransfer;
  wire             performance_counter_control_slave_grant_vector;
  wire             performance_counter_control_slave_in_a_read_cycle;
  wire             performance_counter_control_slave_in_a_write_cycle;
  wire             performance_counter_control_slave_master_qreq_vector;
  wire             performance_counter_control_slave_non_bursting_master_requests;
  wire    [ 31: 0] performance_counter_control_slave_readdata_from_sa;
  reg              performance_counter_control_slave_reg_firsttransfer;
  wire             performance_counter_control_slave_reset_n;
  reg              performance_counter_control_slave_slavearbiterlockenable;
  wire             performance_counter_control_slave_slavearbiterlockenable2;
  wire             performance_counter_control_slave_unreg_firsttransfer;
  wire             performance_counter_control_slave_waits_for_read;
  wire             performance_counter_control_slave_waits_for_write;
  wire             performance_counter_control_slave_write;
  wire    [ 31: 0] performance_counter_control_slave_writedata;
  wire             slow_peripheral_bridge_m1_arbiterlock;
  wire             slow_peripheral_bridge_m1_arbiterlock2;
  wire             slow_peripheral_bridge_m1_continuerequest;
  wire             slow_peripheral_bridge_m1_granted_performance_counter_control_slave;
  wire             slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave;
  wire             slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave;
  reg              slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register;
  wire             slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register_in;
  wire             slow_peripheral_bridge_m1_requests_performance_counter_control_slave;
  wire             slow_peripheral_bridge_m1_saved_grant_performance_counter_control_slave;
  wire             wait_for_performance_counter_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~performance_counter_control_slave_end_xfer;
    end


  assign performance_counter_control_slave_begins_xfer = ~d1_reasons_to_wait & ((slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave));
  //assign performance_counter_control_slave_readdata_from_sa = performance_counter_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign performance_counter_control_slave_readdata_from_sa = performance_counter_control_slave_readdata;

  assign slow_peripheral_bridge_m1_requests_performance_counter_control_slave = ({slow_peripheral_bridge_m1_address_to_slave[7 : 5] , 5'b0} == 8'h20) & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write);
  //performance_counter_control_slave_arb_share_counter set values, which is an e_mux
  assign performance_counter_control_slave_arb_share_set_values = 1;

  //performance_counter_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign performance_counter_control_slave_non_bursting_master_requests = slow_peripheral_bridge_m1_requests_performance_counter_control_slave;

  //performance_counter_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign performance_counter_control_slave_any_bursting_master_saved_grant = 0;

  //performance_counter_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign performance_counter_control_slave_arb_share_counter_next_value = performance_counter_control_slave_firsttransfer ? (performance_counter_control_slave_arb_share_set_values - 1) : |performance_counter_control_slave_arb_share_counter ? (performance_counter_control_slave_arb_share_counter - 1) : 0;

  //performance_counter_control_slave_allgrants all slave grants, which is an e_mux
  assign performance_counter_control_slave_allgrants = |performance_counter_control_slave_grant_vector;

  //performance_counter_control_slave_end_xfer assignment, which is an e_assign
  assign performance_counter_control_slave_end_xfer = ~(performance_counter_control_slave_waits_for_read | performance_counter_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_performance_counter_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_performance_counter_control_slave = performance_counter_control_slave_end_xfer & (~performance_counter_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //performance_counter_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign performance_counter_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_performance_counter_control_slave & performance_counter_control_slave_allgrants) | (end_xfer_arb_share_counter_term_performance_counter_control_slave & ~performance_counter_control_slave_non_bursting_master_requests);

  //performance_counter_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          performance_counter_control_slave_arb_share_counter <= 0;
      else if (performance_counter_control_slave_arb_counter_enable)
          performance_counter_control_slave_arb_share_counter <= performance_counter_control_slave_arb_share_counter_next_value;
    end


  //performance_counter_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          performance_counter_control_slave_slavearbiterlockenable <= 0;
      else if ((|performance_counter_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_performance_counter_control_slave) | (end_xfer_arb_share_counter_term_performance_counter_control_slave & ~performance_counter_control_slave_non_bursting_master_requests))
          performance_counter_control_slave_slavearbiterlockenable <= |performance_counter_control_slave_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge/m1 performance_counter/control_slave arbiterlock, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock = performance_counter_control_slave_slavearbiterlockenable & slow_peripheral_bridge_m1_continuerequest;

  //performance_counter_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign performance_counter_control_slave_slavearbiterlockenable2 = |performance_counter_control_slave_arb_share_counter_next_value;

  //slow_peripheral_bridge/m1 performance_counter/control_slave arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock2 = performance_counter_control_slave_slavearbiterlockenable2 & slow_peripheral_bridge_m1_continuerequest;

  //performance_counter_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign performance_counter_control_slave_any_continuerequest = 1;

  //slow_peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  assign slow_peripheral_bridge_m1_continuerequest = 1;

  assign slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave = slow_peripheral_bridge_m1_requests_performance_counter_control_slave & ~((slow_peripheral_bridge_m1_read & ((1 < slow_peripheral_bridge_m1_latency_counter))));
  //slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register_in = slow_peripheral_bridge_m1_granted_performance_counter_control_slave & slow_peripheral_bridge_m1_read & ~performance_counter_control_slave_waits_for_read;

  //shift register p1 slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register = {slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register, slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register_in};

  //slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register <= 0;
      else 
        slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register <= p1_slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register;
    end


  //local readdatavalid slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave = slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave_shift_register;

  //performance_counter_control_slave_writedata mux, which is an e_mux
  assign performance_counter_control_slave_writedata = slow_peripheral_bridge_m1_writedata;

  //master is always granted when requested
  assign slow_peripheral_bridge_m1_granted_performance_counter_control_slave = slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave;

  //slow_peripheral_bridge/m1 saved-grant performance_counter/control_slave, which is an e_assign
  assign slow_peripheral_bridge_m1_saved_grant_performance_counter_control_slave = slow_peripheral_bridge_m1_requests_performance_counter_control_slave;

  //allow new arb cycle for performance_counter/control_slave, which is an e_assign
  assign performance_counter_control_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign performance_counter_control_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign performance_counter_control_slave_master_qreq_vector = 1;

  assign performance_counter_control_slave_begintransfer = performance_counter_control_slave_begins_xfer;
  //performance_counter_control_slave_reset_n assignment, which is an e_assign
  assign performance_counter_control_slave_reset_n = reset_n;

  //performance_counter_control_slave_firsttransfer first transaction, which is an e_assign
  assign performance_counter_control_slave_firsttransfer = performance_counter_control_slave_begins_xfer ? performance_counter_control_slave_unreg_firsttransfer : performance_counter_control_slave_reg_firsttransfer;

  //performance_counter_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign performance_counter_control_slave_unreg_firsttransfer = ~(performance_counter_control_slave_slavearbiterlockenable & performance_counter_control_slave_any_continuerequest);

  //performance_counter_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          performance_counter_control_slave_reg_firsttransfer <= 1'b1;
      else if (performance_counter_control_slave_begins_xfer)
          performance_counter_control_slave_reg_firsttransfer <= performance_counter_control_slave_unreg_firsttransfer;
    end


  //performance_counter_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign performance_counter_control_slave_beginbursttransfer_internal = performance_counter_control_slave_begins_xfer;

  //performance_counter_control_slave_write assignment, which is an e_mux
  assign performance_counter_control_slave_write = slow_peripheral_bridge_m1_granted_performance_counter_control_slave & slow_peripheral_bridge_m1_write;

  //performance_counter_control_slave_address mux, which is an e_mux
  assign performance_counter_control_slave_address = slow_peripheral_bridge_m1_nativeaddress;

  //d1_performance_counter_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_performance_counter_control_slave_end_xfer <= 1;
      else 
        d1_performance_counter_control_slave_end_xfer <= performance_counter_control_slave_end_xfer;
    end


  //performance_counter_control_slave_waits_for_read in a cycle, which is an e_mux
  assign performance_counter_control_slave_waits_for_read = performance_counter_control_slave_in_a_read_cycle & 0;

  //performance_counter_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign performance_counter_control_slave_in_a_read_cycle = slow_peripheral_bridge_m1_granted_performance_counter_control_slave & slow_peripheral_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = performance_counter_control_slave_in_a_read_cycle;

  //performance_counter_control_slave_waits_for_write in a cycle, which is an e_mux
  assign performance_counter_control_slave_waits_for_write = performance_counter_control_slave_in_a_write_cycle & 0;

  //performance_counter_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign performance_counter_control_slave_in_a_write_cycle = slow_peripheral_bridge_m1_granted_performance_counter_control_slave & slow_peripheral_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = performance_counter_control_slave_in_a_write_cycle;

  assign wait_for_performance_counter_control_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //performance_counter/control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_pipeline_bridge_before_tristate_bridge_s1_module (
                                                                                          // inputs:
                                                                                           clear_fifo,
                                                                                           clk,
                                                                                           data_in,
                                                                                           read,
                                                                                           reset_n,
                                                                                           sync_reset,
                                                                                           write,

                                                                                          // outputs:
                                                                                           data_out,
                                                                                           empty,
                                                                                           fifo_contains_ones_n,
                                                                                           full
                                                                                        )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  wire             full_5;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_4;
  assign empty = !full_0;
  assign full_5 = 0;
  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    0;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_before_tristate_bridge_s1_module (
                                                                                                 // inputs:
                                                                                                  clear_fifo,
                                                                                                  clk,
                                                                                                  data_in,
                                                                                                  read,
                                                                                                  reset_n,
                                                                                                  sync_reset,
                                                                                                  write,

                                                                                                 // outputs:
                                                                                                  data_out,
                                                                                                  empty,
                                                                                                  fifo_contains_ones_n,
                                                                                                  full
                                                                                               )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  wire             full_5;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_4;
  assign empty = !full_0;
  assign full_5 = 0;
  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    0;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_before_tristate_bridge_s1_arbitrator (
                                                              // inputs:
                                                               clk,
                                                               cpu_data_master_address_to_slave,
                                                               cpu_data_master_byteenable,
                                                               cpu_data_master_debugaccess,
                                                               cpu_data_master_latency_counter,
                                                               cpu_data_master_read,
                                                               cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                                               cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register,
                                                               cpu_data_master_write,
                                                               cpu_data_master_writedata,
                                                               cpu_instruction_master_address_to_slave,
                                                               cpu_instruction_master_latency_counter,
                                                               cpu_instruction_master_read,
                                                               cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                                               pipeline_bridge_before_tristate_bridge_s1_endofpacket,
                                                               pipeline_bridge_before_tristate_bridge_s1_readdata,
                                                               pipeline_bridge_before_tristate_bridge_s1_readdatavalid,
                                                               pipeline_bridge_before_tristate_bridge_s1_waitrequest,
                                                               reset_n,

                                                              // outputs:
                                                               cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1,
                                                               cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1,
                                                               cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1,
                                                               cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                                               cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1,
                                                               cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1,
                                                               cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1,
                                                               cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1,
                                                               cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                                               cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1,
                                                               d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer,
                                                               pipeline_bridge_before_tristate_bridge_s1_address,
                                                               pipeline_bridge_before_tristate_bridge_s1_arbiterlock,
                                                               pipeline_bridge_before_tristate_bridge_s1_arbiterlock2,
                                                               pipeline_bridge_before_tristate_bridge_s1_burstcount,
                                                               pipeline_bridge_before_tristate_bridge_s1_byteenable,
                                                               pipeline_bridge_before_tristate_bridge_s1_chipselect,
                                                               pipeline_bridge_before_tristate_bridge_s1_debugaccess,
                                                               pipeline_bridge_before_tristate_bridge_s1_endofpacket_from_sa,
                                                               pipeline_bridge_before_tristate_bridge_s1_nativeaddress,
                                                               pipeline_bridge_before_tristate_bridge_s1_read,
                                                               pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa,
                                                               pipeline_bridge_before_tristate_bridge_s1_reset_n,
                                                               pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa,
                                                               pipeline_bridge_before_tristate_bridge_s1_write,
                                                               pipeline_bridge_before_tristate_bridge_s1_writedata
                                                            )
;

  output           cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1;
  output           cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1;
  output           cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1;
  output           cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  output           cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1;
  output           cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1;
  output           cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1;
  output           cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1;
  output           cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  output           cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1;
  output           d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer;
  output  [ 24: 0] pipeline_bridge_before_tristate_bridge_s1_address;
  output           pipeline_bridge_before_tristate_bridge_s1_arbiterlock;
  output           pipeline_bridge_before_tristate_bridge_s1_arbiterlock2;
  output           pipeline_bridge_before_tristate_bridge_s1_burstcount;
  output  [  3: 0] pipeline_bridge_before_tristate_bridge_s1_byteenable;
  output           pipeline_bridge_before_tristate_bridge_s1_chipselect;
  output           pipeline_bridge_before_tristate_bridge_s1_debugaccess;
  output           pipeline_bridge_before_tristate_bridge_s1_endofpacket_from_sa;
  output  [ 24: 0] pipeline_bridge_before_tristate_bridge_s1_nativeaddress;
  output           pipeline_bridge_before_tristate_bridge_s1_read;
  output  [ 31: 0] pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa;
  output           pipeline_bridge_before_tristate_bridge_s1_reset_n;
  output           pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa;
  output           pipeline_bridge_before_tristate_bridge_s1_write;
  output  [ 31: 0] pipeline_bridge_before_tristate_bridge_s1_writedata;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 28: 0] cpu_instruction_master_address_to_slave;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            pipeline_bridge_before_tristate_bridge_s1_endofpacket;
  input   [ 31: 0] pipeline_bridge_before_tristate_bridge_s1_readdata;
  input            pipeline_bridge_before_tristate_bridge_s1_readdatavalid;
  input            pipeline_bridge_before_tristate_bridge_s1_waitrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_data_master_rdv_fifo_empty_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_data_master_rdv_fifo_output_from_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  wire             cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_data_master_saved_grant_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_rdv_fifo_output_from_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  wire             cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_saved_grant_pipeline_bridge_before_tristate_bridge_s1;
  reg              d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_bridge_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_data_master_granted_slave_pipeline_bridge_before_tristate_bridge_s1;
  reg              last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_before_tristate_bridge_s1;
  wire    [ 24: 0] pipeline_bridge_before_tristate_bridge_s1_address;
  wire             pipeline_bridge_before_tristate_bridge_s1_allgrants;
  wire             pipeline_bridge_before_tristate_bridge_s1_allow_new_arb_cycle;
  wire             pipeline_bridge_before_tristate_bridge_s1_any_bursting_master_saved_grant;
  wire             pipeline_bridge_before_tristate_bridge_s1_any_continuerequest;
  reg     [  1: 0] pipeline_bridge_before_tristate_bridge_s1_arb_addend;
  wire             pipeline_bridge_before_tristate_bridge_s1_arb_counter_enable;
  reg              pipeline_bridge_before_tristate_bridge_s1_arb_share_counter;
  wire             pipeline_bridge_before_tristate_bridge_s1_arb_share_counter_next_value;
  wire             pipeline_bridge_before_tristate_bridge_s1_arb_share_set_values;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_s1_arb_winner;
  wire             pipeline_bridge_before_tristate_bridge_s1_arbiterlock;
  wire             pipeline_bridge_before_tristate_bridge_s1_arbiterlock2;
  wire             pipeline_bridge_before_tristate_bridge_s1_arbitration_holdoff_internal;
  wire             pipeline_bridge_before_tristate_bridge_s1_beginbursttransfer_internal;
  wire             pipeline_bridge_before_tristate_bridge_s1_begins_xfer;
  wire             pipeline_bridge_before_tristate_bridge_s1_burstcount;
  wire    [  3: 0] pipeline_bridge_before_tristate_bridge_s1_byteenable;
  wire             pipeline_bridge_before_tristate_bridge_s1_chipselect;
  wire    [  3: 0] pipeline_bridge_before_tristate_bridge_s1_chosen_master_double_vector;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_s1_chosen_master_rot_left;
  wire             pipeline_bridge_before_tristate_bridge_s1_debugaccess;
  wire             pipeline_bridge_before_tristate_bridge_s1_end_xfer;
  wire             pipeline_bridge_before_tristate_bridge_s1_endofpacket_from_sa;
  wire             pipeline_bridge_before_tristate_bridge_s1_firsttransfer;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_s1_grant_vector;
  wire             pipeline_bridge_before_tristate_bridge_s1_in_a_read_cycle;
  wire             pipeline_bridge_before_tristate_bridge_s1_in_a_write_cycle;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_s1_master_qreq_vector;
  wire             pipeline_bridge_before_tristate_bridge_s1_move_on_to_next_transaction;
  wire    [ 24: 0] pipeline_bridge_before_tristate_bridge_s1_nativeaddress;
  wire             pipeline_bridge_before_tristate_bridge_s1_non_bursting_master_requests;
  wire             pipeline_bridge_before_tristate_bridge_s1_read;
  wire    [ 31: 0] pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa;
  wire             pipeline_bridge_before_tristate_bridge_s1_readdatavalid_from_sa;
  reg              pipeline_bridge_before_tristate_bridge_s1_reg_firsttransfer;
  wire             pipeline_bridge_before_tristate_bridge_s1_reset_n;
  reg     [  1: 0] pipeline_bridge_before_tristate_bridge_s1_saved_chosen_master_vector;
  reg              pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable;
  wire             pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable2;
  wire             pipeline_bridge_before_tristate_bridge_s1_unreg_firsttransfer;
  wire             pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa;
  wire             pipeline_bridge_before_tristate_bridge_s1_waits_for_read;
  wire             pipeline_bridge_before_tristate_bridge_s1_waits_for_write;
  wire             pipeline_bridge_before_tristate_bridge_s1_write;
  wire    [ 31: 0] pipeline_bridge_before_tristate_bridge_s1_writedata;
  wire    [ 28: 0] shifted_address_to_pipeline_bridge_before_tristate_bridge_s1_from_cpu_data_master;
  wire    [ 28: 0] shifted_address_to_pipeline_bridge_before_tristate_bridge_s1_from_cpu_instruction_master;
  wire             wait_for_pipeline_bridge_before_tristate_bridge_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pipeline_bridge_before_tristate_bridge_s1_end_xfer;
    end


  assign pipeline_bridge_before_tristate_bridge_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1 | cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1));
  //assign pipeline_bridge_before_tristate_bridge_s1_readdatavalid_from_sa = pipeline_bridge_before_tristate_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_readdatavalid_from_sa = pipeline_bridge_before_tristate_bridge_s1_readdatavalid;

  //assign pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa = pipeline_bridge_before_tristate_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa = pipeline_bridge_before_tristate_bridge_s1_readdata;

  assign cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1 = ({cpu_data_master_address_to_slave[28 : 27] , 27'b0} == 29'h10000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa = pipeline_bridge_before_tristate_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa = pipeline_bridge_before_tristate_bridge_s1_waitrequest;

  //pipeline_bridge_before_tristate_bridge_s1_arb_share_counter set values, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_arb_share_set_values = 1;

  //pipeline_bridge_before_tristate_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_non_bursting_master_requests = cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1 |
    cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1 |
    cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1 |
    cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1 |
    cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1 |
    cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1;

  //pipeline_bridge_before_tristate_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_any_bursting_master_saved_grant = 0;

  //pipeline_bridge_before_tristate_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_arb_share_counter_next_value = pipeline_bridge_before_tristate_bridge_s1_firsttransfer ? (pipeline_bridge_before_tristate_bridge_s1_arb_share_set_values - 1) : |pipeline_bridge_before_tristate_bridge_s1_arb_share_counter ? (pipeline_bridge_before_tristate_bridge_s1_arb_share_counter - 1) : 0;

  //pipeline_bridge_before_tristate_bridge_s1_allgrants all slave grants, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_allgrants = (|pipeline_bridge_before_tristate_bridge_s1_grant_vector) |
    (|pipeline_bridge_before_tristate_bridge_s1_grant_vector) |
    (|pipeline_bridge_before_tristate_bridge_s1_grant_vector) |
    (|pipeline_bridge_before_tristate_bridge_s1_grant_vector) |
    (|pipeline_bridge_before_tristate_bridge_s1_grant_vector) |
    (|pipeline_bridge_before_tristate_bridge_s1_grant_vector);

  //pipeline_bridge_before_tristate_bridge_s1_end_xfer assignment, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_end_xfer = ~(pipeline_bridge_before_tristate_bridge_s1_waits_for_read | pipeline_bridge_before_tristate_bridge_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_bridge_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_bridge_s1 = pipeline_bridge_before_tristate_bridge_s1_end_xfer & (~pipeline_bridge_before_tristate_bridge_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pipeline_bridge_before_tristate_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_bridge_s1 & pipeline_bridge_before_tristate_bridge_s1_allgrants) | (end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_bridge_s1 & ~pipeline_bridge_before_tristate_bridge_s1_non_bursting_master_requests);

  //pipeline_bridge_before_tristate_bridge_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_s1_arb_share_counter <= 0;
      else if (pipeline_bridge_before_tristate_bridge_s1_arb_counter_enable)
          pipeline_bridge_before_tristate_bridge_s1_arb_share_counter <= pipeline_bridge_before_tristate_bridge_s1_arb_share_counter_next_value;
    end


  //pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable <= 0;
      else if ((|pipeline_bridge_before_tristate_bridge_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_bridge_s1) | (end_xfer_arb_share_counter_term_pipeline_bridge_before_tristate_bridge_s1 & ~pipeline_bridge_before_tristate_bridge_s1_non_bursting_master_requests))
          pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable <= |pipeline_bridge_before_tristate_bridge_s1_arb_share_counter_next_value;
    end


  //cpu/data_master pipeline_bridge_before_tristate_bridge/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable2 = |pipeline_bridge_before_tristate_bridge_s1_arb_share_counter_next_value;

  //cpu/data_master pipeline_bridge_before_tristate_bridge/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //cpu/instruction_master pipeline_bridge_before_tristate_bridge/s1 arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //cpu/instruction_master pipeline_bridge_before_tristate_bridge/s1 arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //cpu/instruction_master granted pipeline_bridge_before_tristate_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_before_tristate_bridge_s1 <= 0;
      else 
        last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_before_tristate_bridge_s1 <= cpu_instruction_master_saved_grant_pipeline_bridge_before_tristate_bridge_s1 ? 1 : (pipeline_bridge_before_tristate_bridge_s1_arbitration_holdoff_internal | ~cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1) ? 0 : last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_before_tristate_bridge_s1;
    end


  //cpu_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_instruction_master_continuerequest = last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_before_tristate_bridge_s1 & cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1;

  //pipeline_bridge_before_tristate_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_any_continuerequest = cpu_instruction_master_continuerequest |
    cpu_data_master_continuerequest;

  assign cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1 = cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register))) | cpu_instruction_master_arbiterlock);
  //unique name for pipeline_bridge_before_tristate_bridge_s1_move_on_to_next_transaction, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_move_on_to_next_transaction = pipeline_bridge_before_tristate_bridge_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_pipeline_bridge_before_tristate_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_pipeline_bridge_before_tristate_bridge_s1_module rdv_fifo_for_cpu_data_master_to_pipeline_bridge_before_tristate_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1),
      .data_out             (cpu_data_master_rdv_fifo_output_from_pipeline_bridge_before_tristate_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_pipeline_bridge_before_tristate_bridge_s1),
      .full                 (),
      .read                 (pipeline_bridge_before_tristate_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pipeline_bridge_before_tristate_bridge_s1_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register = ~cpu_data_master_rdv_fifo_empty_pipeline_bridge_before_tristate_bridge_s1;
  //local readdatavalid cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1 = (pipeline_bridge_before_tristate_bridge_s1_readdatavalid_from_sa & cpu_data_master_rdv_fifo_output_from_pipeline_bridge_before_tristate_bridge_s1) & ~ cpu_data_master_rdv_fifo_empty_pipeline_bridge_before_tristate_bridge_s1;

  //pipeline_bridge_before_tristate_bridge_s1_writedata mux, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_writedata = cpu_data_master_writedata;

  //assign pipeline_bridge_before_tristate_bridge_s1_endofpacket_from_sa = pipeline_bridge_before_tristate_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_endofpacket_from_sa = pipeline_bridge_before_tristate_bridge_s1_endofpacket;

  assign cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1 = (({cpu_instruction_master_address_to_slave[28 : 27] , 27'b0} == 29'h10000000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //cpu/data_master granted pipeline_bridge_before_tristate_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_data_master_granted_slave_pipeline_bridge_before_tristate_bridge_s1 <= 0;
      else 
        last_cycle_cpu_data_master_granted_slave_pipeline_bridge_before_tristate_bridge_s1 <= cpu_data_master_saved_grant_pipeline_bridge_before_tristate_bridge_s1 ? 1 : (pipeline_bridge_before_tristate_bridge_s1_arbitration_holdoff_internal | ~cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1) ? 0 : last_cycle_cpu_data_master_granted_slave_pipeline_bridge_before_tristate_bridge_s1;
    end


  //cpu_data_master_continuerequest continued request, which is an e_mux
  assign cpu_data_master_continuerequest = last_cycle_cpu_data_master_granted_slave_pipeline_bridge_before_tristate_bridge_s1 & cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1;

  assign cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1 = cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1 & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register))) | cpu_data_master_arbiterlock);
  //rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_before_tristate_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_before_tristate_bridge_s1_module rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_before_tristate_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_pipeline_bridge_before_tristate_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_before_tristate_bridge_s1),
      .full                 (),
      .read                 (pipeline_bridge_before_tristate_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pipeline_bridge_before_tristate_bridge_s1_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register = ~cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_before_tristate_bridge_s1;
  //local readdatavalid cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1, which is an e_mux
  assign cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1 = (pipeline_bridge_before_tristate_bridge_s1_readdatavalid_from_sa & cpu_instruction_master_rdv_fifo_output_from_pipeline_bridge_before_tristate_bridge_s1) & ~ cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_before_tristate_bridge_s1;

  //allow new arb cycle for pipeline_bridge_before_tristate_bridge/s1, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_allow_new_arb_cycle = ~cpu_data_master_arbiterlock & ~cpu_instruction_master_arbiterlock;

  //cpu/instruction_master assignment into master qualified-requests vector for pipeline_bridge_before_tristate_bridge/s1, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_master_qreq_vector[0] = cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1;

  //cpu/instruction_master grant pipeline_bridge_before_tristate_bridge/s1, which is an e_assign
  assign cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1 = pipeline_bridge_before_tristate_bridge_s1_grant_vector[0];

  //cpu/instruction_master saved-grant pipeline_bridge_before_tristate_bridge/s1, which is an e_assign
  assign cpu_instruction_master_saved_grant_pipeline_bridge_before_tristate_bridge_s1 = pipeline_bridge_before_tristate_bridge_s1_arb_winner[0] && cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1;

  //cpu/data_master assignment into master qualified-requests vector for pipeline_bridge_before_tristate_bridge/s1, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_master_qreq_vector[1] = cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1;

  //cpu/data_master grant pipeline_bridge_before_tristate_bridge/s1, which is an e_assign
  assign cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1 = pipeline_bridge_before_tristate_bridge_s1_grant_vector[1];

  //cpu/data_master saved-grant pipeline_bridge_before_tristate_bridge/s1, which is an e_assign
  assign cpu_data_master_saved_grant_pipeline_bridge_before_tristate_bridge_s1 = pipeline_bridge_before_tristate_bridge_s1_arb_winner[1] && cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1;

  //pipeline_bridge_before_tristate_bridge/s1 chosen-master double-vector, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_chosen_master_double_vector = {pipeline_bridge_before_tristate_bridge_s1_master_qreq_vector, pipeline_bridge_before_tristate_bridge_s1_master_qreq_vector} & ({~pipeline_bridge_before_tristate_bridge_s1_master_qreq_vector, ~pipeline_bridge_before_tristate_bridge_s1_master_qreq_vector} + pipeline_bridge_before_tristate_bridge_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign pipeline_bridge_before_tristate_bridge_s1_arb_winner = (pipeline_bridge_before_tristate_bridge_s1_allow_new_arb_cycle & | pipeline_bridge_before_tristate_bridge_s1_grant_vector) ? pipeline_bridge_before_tristate_bridge_s1_grant_vector : pipeline_bridge_before_tristate_bridge_s1_saved_chosen_master_vector;

  //saved pipeline_bridge_before_tristate_bridge_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_s1_saved_chosen_master_vector <= 0;
      else if (pipeline_bridge_before_tristate_bridge_s1_allow_new_arb_cycle)
          pipeline_bridge_before_tristate_bridge_s1_saved_chosen_master_vector <= |pipeline_bridge_before_tristate_bridge_s1_grant_vector ? pipeline_bridge_before_tristate_bridge_s1_grant_vector : pipeline_bridge_before_tristate_bridge_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign pipeline_bridge_before_tristate_bridge_s1_grant_vector = {(pipeline_bridge_before_tristate_bridge_s1_chosen_master_double_vector[1] | pipeline_bridge_before_tristate_bridge_s1_chosen_master_double_vector[3]),
    (pipeline_bridge_before_tristate_bridge_s1_chosen_master_double_vector[0] | pipeline_bridge_before_tristate_bridge_s1_chosen_master_double_vector[2])};

  //pipeline_bridge_before_tristate_bridge/s1 chosen master rotated left, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_chosen_master_rot_left = (pipeline_bridge_before_tristate_bridge_s1_arb_winner << 1) ? (pipeline_bridge_before_tristate_bridge_s1_arb_winner << 1) : 1;

  //pipeline_bridge_before_tristate_bridge/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_s1_arb_addend <= 1;
      else if (|pipeline_bridge_before_tristate_bridge_s1_grant_vector)
          pipeline_bridge_before_tristate_bridge_s1_arb_addend <= pipeline_bridge_before_tristate_bridge_s1_end_xfer? pipeline_bridge_before_tristate_bridge_s1_chosen_master_rot_left : pipeline_bridge_before_tristate_bridge_s1_grant_vector;
    end


  //pipeline_bridge_before_tristate_bridge_s1_reset_n assignment, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_reset_n = reset_n;

  assign pipeline_bridge_before_tristate_bridge_s1_chipselect = cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1 | cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1;
  //pipeline_bridge_before_tristate_bridge_s1_firsttransfer first transaction, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_firsttransfer = pipeline_bridge_before_tristate_bridge_s1_begins_xfer ? pipeline_bridge_before_tristate_bridge_s1_unreg_firsttransfer : pipeline_bridge_before_tristate_bridge_s1_reg_firsttransfer;

  //pipeline_bridge_before_tristate_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_unreg_firsttransfer = ~(pipeline_bridge_before_tristate_bridge_s1_slavearbiterlockenable & pipeline_bridge_before_tristate_bridge_s1_any_continuerequest);

  //pipeline_bridge_before_tristate_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_s1_reg_firsttransfer <= 1'b1;
      else if (pipeline_bridge_before_tristate_bridge_s1_begins_xfer)
          pipeline_bridge_before_tristate_bridge_s1_reg_firsttransfer <= pipeline_bridge_before_tristate_bridge_s1_unreg_firsttransfer;
    end


  //pipeline_bridge_before_tristate_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_beginbursttransfer_internal = pipeline_bridge_before_tristate_bridge_s1_begins_xfer;

  //pipeline_bridge_before_tristate_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_arbitration_holdoff_internal = pipeline_bridge_before_tristate_bridge_s1_begins_xfer & pipeline_bridge_before_tristate_bridge_s1_firsttransfer;

  //pipeline_bridge_before_tristate_bridge_s1_read assignment, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_read = (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1 & cpu_instruction_master_read);

  //pipeline_bridge_before_tristate_bridge_s1_write assignment, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_write = cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1 & cpu_data_master_write;

  assign shifted_address_to_pipeline_bridge_before_tristate_bridge_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //pipeline_bridge_before_tristate_bridge_s1_address mux, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_address = (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1)? (shifted_address_to_pipeline_bridge_before_tristate_bridge_s1_from_cpu_data_master >> 2) :
    (shifted_address_to_pipeline_bridge_before_tristate_bridge_s1_from_cpu_instruction_master >> 2);

  assign shifted_address_to_pipeline_bridge_before_tristate_bridge_s1_from_cpu_instruction_master = cpu_instruction_master_address_to_slave;
  //slaveid pipeline_bridge_before_tristate_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_nativeaddress = (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1)? (cpu_data_master_address_to_slave >> 2) :
    (cpu_instruction_master_address_to_slave >> 2);

  //d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer <= 1;
      else 
        d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer <= pipeline_bridge_before_tristate_bridge_s1_end_xfer;
    end


  //pipeline_bridge_before_tristate_bridge_s1_waits_for_read in a cycle, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_waits_for_read = pipeline_bridge_before_tristate_bridge_s1_in_a_read_cycle & pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa;

  //pipeline_bridge_before_tristate_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_in_a_read_cycle = (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1 & cpu_data_master_read) | (cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1 & cpu_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pipeline_bridge_before_tristate_bridge_s1_in_a_read_cycle;

  //pipeline_bridge_before_tristate_bridge_s1_waits_for_write in a cycle, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_waits_for_write = pipeline_bridge_before_tristate_bridge_s1_in_a_write_cycle & pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa;

  //pipeline_bridge_before_tristate_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_s1_in_a_write_cycle = cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pipeline_bridge_before_tristate_bridge_s1_in_a_write_cycle;

  assign wait_for_pipeline_bridge_before_tristate_bridge_s1_counter = 0;
  //pipeline_bridge_before_tristate_bridge_s1_byteenable byte enable port mux, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_byteenable = (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_burstcount = 1;

  //pipeline_bridge_before_tristate_bridge/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_arbiterlock = (cpu_data_master_arbiterlock)? cpu_data_master_arbiterlock :
    cpu_instruction_master_arbiterlock;

  //pipeline_bridge_before_tristate_bridge/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_arbiterlock2 = (cpu_data_master_arbiterlock2)? cpu_data_master_arbiterlock2 :
    cpu_instruction_master_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_s1_debugaccess = (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pipeline_bridge_before_tristate_bridge/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1 + cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_saved_grant_pipeline_bridge_before_tristate_bridge_s1 + cpu_instruction_master_saved_grant_pipeline_bridge_before_tristate_bridge_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_before_tristate_bridge_m1_arbitrator (
                                                              // inputs:
                                                               clk,
                                                               d1_flash_tristate_bridge_avalon_slave_end_xfer,
                                                               ext_flash_s1_wait_counter_eq_0,
                                                               incoming_flash_tristate_bridge_data,
                                                               incoming_flash_tristate_bridge_data_with_Xs_converted_to_0,
                                                               max2_s1_wait_counter_eq_0,
                                                               pipeline_bridge_before_tristate_bridge_m1_address,
                                                               pipeline_bridge_before_tristate_bridge_m1_burstcount,
                                                               pipeline_bridge_before_tristate_bridge_m1_byteenable,
                                                               pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1,
                                                               pipeline_bridge_before_tristate_bridge_m1_chipselect,
                                                               pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1,
                                                               pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1,
                                                               pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1,
                                                               pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1,
                                                               pipeline_bridge_before_tristate_bridge_m1_read,
                                                               pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1,
                                                               pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1,
                                                               pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1,
                                                               pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1,
                                                               pipeline_bridge_before_tristate_bridge_m1_write,
                                                               pipeline_bridge_before_tristate_bridge_m1_writedata,
                                                               reset_n,

                                                              // outputs:
                                                               pipeline_bridge_before_tristate_bridge_m1_address_to_slave,
                                                               pipeline_bridge_before_tristate_bridge_m1_dbs_address,
                                                               pipeline_bridge_before_tristate_bridge_m1_dbs_write_16,
                                                               pipeline_bridge_before_tristate_bridge_m1_latency_counter,
                                                               pipeline_bridge_before_tristate_bridge_m1_readdata,
                                                               pipeline_bridge_before_tristate_bridge_m1_readdatavalid,
                                                               pipeline_bridge_before_tristate_bridge_m1_waitrequest
                                                            )
;

  output  [ 26: 0] pipeline_bridge_before_tristate_bridge_m1_address_to_slave;
  output  [  1: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_address;
  output  [ 15: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_write_16;
  output  [  1: 0] pipeline_bridge_before_tristate_bridge_m1_latency_counter;
  output  [ 31: 0] pipeline_bridge_before_tristate_bridge_m1_readdata;
  output           pipeline_bridge_before_tristate_bridge_m1_readdatavalid;
  output           pipeline_bridge_before_tristate_bridge_m1_waitrequest;
  input            clk;
  input            d1_flash_tristate_bridge_avalon_slave_end_xfer;
  input            ext_flash_s1_wait_counter_eq_0;
  input   [ 31: 0] incoming_flash_tristate_bridge_data;
  input   [ 15: 0] incoming_flash_tristate_bridge_data_with_Xs_converted_to_0;
  input            max2_s1_wait_counter_eq_0;
  input   [ 26: 0] pipeline_bridge_before_tristate_bridge_m1_address;
  input            pipeline_bridge_before_tristate_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_before_tristate_bridge_m1_byteenable;
  input   [  1: 0] pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1;
  input            pipeline_bridge_before_tristate_bridge_m1_chipselect;
  input            pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1;
  input            pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1;
  input            pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1;
  input            pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1;
  input            pipeline_bridge_before_tristate_bridge_m1_read;
  input            pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1;
  input            pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1;
  input            pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1;
  input            pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1;
  input            pipeline_bridge_before_tristate_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_before_tristate_bridge_m1_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire    [  1: 0] p1_pipeline_bridge_before_tristate_bridge_m1_latency_counter;
  reg     [ 26: 0] pipeline_bridge_before_tristate_bridge_m1_address_last_time;
  wire    [ 26: 0] pipeline_bridge_before_tristate_bridge_m1_address_to_slave;
  reg              pipeline_bridge_before_tristate_bridge_m1_burstcount_last_time;
  reg     [  3: 0] pipeline_bridge_before_tristate_bridge_m1_byteenable_last_time;
  reg              pipeline_bridge_before_tristate_bridge_m1_chipselect_last_time;
  reg     [  1: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_address;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_increment;
  reg     [  1: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_rdv_counter;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_rdv_counter_inc;
  wire    [ 15: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_write_16;
  wire             pipeline_bridge_before_tristate_bridge_m1_is_granted_some_slave;
  reg     [  1: 0] pipeline_bridge_before_tristate_bridge_m1_latency_counter;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_m1_next_dbs_rdv_counter;
  reg              pipeline_bridge_before_tristate_bridge_m1_read_but_no_slave_selected;
  reg              pipeline_bridge_before_tristate_bridge_m1_read_last_time;
  wire    [ 31: 0] pipeline_bridge_before_tristate_bridge_m1_readdata;
  wire             pipeline_bridge_before_tristate_bridge_m1_readdatavalid;
  wire             pipeline_bridge_before_tristate_bridge_m1_run;
  wire             pipeline_bridge_before_tristate_bridge_m1_waitrequest;
  reg              pipeline_bridge_before_tristate_bridge_m1_write_last_time;
  reg     [ 31: 0] pipeline_bridge_before_tristate_bridge_m1_writedata_last_time;
  wire             pre_dbs_count_enable;
  wire             pre_flush_pipeline_bridge_before_tristate_bridge_m1_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1 | ~pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1) & ((pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1 | ((pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect) & !pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1 & pipeline_bridge_before_tristate_bridge_m1_dbs_address[1]) | ~pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1)) & ((~pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1 | ~pipeline_bridge_before_tristate_bridge_m1_chipselect | (1 & ((max2_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer)) & pipeline_bridge_before_tristate_bridge_m1_chipselect))) & ((~pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1 | ~pipeline_bridge_before_tristate_bridge_m1_chipselect | (1 & ((max2_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer)) & pipeline_bridge_before_tristate_bridge_m1_chipselect))) & ((~pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1 | ~(pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect) | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer)) & (pipeline_bridge_before_tristate_bridge_m1_dbs_address[1]) & (pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect)))) & ((~pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1 | ~(pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect) | (1 & ((ext_flash_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer)) & (pipeline_bridge_before_tristate_bridge_m1_dbs_address[1]) & (pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect))));

  //cascaded wait assignment, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_m1_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign pipeline_bridge_before_tristate_bridge_m1_address_to_slave = pipeline_bridge_before_tristate_bridge_m1_address[26 : 0];

  //pipeline_bridge_before_tristate_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_read_but_no_slave_selected <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_read_but_no_slave_selected <= (pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect) & pipeline_bridge_before_tristate_bridge_m1_run & ~pipeline_bridge_before_tristate_bridge_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_m1_is_granted_some_slave = pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1 |
    pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_pipeline_bridge_before_tristate_bridge_m1_readdatavalid = pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1 |
    (pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1 & dbs_rdv_counter_overflow);

  //latent slave read data valid which is not flushed, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_m1_readdatavalid = pipeline_bridge_before_tristate_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_before_tristate_bridge_m1_readdatavalid |
    pipeline_bridge_before_tristate_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_before_tristate_bridge_m1_readdatavalid;

  //pipeline_bridge_before_tristate_bridge/m1 readdata mux, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_m1_readdata = ({32 {~pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1}} | incoming_flash_tristate_bridge_data) &
    ({32 {~pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1}} | {incoming_flash_tristate_bridge_data_with_Xs_converted_to_0[15 : 0],
    dbs_latent_16_reg_segment_0});

  //actual waitrequest port, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_m1_waitrequest = ~pipeline_bridge_before_tristate_bridge_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_latency_counter <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_latency_counter <= p1_pipeline_bridge_before_tristate_bridge_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_pipeline_bridge_before_tristate_bridge_m1_latency_counter = ((pipeline_bridge_before_tristate_bridge_m1_run & (pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect)))? latency_load_value :
    (pipeline_bridge_before_tristate_bridge_m1_latency_counter)? pipeline_bridge_before_tristate_bridge_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({2 {pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1}} & 2) |
    ({2 {pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1}} & 2);

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (((~0) & pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1 & (pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect) & !pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1)) |
    ((pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1 & (pipeline_bridge_before_tristate_bridge_m1_read & pipeline_bridge_before_tristate_bridge_m1_chipselect) & 1 & 1 & ({ext_flash_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer}))) |
    ((pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1 & (pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect) & 1 & 1 & ({ext_flash_s1_wait_counter_eq_0 & ~d1_flash_tristate_bridge_avalon_slave_end_xfer})));

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = incoming_flash_tristate_bridge_data_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((pipeline_bridge_before_tristate_bridge_m1_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //mux write dbs 1, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_m1_dbs_write_16 = (pipeline_bridge_before_tristate_bridge_m1_dbs_address[1])? pipeline_bridge_before_tristate_bridge_m1_writedata[31 : 16] :
    pipeline_bridge_before_tristate_bridge_m1_writedata[15 : 0];

  //dbs count increment, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_m1_dbs_increment = (pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = pipeline_bridge_before_tristate_bridge_m1_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = pipeline_bridge_before_tristate_bridge_m1_dbs_address + pipeline_bridge_before_tristate_bridge_m1_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_dbs_address <= 0;
      else if (dbs_count_enable)
          pipeline_bridge_before_tristate_bridge_m1_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign pipeline_bridge_before_tristate_bridge_m1_next_dbs_rdv_counter = pipeline_bridge_before_tristate_bridge_m1_dbs_rdv_counter + pipeline_bridge_before_tristate_bridge_m1_dbs_rdv_counter_inc;

  //pipeline_bridge_before_tristate_bridge_m1_rdv_inc_mux, which is an e_mux
  assign pipeline_bridge_before_tristate_bridge_m1_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          pipeline_bridge_before_tristate_bridge_m1_dbs_rdv_counter <= pipeline_bridge_before_tristate_bridge_m1_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = pipeline_bridge_before_tristate_bridge_m1_dbs_rdv_counter[1] & ~pipeline_bridge_before_tristate_bridge_m1_next_dbs_rdv_counter[1];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pipeline_bridge_before_tristate_bridge_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_address_last_time <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_address_last_time <= pipeline_bridge_before_tristate_bridge_m1_address;
    end


  //pipeline_bridge_before_tristate_bridge/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= pipeline_bridge_before_tristate_bridge_m1_waitrequest & pipeline_bridge_before_tristate_bridge_m1_chipselect;
    end


  //pipeline_bridge_before_tristate_bridge_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_before_tristate_bridge_m1_address != pipeline_bridge_before_tristate_bridge_m1_address_last_time))
        begin
          $write("%0d ns: pipeline_bridge_before_tristate_bridge_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_before_tristate_bridge_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_chipselect_last_time <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_chipselect_last_time <= pipeline_bridge_before_tristate_bridge_m1_chipselect;
    end


  //pipeline_bridge_before_tristate_bridge_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_before_tristate_bridge_m1_chipselect != pipeline_bridge_before_tristate_bridge_m1_chipselect_last_time))
        begin
          $write("%0d ns: pipeline_bridge_before_tristate_bridge_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_before_tristate_bridge_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_burstcount_last_time <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_burstcount_last_time <= pipeline_bridge_before_tristate_bridge_m1_burstcount;
    end


  //pipeline_bridge_before_tristate_bridge_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_before_tristate_bridge_m1_burstcount != pipeline_bridge_before_tristate_bridge_m1_burstcount_last_time))
        begin
          $write("%0d ns: pipeline_bridge_before_tristate_bridge_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_before_tristate_bridge_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_byteenable_last_time <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_byteenable_last_time <= pipeline_bridge_before_tristate_bridge_m1_byteenable;
    end


  //pipeline_bridge_before_tristate_bridge_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_before_tristate_bridge_m1_byteenable != pipeline_bridge_before_tristate_bridge_m1_byteenable_last_time))
        begin
          $write("%0d ns: pipeline_bridge_before_tristate_bridge_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_before_tristate_bridge_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_read_last_time <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_read_last_time <= pipeline_bridge_before_tristate_bridge_m1_read;
    end


  //pipeline_bridge_before_tristate_bridge_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_before_tristate_bridge_m1_read != pipeline_bridge_before_tristate_bridge_m1_read_last_time))
        begin
          $write("%0d ns: pipeline_bridge_before_tristate_bridge_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_before_tristate_bridge_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_write_last_time <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_write_last_time <= pipeline_bridge_before_tristate_bridge_m1_write;
    end


  //pipeline_bridge_before_tristate_bridge_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_before_tristate_bridge_m1_write != pipeline_bridge_before_tristate_bridge_m1_write_last_time))
        begin
          $write("%0d ns: pipeline_bridge_before_tristate_bridge_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_before_tristate_bridge_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_before_tristate_bridge_m1_writedata_last_time <= 0;
      else 
        pipeline_bridge_before_tristate_bridge_m1_writedata_last_time <= pipeline_bridge_before_tristate_bridge_m1_writedata;
    end


  //pipeline_bridge_before_tristate_bridge_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_before_tristate_bridge_m1_writedata != pipeline_bridge_before_tristate_bridge_m1_writedata_last_time) & (pipeline_bridge_before_tristate_bridge_m1_write & pipeline_bridge_before_tristate_bridge_m1_chipselect))
        begin
          $write("%0d ns: pipeline_bridge_before_tristate_bridge_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_before_tristate_bridge_bridge_arbitrator 
;



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pll_s1_arbitrator (
                           // inputs:
                            clk,
                            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave,
                            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_nativeaddress,
                            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read,
                            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write,
                            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata,
                            pll_s1_readdata,
                            pll_s1_resetrequest,
                            reset_n,

                           // outputs:
                            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1,
                            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1,
                            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_data_valid_pll_s1,
                            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1,
                            d1_pll_s1_end_xfer,
                            pll_s1_address,
                            pll_s1_chipselect,
                            pll_s1_read,
                            pll_s1_readdata_from_sa,
                            pll_s1_reset_n,
                            pll_s1_resetrequest_from_sa,
                            pll_s1_write,
                            pll_s1_writedata
                         )
;

  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_data_valid_pll_s1;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1;
  output           d1_pll_s1_end_xfer;
  output  [  2: 0] pll_s1_address;
  output           pll_s1_chipselect;
  output           pll_s1_read;
  output  [ 15: 0] pll_s1_readdata_from_sa;
  output           pll_s1_reset_n;
  output           pll_s1_resetrequest_from_sa;
  output           pll_s1_write;
  output  [ 15: 0] pll_s1_writedata;
  input            clk;
  input   [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave;
  input   [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_nativeaddress;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata;
  input   [ 15: 0] pll_s1_readdata;
  input            pll_s1_resetrequest;
  input            reset_n;

  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_arbiterlock;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_arbiterlock2;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_continuerequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_data_valid_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_saved_grant_pll_s1;
  reg              d1_pll_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pll_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  2: 0] pll_s1_address;
  wire             pll_s1_allgrants;
  wire             pll_s1_allow_new_arb_cycle;
  wire             pll_s1_any_bursting_master_saved_grant;
  wire             pll_s1_any_continuerequest;
  wire             pll_s1_arb_counter_enable;
  reg              pll_s1_arb_share_counter;
  wire             pll_s1_arb_share_counter_next_value;
  wire             pll_s1_arb_share_set_values;
  wire             pll_s1_beginbursttransfer_internal;
  wire             pll_s1_begins_xfer;
  wire             pll_s1_chipselect;
  wire             pll_s1_end_xfer;
  wire             pll_s1_firsttransfer;
  wire             pll_s1_grant_vector;
  wire             pll_s1_in_a_read_cycle;
  wire             pll_s1_in_a_write_cycle;
  wire             pll_s1_master_qreq_vector;
  wire             pll_s1_non_bursting_master_requests;
  wire             pll_s1_read;
  wire    [ 15: 0] pll_s1_readdata_from_sa;
  reg              pll_s1_reg_firsttransfer;
  wire             pll_s1_reset_n;
  wire             pll_s1_resetrequest_from_sa;
  reg              pll_s1_slavearbiterlockenable;
  wire             pll_s1_slavearbiterlockenable2;
  wire             pll_s1_unreg_firsttransfer;
  wire             pll_s1_waits_for_read;
  wire             pll_s1_waits_for_write;
  wire             pll_s1_write;
  wire    [ 15: 0] pll_s1_writedata;
  wire             wait_for_pll_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pll_s1_end_xfer;
    end


  assign pll_s1_begins_xfer = ~d1_reasons_to_wait & ((cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1));
  //assign pll_s1_readdata_from_sa = pll_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pll_s1_readdata_from_sa = pll_s1_readdata;

  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1 = (1) & (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read | cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write);
  //pll_s1_arb_share_counter set values, which is an e_mux
  assign pll_s1_arb_share_set_values = 1;

  //pll_s1_non_bursting_master_requests mux, which is an e_mux
  assign pll_s1_non_bursting_master_requests = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1;

  //pll_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pll_s1_any_bursting_master_saved_grant = 0;

  //pll_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pll_s1_arb_share_counter_next_value = pll_s1_firsttransfer ? (pll_s1_arb_share_set_values - 1) : |pll_s1_arb_share_counter ? (pll_s1_arb_share_counter - 1) : 0;

  //pll_s1_allgrants all slave grants, which is an e_mux
  assign pll_s1_allgrants = |pll_s1_grant_vector;

  //pll_s1_end_xfer assignment, which is an e_assign
  assign pll_s1_end_xfer = ~(pll_s1_waits_for_read | pll_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pll_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pll_s1 = pll_s1_end_xfer & (~pll_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pll_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pll_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pll_s1 & pll_s1_allgrants) | (end_xfer_arb_share_counter_term_pll_s1 & ~pll_s1_non_bursting_master_requests);

  //pll_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pll_s1_arb_share_counter <= 0;
      else if (pll_s1_arb_counter_enable)
          pll_s1_arb_share_counter <= pll_s1_arb_share_counter_next_value;
    end


  //pll_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pll_s1_slavearbiterlockenable <= 0;
      else if ((|pll_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pll_s1) | (end_xfer_arb_share_counter_term_pll_s1 & ~pll_s1_non_bursting_master_requests))
          pll_s1_slavearbiterlockenable <= |pll_s1_arb_share_counter_next_value;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_0/out pll/s1 arbiterlock, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_arbiterlock = pll_s1_slavearbiterlockenable & cycloneIII_3c120_niosII_standard_sopc_clock_0_out_continuerequest;

  //pll_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pll_s1_slavearbiterlockenable2 = |pll_s1_arb_share_counter_next_value;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0/out pll/s1 arbiterlock2, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_arbiterlock2 = pll_s1_slavearbiterlockenable2 & cycloneIII_3c120_niosII_standard_sopc_clock_0_out_continuerequest;

  //pll_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign pll_s1_any_continuerequest = 1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_continuerequest continued request, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_continuerequest = 1;

  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1 = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1;
  //pll_s1_writedata mux, which is an e_mux
  assign pll_s1_writedata = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata;

  //master is always granted when requested
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1 = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0/out saved-grant pll/s1, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_saved_grant_pll_s1 = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1;

  //allow new arb cycle for pll/s1, which is an e_assign
  assign pll_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign pll_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign pll_s1_master_qreq_vector = 1;

  //pll_s1_reset_n assignment, which is an e_assign
  assign pll_s1_reset_n = reset_n;

  //assign pll_s1_resetrequest_from_sa = pll_s1_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pll_s1_resetrequest_from_sa = pll_s1_resetrequest;

  assign pll_s1_chipselect = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1;
  //pll_s1_firsttransfer first transaction, which is an e_assign
  assign pll_s1_firsttransfer = pll_s1_begins_xfer ? pll_s1_unreg_firsttransfer : pll_s1_reg_firsttransfer;

  //pll_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pll_s1_unreg_firsttransfer = ~(pll_s1_slavearbiterlockenable & pll_s1_any_continuerequest);

  //pll_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pll_s1_reg_firsttransfer <= 1'b1;
      else if (pll_s1_begins_xfer)
          pll_s1_reg_firsttransfer <= pll_s1_unreg_firsttransfer;
    end


  //pll_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pll_s1_beginbursttransfer_internal = pll_s1_begins_xfer;

  //pll_s1_read assignment, which is an e_mux
  assign pll_s1_read = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read;

  //pll_s1_write assignment, which is an e_mux
  assign pll_s1_write = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write;

  //pll_s1_address mux, which is an e_mux
  assign pll_s1_address = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_nativeaddress;

  //d1_pll_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pll_s1_end_xfer <= 1;
      else 
        d1_pll_s1_end_xfer <= pll_s1_end_xfer;
    end


  //pll_s1_waits_for_read in a cycle, which is an e_mux
  assign pll_s1_waits_for_read = pll_s1_in_a_read_cycle & pll_s1_begins_xfer;

  //pll_s1_in_a_read_cycle assignment, which is an e_assign
  assign pll_s1_in_a_read_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pll_s1_in_a_read_cycle;

  //pll_s1_waits_for_write in a cycle, which is an e_mux
  assign pll_s1_waits_for_write = pll_s1_in_a_write_cycle & 0;

  //pll_s1_in_a_write_cycle assignment, which is an e_assign
  assign pll_s1_in_a_write_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pll_s1_in_a_write_cycle;

  assign wait_for_pll_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pll/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_csr_arbitrator (
                                 // inputs:
                                  clk,
                                  cpu_data_master_address_to_slave,
                                  cpu_data_master_latency_counter,
                                  cpu_data_master_read,
                                  cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                  cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                  cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register,
                                  cpu_data_master_write,
                                  cpu_data_master_writedata,
                                  reset_n,
                                  sgdma_rx_csr_irq,
                                  sgdma_rx_csr_readdata,

                                 // outputs:
                                  cpu_data_master_granted_sgdma_rx_csr,
                                  cpu_data_master_qualified_request_sgdma_rx_csr,
                                  cpu_data_master_read_data_valid_sgdma_rx_csr,
                                  cpu_data_master_requests_sgdma_rx_csr,
                                  d1_sgdma_rx_csr_end_xfer,
                                  sgdma_rx_csr_address,
                                  sgdma_rx_csr_chipselect,
                                  sgdma_rx_csr_irq_from_sa,
                                  sgdma_rx_csr_read,
                                  sgdma_rx_csr_readdata_from_sa,
                                  sgdma_rx_csr_reset_n,
                                  sgdma_rx_csr_write,
                                  sgdma_rx_csr_writedata
                               )
;

  output           cpu_data_master_granted_sgdma_rx_csr;
  output           cpu_data_master_qualified_request_sgdma_rx_csr;
  output           cpu_data_master_read_data_valid_sgdma_rx_csr;
  output           cpu_data_master_requests_sgdma_rx_csr;
  output           d1_sgdma_rx_csr_end_xfer;
  output  [  3: 0] sgdma_rx_csr_address;
  output           sgdma_rx_csr_chipselect;
  output           sgdma_rx_csr_irq_from_sa;
  output           sgdma_rx_csr_read;
  output  [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  output           sgdma_rx_csr_reset_n;
  output           sgdma_rx_csr_write;
  output  [ 31: 0] sgdma_rx_csr_writedata;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input            sgdma_rx_csr_irq;
  input   [ 31: 0] sgdma_rx_csr_readdata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_sgdma_rx_csr;
  wire             cpu_data_master_qualified_request_sgdma_rx_csr;
  wire             cpu_data_master_read_data_valid_sgdma_rx_csr;
  wire             cpu_data_master_requests_sgdma_rx_csr;
  wire             cpu_data_master_saved_grant_sgdma_rx_csr;
  reg              d1_reasons_to_wait;
  reg              d1_sgdma_rx_csr_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sgdma_rx_csr;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  3: 0] sgdma_rx_csr_address;
  wire             sgdma_rx_csr_allgrants;
  wire             sgdma_rx_csr_allow_new_arb_cycle;
  wire             sgdma_rx_csr_any_bursting_master_saved_grant;
  wire             sgdma_rx_csr_any_continuerequest;
  wire             sgdma_rx_csr_arb_counter_enable;
  reg              sgdma_rx_csr_arb_share_counter;
  wire             sgdma_rx_csr_arb_share_counter_next_value;
  wire             sgdma_rx_csr_arb_share_set_values;
  wire             sgdma_rx_csr_beginbursttransfer_internal;
  wire             sgdma_rx_csr_begins_xfer;
  wire             sgdma_rx_csr_chipselect;
  wire             sgdma_rx_csr_end_xfer;
  wire             sgdma_rx_csr_firsttransfer;
  wire             sgdma_rx_csr_grant_vector;
  wire             sgdma_rx_csr_in_a_read_cycle;
  wire             sgdma_rx_csr_in_a_write_cycle;
  wire             sgdma_rx_csr_irq_from_sa;
  wire             sgdma_rx_csr_master_qreq_vector;
  wire             sgdma_rx_csr_non_bursting_master_requests;
  wire             sgdma_rx_csr_read;
  wire    [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  reg              sgdma_rx_csr_reg_firsttransfer;
  wire             sgdma_rx_csr_reset_n;
  reg              sgdma_rx_csr_slavearbiterlockenable;
  wire             sgdma_rx_csr_slavearbiterlockenable2;
  wire             sgdma_rx_csr_unreg_firsttransfer;
  wire             sgdma_rx_csr_waits_for_read;
  wire             sgdma_rx_csr_waits_for_write;
  wire             sgdma_rx_csr_write;
  wire    [ 31: 0] sgdma_rx_csr_writedata;
  wire    [ 28: 0] shifted_address_to_sgdma_rx_csr_from_cpu_data_master;
  wire             wait_for_sgdma_rx_csr_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sgdma_rx_csr_end_xfer;
    end


  assign sgdma_rx_csr_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_sgdma_rx_csr));
  //assign sgdma_rx_csr_readdata_from_sa = sgdma_rx_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_rx_csr_readdata_from_sa = sgdma_rx_csr_readdata;

  assign cpu_data_master_requests_sgdma_rx_csr = ({cpu_data_master_address_to_slave[28 : 6] , 6'b0} == 29'h1002000) & (cpu_data_master_read | cpu_data_master_write);
  //sgdma_rx_csr_arb_share_counter set values, which is an e_mux
  assign sgdma_rx_csr_arb_share_set_values = 1;

  //sgdma_rx_csr_non_bursting_master_requests mux, which is an e_mux
  assign sgdma_rx_csr_non_bursting_master_requests = cpu_data_master_requests_sgdma_rx_csr;

  //sgdma_rx_csr_any_bursting_master_saved_grant mux, which is an e_mux
  assign sgdma_rx_csr_any_bursting_master_saved_grant = 0;

  //sgdma_rx_csr_arb_share_counter_next_value assignment, which is an e_assign
  assign sgdma_rx_csr_arb_share_counter_next_value = sgdma_rx_csr_firsttransfer ? (sgdma_rx_csr_arb_share_set_values - 1) : |sgdma_rx_csr_arb_share_counter ? (sgdma_rx_csr_arb_share_counter - 1) : 0;

  //sgdma_rx_csr_allgrants all slave grants, which is an e_mux
  assign sgdma_rx_csr_allgrants = |sgdma_rx_csr_grant_vector;

  //sgdma_rx_csr_end_xfer assignment, which is an e_assign
  assign sgdma_rx_csr_end_xfer = ~(sgdma_rx_csr_waits_for_read | sgdma_rx_csr_waits_for_write);

  //end_xfer_arb_share_counter_term_sgdma_rx_csr arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sgdma_rx_csr = sgdma_rx_csr_end_xfer & (~sgdma_rx_csr_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sgdma_rx_csr_arb_share_counter arbitration counter enable, which is an e_assign
  assign sgdma_rx_csr_arb_counter_enable = (end_xfer_arb_share_counter_term_sgdma_rx_csr & sgdma_rx_csr_allgrants) | (end_xfer_arb_share_counter_term_sgdma_rx_csr & ~sgdma_rx_csr_non_bursting_master_requests);

  //sgdma_rx_csr_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_csr_arb_share_counter <= 0;
      else if (sgdma_rx_csr_arb_counter_enable)
          sgdma_rx_csr_arb_share_counter <= sgdma_rx_csr_arb_share_counter_next_value;
    end


  //sgdma_rx_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_csr_slavearbiterlockenable <= 0;
      else if ((|sgdma_rx_csr_master_qreq_vector & end_xfer_arb_share_counter_term_sgdma_rx_csr) | (end_xfer_arb_share_counter_term_sgdma_rx_csr & ~sgdma_rx_csr_non_bursting_master_requests))
          sgdma_rx_csr_slavearbiterlockenable <= |sgdma_rx_csr_arb_share_counter_next_value;
    end


  //cpu/data_master sgdma_rx/csr arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = sgdma_rx_csr_slavearbiterlockenable & cpu_data_master_continuerequest;

  //sgdma_rx_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sgdma_rx_csr_slavearbiterlockenable2 = |sgdma_rx_csr_arb_share_counter_next_value;

  //cpu/data_master sgdma_rx/csr arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = sgdma_rx_csr_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //sgdma_rx_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sgdma_rx_csr_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_sgdma_rx_csr = cpu_data_master_requests_sgdma_rx_csr & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_sgdma_rx_csr, which is an e_mux
  assign cpu_data_master_read_data_valid_sgdma_rx_csr = cpu_data_master_granted_sgdma_rx_csr & cpu_data_master_read & ~sgdma_rx_csr_waits_for_read;

  //sgdma_rx_csr_writedata mux, which is an e_mux
  assign sgdma_rx_csr_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_sgdma_rx_csr = cpu_data_master_qualified_request_sgdma_rx_csr;

  //cpu/data_master saved-grant sgdma_rx/csr, which is an e_assign
  assign cpu_data_master_saved_grant_sgdma_rx_csr = cpu_data_master_requests_sgdma_rx_csr;

  //allow new arb cycle for sgdma_rx/csr, which is an e_assign
  assign sgdma_rx_csr_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sgdma_rx_csr_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sgdma_rx_csr_master_qreq_vector = 1;

  //sgdma_rx_csr_reset_n assignment, which is an e_assign
  assign sgdma_rx_csr_reset_n = reset_n;

  assign sgdma_rx_csr_chipselect = cpu_data_master_granted_sgdma_rx_csr;
  //sgdma_rx_csr_firsttransfer first transaction, which is an e_assign
  assign sgdma_rx_csr_firsttransfer = sgdma_rx_csr_begins_xfer ? sgdma_rx_csr_unreg_firsttransfer : sgdma_rx_csr_reg_firsttransfer;

  //sgdma_rx_csr_unreg_firsttransfer first transaction, which is an e_assign
  assign sgdma_rx_csr_unreg_firsttransfer = ~(sgdma_rx_csr_slavearbiterlockenable & sgdma_rx_csr_any_continuerequest);

  //sgdma_rx_csr_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_csr_reg_firsttransfer <= 1'b1;
      else if (sgdma_rx_csr_begins_xfer)
          sgdma_rx_csr_reg_firsttransfer <= sgdma_rx_csr_unreg_firsttransfer;
    end


  //sgdma_rx_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sgdma_rx_csr_beginbursttransfer_internal = sgdma_rx_csr_begins_xfer;

  //sgdma_rx_csr_read assignment, which is an e_mux
  assign sgdma_rx_csr_read = cpu_data_master_granted_sgdma_rx_csr & cpu_data_master_read;

  //sgdma_rx_csr_write assignment, which is an e_mux
  assign sgdma_rx_csr_write = cpu_data_master_granted_sgdma_rx_csr & cpu_data_master_write;

  assign shifted_address_to_sgdma_rx_csr_from_cpu_data_master = cpu_data_master_address_to_slave;
  //sgdma_rx_csr_address mux, which is an e_mux
  assign sgdma_rx_csr_address = shifted_address_to_sgdma_rx_csr_from_cpu_data_master >> 2;

  //d1_sgdma_rx_csr_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sgdma_rx_csr_end_xfer <= 1;
      else 
        d1_sgdma_rx_csr_end_xfer <= sgdma_rx_csr_end_xfer;
    end


  //sgdma_rx_csr_waits_for_read in a cycle, which is an e_mux
  assign sgdma_rx_csr_waits_for_read = sgdma_rx_csr_in_a_read_cycle & sgdma_rx_csr_begins_xfer;

  //sgdma_rx_csr_in_a_read_cycle assignment, which is an e_assign
  assign sgdma_rx_csr_in_a_read_cycle = cpu_data_master_granted_sgdma_rx_csr & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sgdma_rx_csr_in_a_read_cycle;

  //sgdma_rx_csr_waits_for_write in a cycle, which is an e_mux
  assign sgdma_rx_csr_waits_for_write = sgdma_rx_csr_in_a_write_cycle & 0;

  //sgdma_rx_csr_in_a_write_cycle assignment, which is an e_assign
  assign sgdma_rx_csr_in_a_write_cycle = cpu_data_master_granted_sgdma_rx_csr & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sgdma_rx_csr_in_a_write_cycle;

  assign wait_for_sgdma_rx_csr_counter = 0;
  //assign sgdma_rx_csr_irq_from_sa = sgdma_rx_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_rx_csr_irq_from_sa = sgdma_rx_csr_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx/csr enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_in_arbitrator (
                                // inputs:
                                 clk,
                                 reset_n,
                                 sgdma_rx_in_ready,
                                 tse_mac_receive_data,
                                 tse_mac_receive_empty,
                                 tse_mac_receive_endofpacket,
                                 tse_mac_receive_error,
                                 tse_mac_receive_startofpacket,
                                 tse_mac_receive_valid,

                                // outputs:
                                 sgdma_rx_in_data,
                                 sgdma_rx_in_empty,
                                 sgdma_rx_in_endofpacket,
                                 sgdma_rx_in_error,
                                 sgdma_rx_in_ready_from_sa,
                                 sgdma_rx_in_startofpacket,
                                 sgdma_rx_in_valid
                              )
;

  output  [ 31: 0] sgdma_rx_in_data;
  output  [  1: 0] sgdma_rx_in_empty;
  output           sgdma_rx_in_endofpacket;
  output  [  5: 0] sgdma_rx_in_error;
  output           sgdma_rx_in_ready_from_sa;
  output           sgdma_rx_in_startofpacket;
  output           sgdma_rx_in_valid;
  input            clk;
  input            reset_n;
  input            sgdma_rx_in_ready;
  input   [ 31: 0] tse_mac_receive_data;
  input   [  1: 0] tse_mac_receive_empty;
  input            tse_mac_receive_endofpacket;
  input   [  5: 0] tse_mac_receive_error;
  input            tse_mac_receive_startofpacket;
  input            tse_mac_receive_valid;

  wire    [ 31: 0] sgdma_rx_in_data;
  wire    [  1: 0] sgdma_rx_in_empty;
  wire             sgdma_rx_in_endofpacket;
  wire    [  5: 0] sgdma_rx_in_error;
  wire             sgdma_rx_in_ready_from_sa;
  wire             sgdma_rx_in_startofpacket;
  wire             sgdma_rx_in_valid;
  //mux sgdma_rx_in_data, which is an e_mux
  assign sgdma_rx_in_data = tse_mac_receive_data;

  //mux sgdma_rx_in_empty, which is an e_mux
  assign sgdma_rx_in_empty = tse_mac_receive_empty;

  //mux sgdma_rx_in_endofpacket, which is an e_mux
  assign sgdma_rx_in_endofpacket = tse_mac_receive_endofpacket;

  //mux sgdma_rx_in_error, which is an e_mux
  assign sgdma_rx_in_error = tse_mac_receive_error;

  //assign sgdma_rx_in_ready_from_sa = sgdma_rx_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_rx_in_ready_from_sa = sgdma_rx_in_ready;

  //mux sgdma_rx_in_startofpacket, which is an e_mux
  assign sgdma_rx_in_startofpacket = tse_mac_receive_startofpacket;

  //mux sgdma_rx_in_valid, which is an e_mux
  assign sgdma_rx_in_valid = tse_mac_receive_valid;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_descriptor_read_arbitrator (
                                             // inputs:
                                              clk,
                                              d1_descriptor_memory_s1_end_xfer,
                                              descriptor_memory_s1_readdata_from_sa,
                                              reset_n,
                                              sgdma_rx_descriptor_read_address,
                                              sgdma_rx_descriptor_read_granted_descriptor_memory_s1,
                                              sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1,
                                              sgdma_rx_descriptor_read_read,
                                              sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1,
                                              sgdma_rx_descriptor_read_requests_descriptor_memory_s1,

                                             // outputs:
                                              sgdma_rx_descriptor_read_address_to_slave,
                                              sgdma_rx_descriptor_read_latency_counter,
                                              sgdma_rx_descriptor_read_readdata,
                                              sgdma_rx_descriptor_read_readdatavalid,
                                              sgdma_rx_descriptor_read_waitrequest
                                           )
;

  output  [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  output           sgdma_rx_descriptor_read_latency_counter;
  output  [ 31: 0] sgdma_rx_descriptor_read_readdata;
  output           sgdma_rx_descriptor_read_readdatavalid;
  output           sgdma_rx_descriptor_read_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s1_end_xfer;
  input   [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_descriptor_read_address;
  input            sgdma_rx_descriptor_read_granted_descriptor_memory_s1;
  input            sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;
  input            sgdma_rx_descriptor_read_read;
  input            sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;
  input            sgdma_rx_descriptor_read_requests_descriptor_memory_s1;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_sgdma_rx_descriptor_read_latency_counter;
  wire             pre_flush_sgdma_rx_descriptor_read_readdatavalid;
  wire             r_0;
  reg     [ 31: 0] sgdma_rx_descriptor_read_address_last_time;
  wire    [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  wire             sgdma_rx_descriptor_read_is_granted_some_slave;
  reg              sgdma_rx_descriptor_read_latency_counter;
  reg              sgdma_rx_descriptor_read_read_but_no_slave_selected;
  reg              sgdma_rx_descriptor_read_read_last_time;
  wire    [ 31: 0] sgdma_rx_descriptor_read_readdata;
  wire             sgdma_rx_descriptor_read_readdatavalid;
  wire             sgdma_rx_descriptor_read_run;
  wire             sgdma_rx_descriptor_read_waitrequest;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 | ~sgdma_rx_descriptor_read_requests_descriptor_memory_s1) & (sgdma_rx_descriptor_read_granted_descriptor_memory_s1 | ~sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1) & ((~sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 | ~(sgdma_rx_descriptor_read_read) | (1 & (sgdma_rx_descriptor_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_rx_descriptor_read_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_rx_descriptor_read_address_to_slave = {20'b1000000000000,
    sgdma_rx_descriptor_read_address[11 : 0]};

  //sgdma_rx_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_read_but_no_slave_selected <= 0;
      else 
        sgdma_rx_descriptor_read_read_but_no_slave_selected <= sgdma_rx_descriptor_read_read & sgdma_rx_descriptor_read_run & ~sgdma_rx_descriptor_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign sgdma_rx_descriptor_read_is_granted_some_slave = sgdma_rx_descriptor_read_granted_descriptor_memory_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_sgdma_rx_descriptor_read_readdatavalid = sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign sgdma_rx_descriptor_read_readdatavalid = sgdma_rx_descriptor_read_read_but_no_slave_selected |
    pre_flush_sgdma_rx_descriptor_read_readdatavalid;

  //sgdma_rx/descriptor_read readdata mux, which is an e_mux
  assign sgdma_rx_descriptor_read_readdata = descriptor_memory_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign sgdma_rx_descriptor_read_waitrequest = ~sgdma_rx_descriptor_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_latency_counter <= 0;
      else 
        sgdma_rx_descriptor_read_latency_counter <= p1_sgdma_rx_descriptor_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_sgdma_rx_descriptor_read_latency_counter = ((sgdma_rx_descriptor_read_run & sgdma_rx_descriptor_read_read))? latency_load_value :
    (sgdma_rx_descriptor_read_latency_counter)? sgdma_rx_descriptor_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {sgdma_rx_descriptor_read_requests_descriptor_memory_s1}} & 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx_descriptor_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_address_last_time <= 0;
      else 
        sgdma_rx_descriptor_read_address_last_time <= sgdma_rx_descriptor_read_address;
    end


  //sgdma_rx/descriptor_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_rx_descriptor_read_waitrequest & (sgdma_rx_descriptor_read_read);
    end


  //sgdma_rx_descriptor_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_read_address != sgdma_rx_descriptor_read_address_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_descriptor_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_read_read_last_time <= 0;
      else 
        sgdma_rx_descriptor_read_read_last_time <= sgdma_rx_descriptor_read_read;
    end


  //sgdma_rx_descriptor_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_read_read != sgdma_rx_descriptor_read_read_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_descriptor_write_arbitrator (
                                              // inputs:
                                               clk,
                                               d1_descriptor_memory_s1_end_xfer,
                                               reset_n,
                                               sgdma_rx_descriptor_write_address,
                                               sgdma_rx_descriptor_write_granted_descriptor_memory_s1,
                                               sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1,
                                               sgdma_rx_descriptor_write_requests_descriptor_memory_s1,
                                               sgdma_rx_descriptor_write_write,
                                               sgdma_rx_descriptor_write_writedata,

                                              // outputs:
                                               sgdma_rx_descriptor_write_address_to_slave,
                                               sgdma_rx_descriptor_write_waitrequest
                                            )
;

  output  [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  output           sgdma_rx_descriptor_write_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s1_end_xfer;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_descriptor_write_address;
  input            sgdma_rx_descriptor_write_granted_descriptor_memory_s1;
  input            sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;
  input            sgdma_rx_descriptor_write_requests_descriptor_memory_s1;
  input            sgdma_rx_descriptor_write_write;
  input   [ 31: 0] sgdma_rx_descriptor_write_writedata;

  reg              active_and_waiting_last_time;
  wire             r_0;
  reg     [ 31: 0] sgdma_rx_descriptor_write_address_last_time;
  wire    [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  wire             sgdma_rx_descriptor_write_run;
  wire             sgdma_rx_descriptor_write_waitrequest;
  reg              sgdma_rx_descriptor_write_write_last_time;
  reg     [ 31: 0] sgdma_rx_descriptor_write_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 | ~sgdma_rx_descriptor_write_requests_descriptor_memory_s1) & (sgdma_rx_descriptor_write_granted_descriptor_memory_s1 | ~sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1) & ((~sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 | ~(sgdma_rx_descriptor_write_write) | (1 & (sgdma_rx_descriptor_write_write))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_rx_descriptor_write_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_rx_descriptor_write_address_to_slave = {20'b1000000000000,
    sgdma_rx_descriptor_write_address[11 : 0]};

  //actual waitrequest port, which is an e_assign
  assign sgdma_rx_descriptor_write_waitrequest = ~sgdma_rx_descriptor_write_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx_descriptor_write_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_write_address_last_time <= 0;
      else 
        sgdma_rx_descriptor_write_address_last_time <= sgdma_rx_descriptor_write_address;
    end


  //sgdma_rx/descriptor_write waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_rx_descriptor_write_waitrequest & (sgdma_rx_descriptor_write_write);
    end


  //sgdma_rx_descriptor_write_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_write_address != sgdma_rx_descriptor_write_address_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_write_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_descriptor_write_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_write_write_last_time <= 0;
      else 
        sgdma_rx_descriptor_write_write_last_time <= sgdma_rx_descriptor_write_write;
    end


  //sgdma_rx_descriptor_write_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_write_write != sgdma_rx_descriptor_write_write_last_time))
        begin
          $write("%0d ns: sgdma_rx_descriptor_write_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_descriptor_write_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_descriptor_write_writedata_last_time <= 0;
      else 
        sgdma_rx_descriptor_write_writedata_last_time <= sgdma_rx_descriptor_write_writedata;
    end


  //sgdma_rx_descriptor_write_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_descriptor_write_writedata != sgdma_rx_descriptor_write_writedata_last_time) & sgdma_rx_descriptor_write_write)
        begin
          $write("%0d ns: sgdma_rx_descriptor_write_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_rx_m_write_arbitrator (
                                     // inputs:
                                      clk,
                                      cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
                                      d1_cpu_ddr_clock_bridge_s1_end_xfer,
                                      reset_n,
                                      sgdma_rx_m_write_address,
                                      sgdma_rx_m_write_byteenable,
                                      sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1,
                                      sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1,
                                      sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1,
                                      sgdma_rx_m_write_write,
                                      sgdma_rx_m_write_writedata,

                                     // outputs:
                                      sgdma_rx_m_write_address_to_slave,
                                      sgdma_rx_m_write_waitrequest
                                   )
;

  output  [ 31: 0] sgdma_rx_m_write_address_to_slave;
  output           sgdma_rx_m_write_waitrequest;
  input            clk;
  input            cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  input            d1_cpu_ddr_clock_bridge_s1_end_xfer;
  input            reset_n;
  input   [ 31: 0] sgdma_rx_m_write_address;
  input   [  3: 0] sgdma_rx_m_write_byteenable;
  input            sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1;
  input            sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1;
  input            sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1;
  input            sgdma_rx_m_write_write;
  input   [ 31: 0] sgdma_rx_m_write_writedata;

  reg              active_and_waiting_last_time;
  wire             r_0;
  reg     [ 31: 0] sgdma_rx_m_write_address_last_time;
  wire    [ 31: 0] sgdma_rx_m_write_address_to_slave;
  reg     [  3: 0] sgdma_rx_m_write_byteenable_last_time;
  wire             sgdma_rx_m_write_run;
  wire             sgdma_rx_m_write_waitrequest;
  reg              sgdma_rx_m_write_write_last_time;
  reg     [ 31: 0] sgdma_rx_m_write_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1 | ~sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1) & (sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1 | ~sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1) & ((~sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1 | ~(sgdma_rx_m_write_write) | (1 & ~cpu_ddr_clock_bridge_s1_waitrequest_from_sa & (sgdma_rx_m_write_write))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_rx_m_write_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_rx_m_write_address_to_slave = {6'b111,
    sgdma_rx_m_write_address[25 : 0]};

  //actual waitrequest port, which is an e_assign
  assign sgdma_rx_m_write_waitrequest = ~sgdma_rx_m_write_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_rx_m_write_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_address_last_time <= 0;
      else 
        sgdma_rx_m_write_address_last_time <= sgdma_rx_m_write_address;
    end


  //sgdma_rx/m_write waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_rx_m_write_waitrequest & (sgdma_rx_m_write_write);
    end


  //sgdma_rx_m_write_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_address != sgdma_rx_m_write_address_last_time))
        begin
          $write("%0d ns: sgdma_rx_m_write_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_m_write_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_byteenable_last_time <= 0;
      else 
        sgdma_rx_m_write_byteenable_last_time <= sgdma_rx_m_write_byteenable;
    end


  //sgdma_rx_m_write_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_byteenable != sgdma_rx_m_write_byteenable_last_time))
        begin
          $write("%0d ns: sgdma_rx_m_write_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_m_write_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_write_last_time <= 0;
      else 
        sgdma_rx_m_write_write_last_time <= sgdma_rx_m_write_write;
    end


  //sgdma_rx_m_write_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_write != sgdma_rx_m_write_write_last_time))
        begin
          $write("%0d ns: sgdma_rx_m_write_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_rx_m_write_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_rx_m_write_writedata_last_time <= 0;
      else 
        sgdma_rx_m_write_writedata_last_time <= sgdma_rx_m_write_writedata;
    end


  //sgdma_rx_m_write_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_rx_m_write_writedata != sgdma_rx_m_write_writedata_last_time) & sgdma_rx_m_write_write)
        begin
          $write("%0d ns: sgdma_rx_m_write_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_csr_arbitrator (
                                 // inputs:
                                  clk,
                                  cpu_data_master_address_to_slave,
                                  cpu_data_master_latency_counter,
                                  cpu_data_master_read,
                                  cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                  cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                  cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register,
                                  cpu_data_master_write,
                                  cpu_data_master_writedata,
                                  reset_n,
                                  sgdma_tx_csr_irq,
                                  sgdma_tx_csr_readdata,

                                 // outputs:
                                  cpu_data_master_granted_sgdma_tx_csr,
                                  cpu_data_master_qualified_request_sgdma_tx_csr,
                                  cpu_data_master_read_data_valid_sgdma_tx_csr,
                                  cpu_data_master_requests_sgdma_tx_csr,
                                  d1_sgdma_tx_csr_end_xfer,
                                  sgdma_tx_csr_address,
                                  sgdma_tx_csr_chipselect,
                                  sgdma_tx_csr_irq_from_sa,
                                  sgdma_tx_csr_read,
                                  sgdma_tx_csr_readdata_from_sa,
                                  sgdma_tx_csr_reset_n,
                                  sgdma_tx_csr_write,
                                  sgdma_tx_csr_writedata
                               )
;

  output           cpu_data_master_granted_sgdma_tx_csr;
  output           cpu_data_master_qualified_request_sgdma_tx_csr;
  output           cpu_data_master_read_data_valid_sgdma_tx_csr;
  output           cpu_data_master_requests_sgdma_tx_csr;
  output           d1_sgdma_tx_csr_end_xfer;
  output  [  3: 0] sgdma_tx_csr_address;
  output           sgdma_tx_csr_chipselect;
  output           sgdma_tx_csr_irq_from_sa;
  output           sgdma_tx_csr_read;
  output  [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  output           sgdma_tx_csr_reset_n;
  output           sgdma_tx_csr_write;
  output  [ 31: 0] sgdma_tx_csr_writedata;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input            sgdma_tx_csr_irq;
  input   [ 31: 0] sgdma_tx_csr_readdata;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_sgdma_tx_csr;
  wire             cpu_data_master_qualified_request_sgdma_tx_csr;
  wire             cpu_data_master_read_data_valid_sgdma_tx_csr;
  wire             cpu_data_master_requests_sgdma_tx_csr;
  wire             cpu_data_master_saved_grant_sgdma_tx_csr;
  reg              d1_reasons_to_wait;
  reg              d1_sgdma_tx_csr_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sgdma_tx_csr;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  3: 0] sgdma_tx_csr_address;
  wire             sgdma_tx_csr_allgrants;
  wire             sgdma_tx_csr_allow_new_arb_cycle;
  wire             sgdma_tx_csr_any_bursting_master_saved_grant;
  wire             sgdma_tx_csr_any_continuerequest;
  wire             sgdma_tx_csr_arb_counter_enable;
  reg              sgdma_tx_csr_arb_share_counter;
  wire             sgdma_tx_csr_arb_share_counter_next_value;
  wire             sgdma_tx_csr_arb_share_set_values;
  wire             sgdma_tx_csr_beginbursttransfer_internal;
  wire             sgdma_tx_csr_begins_xfer;
  wire             sgdma_tx_csr_chipselect;
  wire             sgdma_tx_csr_end_xfer;
  wire             sgdma_tx_csr_firsttransfer;
  wire             sgdma_tx_csr_grant_vector;
  wire             sgdma_tx_csr_in_a_read_cycle;
  wire             sgdma_tx_csr_in_a_write_cycle;
  wire             sgdma_tx_csr_irq_from_sa;
  wire             sgdma_tx_csr_master_qreq_vector;
  wire             sgdma_tx_csr_non_bursting_master_requests;
  wire             sgdma_tx_csr_read;
  wire    [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  reg              sgdma_tx_csr_reg_firsttransfer;
  wire             sgdma_tx_csr_reset_n;
  reg              sgdma_tx_csr_slavearbiterlockenable;
  wire             sgdma_tx_csr_slavearbiterlockenable2;
  wire             sgdma_tx_csr_unreg_firsttransfer;
  wire             sgdma_tx_csr_waits_for_read;
  wire             sgdma_tx_csr_waits_for_write;
  wire             sgdma_tx_csr_write;
  wire    [ 31: 0] sgdma_tx_csr_writedata;
  wire    [ 28: 0] shifted_address_to_sgdma_tx_csr_from_cpu_data_master;
  wire             wait_for_sgdma_tx_csr_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sgdma_tx_csr_end_xfer;
    end


  assign sgdma_tx_csr_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_sgdma_tx_csr));
  //assign sgdma_tx_csr_readdata_from_sa = sgdma_tx_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_tx_csr_readdata_from_sa = sgdma_tx_csr_readdata;

  assign cpu_data_master_requests_sgdma_tx_csr = ({cpu_data_master_address_to_slave[28 : 6] , 6'b0} == 29'h1002400) & (cpu_data_master_read | cpu_data_master_write);
  //sgdma_tx_csr_arb_share_counter set values, which is an e_mux
  assign sgdma_tx_csr_arb_share_set_values = 1;

  //sgdma_tx_csr_non_bursting_master_requests mux, which is an e_mux
  assign sgdma_tx_csr_non_bursting_master_requests = cpu_data_master_requests_sgdma_tx_csr;

  //sgdma_tx_csr_any_bursting_master_saved_grant mux, which is an e_mux
  assign sgdma_tx_csr_any_bursting_master_saved_grant = 0;

  //sgdma_tx_csr_arb_share_counter_next_value assignment, which is an e_assign
  assign sgdma_tx_csr_arb_share_counter_next_value = sgdma_tx_csr_firsttransfer ? (sgdma_tx_csr_arb_share_set_values - 1) : |sgdma_tx_csr_arb_share_counter ? (sgdma_tx_csr_arb_share_counter - 1) : 0;

  //sgdma_tx_csr_allgrants all slave grants, which is an e_mux
  assign sgdma_tx_csr_allgrants = |sgdma_tx_csr_grant_vector;

  //sgdma_tx_csr_end_xfer assignment, which is an e_assign
  assign sgdma_tx_csr_end_xfer = ~(sgdma_tx_csr_waits_for_read | sgdma_tx_csr_waits_for_write);

  //end_xfer_arb_share_counter_term_sgdma_tx_csr arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sgdma_tx_csr = sgdma_tx_csr_end_xfer & (~sgdma_tx_csr_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sgdma_tx_csr_arb_share_counter arbitration counter enable, which is an e_assign
  assign sgdma_tx_csr_arb_counter_enable = (end_xfer_arb_share_counter_term_sgdma_tx_csr & sgdma_tx_csr_allgrants) | (end_xfer_arb_share_counter_term_sgdma_tx_csr & ~sgdma_tx_csr_non_bursting_master_requests);

  //sgdma_tx_csr_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_csr_arb_share_counter <= 0;
      else if (sgdma_tx_csr_arb_counter_enable)
          sgdma_tx_csr_arb_share_counter <= sgdma_tx_csr_arb_share_counter_next_value;
    end


  //sgdma_tx_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_csr_slavearbiterlockenable <= 0;
      else if ((|sgdma_tx_csr_master_qreq_vector & end_xfer_arb_share_counter_term_sgdma_tx_csr) | (end_xfer_arb_share_counter_term_sgdma_tx_csr & ~sgdma_tx_csr_non_bursting_master_requests))
          sgdma_tx_csr_slavearbiterlockenable <= |sgdma_tx_csr_arb_share_counter_next_value;
    end


  //cpu/data_master sgdma_tx/csr arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = sgdma_tx_csr_slavearbiterlockenable & cpu_data_master_continuerequest;

  //sgdma_tx_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sgdma_tx_csr_slavearbiterlockenable2 = |sgdma_tx_csr_arb_share_counter_next_value;

  //cpu/data_master sgdma_tx/csr arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = sgdma_tx_csr_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //sgdma_tx_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sgdma_tx_csr_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_sgdma_tx_csr = cpu_data_master_requests_sgdma_tx_csr & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_sgdma_tx_csr, which is an e_mux
  assign cpu_data_master_read_data_valid_sgdma_tx_csr = cpu_data_master_granted_sgdma_tx_csr & cpu_data_master_read & ~sgdma_tx_csr_waits_for_read;

  //sgdma_tx_csr_writedata mux, which is an e_mux
  assign sgdma_tx_csr_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_sgdma_tx_csr = cpu_data_master_qualified_request_sgdma_tx_csr;

  //cpu/data_master saved-grant sgdma_tx/csr, which is an e_assign
  assign cpu_data_master_saved_grant_sgdma_tx_csr = cpu_data_master_requests_sgdma_tx_csr;

  //allow new arb cycle for sgdma_tx/csr, which is an e_assign
  assign sgdma_tx_csr_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sgdma_tx_csr_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sgdma_tx_csr_master_qreq_vector = 1;

  //sgdma_tx_csr_reset_n assignment, which is an e_assign
  assign sgdma_tx_csr_reset_n = reset_n;

  assign sgdma_tx_csr_chipselect = cpu_data_master_granted_sgdma_tx_csr;
  //sgdma_tx_csr_firsttransfer first transaction, which is an e_assign
  assign sgdma_tx_csr_firsttransfer = sgdma_tx_csr_begins_xfer ? sgdma_tx_csr_unreg_firsttransfer : sgdma_tx_csr_reg_firsttransfer;

  //sgdma_tx_csr_unreg_firsttransfer first transaction, which is an e_assign
  assign sgdma_tx_csr_unreg_firsttransfer = ~(sgdma_tx_csr_slavearbiterlockenable & sgdma_tx_csr_any_continuerequest);

  //sgdma_tx_csr_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_csr_reg_firsttransfer <= 1'b1;
      else if (sgdma_tx_csr_begins_xfer)
          sgdma_tx_csr_reg_firsttransfer <= sgdma_tx_csr_unreg_firsttransfer;
    end


  //sgdma_tx_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sgdma_tx_csr_beginbursttransfer_internal = sgdma_tx_csr_begins_xfer;

  //sgdma_tx_csr_read assignment, which is an e_mux
  assign sgdma_tx_csr_read = cpu_data_master_granted_sgdma_tx_csr & cpu_data_master_read;

  //sgdma_tx_csr_write assignment, which is an e_mux
  assign sgdma_tx_csr_write = cpu_data_master_granted_sgdma_tx_csr & cpu_data_master_write;

  assign shifted_address_to_sgdma_tx_csr_from_cpu_data_master = cpu_data_master_address_to_slave;
  //sgdma_tx_csr_address mux, which is an e_mux
  assign sgdma_tx_csr_address = shifted_address_to_sgdma_tx_csr_from_cpu_data_master >> 2;

  //d1_sgdma_tx_csr_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sgdma_tx_csr_end_xfer <= 1;
      else 
        d1_sgdma_tx_csr_end_xfer <= sgdma_tx_csr_end_xfer;
    end


  //sgdma_tx_csr_waits_for_read in a cycle, which is an e_mux
  assign sgdma_tx_csr_waits_for_read = sgdma_tx_csr_in_a_read_cycle & sgdma_tx_csr_begins_xfer;

  //sgdma_tx_csr_in_a_read_cycle assignment, which is an e_assign
  assign sgdma_tx_csr_in_a_read_cycle = cpu_data_master_granted_sgdma_tx_csr & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sgdma_tx_csr_in_a_read_cycle;

  //sgdma_tx_csr_waits_for_write in a cycle, which is an e_mux
  assign sgdma_tx_csr_waits_for_write = sgdma_tx_csr_in_a_write_cycle & 0;

  //sgdma_tx_csr_in_a_write_cycle assignment, which is an e_assign
  assign sgdma_tx_csr_in_a_write_cycle = cpu_data_master_granted_sgdma_tx_csr & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sgdma_tx_csr_in_a_write_cycle;

  assign wait_for_sgdma_tx_csr_counter = 0;
  //assign sgdma_tx_csr_irq_from_sa = sgdma_tx_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sgdma_tx_csr_irq_from_sa = sgdma_tx_csr_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx/csr enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_descriptor_read_arbitrator (
                                             // inputs:
                                              clk,
                                              d1_descriptor_memory_s1_end_xfer,
                                              descriptor_memory_s1_readdata_from_sa,
                                              reset_n,
                                              sgdma_tx_descriptor_read_address,
                                              sgdma_tx_descriptor_read_granted_descriptor_memory_s1,
                                              sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1,
                                              sgdma_tx_descriptor_read_read,
                                              sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1,
                                              sgdma_tx_descriptor_read_requests_descriptor_memory_s1,

                                             // outputs:
                                              sgdma_tx_descriptor_read_address_to_slave,
                                              sgdma_tx_descriptor_read_latency_counter,
                                              sgdma_tx_descriptor_read_readdata,
                                              sgdma_tx_descriptor_read_readdatavalid,
                                              sgdma_tx_descriptor_read_waitrequest
                                           )
;

  output  [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  output           sgdma_tx_descriptor_read_latency_counter;
  output  [ 31: 0] sgdma_tx_descriptor_read_readdata;
  output           sgdma_tx_descriptor_read_readdatavalid;
  output           sgdma_tx_descriptor_read_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s1_end_xfer;
  input   [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_descriptor_read_address;
  input            sgdma_tx_descriptor_read_granted_descriptor_memory_s1;
  input            sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;
  input            sgdma_tx_descriptor_read_read;
  input            sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;
  input            sgdma_tx_descriptor_read_requests_descriptor_memory_s1;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_sgdma_tx_descriptor_read_latency_counter;
  wire             pre_flush_sgdma_tx_descriptor_read_readdatavalid;
  wire             r_0;
  reg     [ 31: 0] sgdma_tx_descriptor_read_address_last_time;
  wire    [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  wire             sgdma_tx_descriptor_read_is_granted_some_slave;
  reg              sgdma_tx_descriptor_read_latency_counter;
  reg              sgdma_tx_descriptor_read_read_but_no_slave_selected;
  reg              sgdma_tx_descriptor_read_read_last_time;
  wire    [ 31: 0] sgdma_tx_descriptor_read_readdata;
  wire             sgdma_tx_descriptor_read_readdatavalid;
  wire             sgdma_tx_descriptor_read_run;
  wire             sgdma_tx_descriptor_read_waitrequest;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 | ~sgdma_tx_descriptor_read_requests_descriptor_memory_s1) & (sgdma_tx_descriptor_read_granted_descriptor_memory_s1 | ~sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1) & ((~sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 | ~(sgdma_tx_descriptor_read_read) | (1 & (sgdma_tx_descriptor_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_tx_descriptor_read_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_tx_descriptor_read_address_to_slave = {20'b1000000000000,
    sgdma_tx_descriptor_read_address[11 : 0]};

  //sgdma_tx_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_read_but_no_slave_selected <= 0;
      else 
        sgdma_tx_descriptor_read_read_but_no_slave_selected <= sgdma_tx_descriptor_read_read & sgdma_tx_descriptor_read_run & ~sgdma_tx_descriptor_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign sgdma_tx_descriptor_read_is_granted_some_slave = sgdma_tx_descriptor_read_granted_descriptor_memory_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_sgdma_tx_descriptor_read_readdatavalid = sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign sgdma_tx_descriptor_read_readdatavalid = sgdma_tx_descriptor_read_read_but_no_slave_selected |
    pre_flush_sgdma_tx_descriptor_read_readdatavalid;

  //sgdma_tx/descriptor_read readdata mux, which is an e_mux
  assign sgdma_tx_descriptor_read_readdata = descriptor_memory_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign sgdma_tx_descriptor_read_waitrequest = ~sgdma_tx_descriptor_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_latency_counter <= 0;
      else 
        sgdma_tx_descriptor_read_latency_counter <= p1_sgdma_tx_descriptor_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_sgdma_tx_descriptor_read_latency_counter = ((sgdma_tx_descriptor_read_run & sgdma_tx_descriptor_read_read))? latency_load_value :
    (sgdma_tx_descriptor_read_latency_counter)? sgdma_tx_descriptor_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {sgdma_tx_descriptor_read_requests_descriptor_memory_s1}} & 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx_descriptor_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_address_last_time <= 0;
      else 
        sgdma_tx_descriptor_read_address_last_time <= sgdma_tx_descriptor_read_address;
    end


  //sgdma_tx/descriptor_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_tx_descriptor_read_waitrequest & (sgdma_tx_descriptor_read_read);
    end


  //sgdma_tx_descriptor_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_read_address != sgdma_tx_descriptor_read_address_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_descriptor_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_read_read_last_time <= 0;
      else 
        sgdma_tx_descriptor_read_read_last_time <= sgdma_tx_descriptor_read_read;
    end


  //sgdma_tx_descriptor_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_read_read != sgdma_tx_descriptor_read_read_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_descriptor_write_arbitrator (
                                              // inputs:
                                               clk,
                                               d1_descriptor_memory_s1_end_xfer,
                                               reset_n,
                                               sgdma_tx_descriptor_write_address,
                                               sgdma_tx_descriptor_write_granted_descriptor_memory_s1,
                                               sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1,
                                               sgdma_tx_descriptor_write_requests_descriptor_memory_s1,
                                               sgdma_tx_descriptor_write_write,
                                               sgdma_tx_descriptor_write_writedata,

                                              // outputs:
                                               sgdma_tx_descriptor_write_address_to_slave,
                                               sgdma_tx_descriptor_write_waitrequest
                                            )
;

  output  [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  output           sgdma_tx_descriptor_write_waitrequest;
  input            clk;
  input            d1_descriptor_memory_s1_end_xfer;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_descriptor_write_address;
  input            sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  input            sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;
  input            sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
  input            sgdma_tx_descriptor_write_write;
  input   [ 31: 0] sgdma_tx_descriptor_write_writedata;

  reg              active_and_waiting_last_time;
  wire             r_0;
  reg     [ 31: 0] sgdma_tx_descriptor_write_address_last_time;
  wire    [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  wire             sgdma_tx_descriptor_write_run;
  wire             sgdma_tx_descriptor_write_waitrequest;
  reg              sgdma_tx_descriptor_write_write_last_time;
  reg     [ 31: 0] sgdma_tx_descriptor_write_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 | ~sgdma_tx_descriptor_write_requests_descriptor_memory_s1) & (sgdma_tx_descriptor_write_granted_descriptor_memory_s1 | ~sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1) & ((~sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 | ~(sgdma_tx_descriptor_write_write) | (1 & (sgdma_tx_descriptor_write_write))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_tx_descriptor_write_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_tx_descriptor_write_address_to_slave = {20'b1000000000000,
    sgdma_tx_descriptor_write_address[11 : 0]};

  //actual waitrequest port, which is an e_assign
  assign sgdma_tx_descriptor_write_waitrequest = ~sgdma_tx_descriptor_write_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx_descriptor_write_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_write_address_last_time <= 0;
      else 
        sgdma_tx_descriptor_write_address_last_time <= sgdma_tx_descriptor_write_address;
    end


  //sgdma_tx/descriptor_write waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_tx_descriptor_write_waitrequest & (sgdma_tx_descriptor_write_write);
    end


  //sgdma_tx_descriptor_write_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_write_address != sgdma_tx_descriptor_write_address_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_write_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_descriptor_write_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_write_write_last_time <= 0;
      else 
        sgdma_tx_descriptor_write_write_last_time <= sgdma_tx_descriptor_write_write;
    end


  //sgdma_tx_descriptor_write_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_write_write != sgdma_tx_descriptor_write_write_last_time))
        begin
          $write("%0d ns: sgdma_tx_descriptor_write_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_descriptor_write_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_descriptor_write_writedata_last_time <= 0;
      else 
        sgdma_tx_descriptor_write_writedata_last_time <= sgdma_tx_descriptor_write_writedata;
    end


  //sgdma_tx_descriptor_write_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_descriptor_write_writedata != sgdma_tx_descriptor_write_writedata_last_time) & sgdma_tx_descriptor_write_write)
        begin
          $write("%0d ns: sgdma_tx_descriptor_write_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_m_read_arbitrator (
                                    // inputs:
                                     clk,
                                     cpu_ddr_clock_bridge_s1_readdata_from_sa,
                                     cpu_ddr_clock_bridge_s1_waitrequest_from_sa,
                                     d1_cpu_ddr_clock_bridge_s1_end_xfer,
                                     reset_n,
                                     sgdma_tx_m_read_address,
                                     sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1,
                                     sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1,
                                     sgdma_tx_m_read_read,
                                     sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1,
                                     sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                     sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1,

                                    // outputs:
                                     sgdma_tx_m_read_address_to_slave,
                                     sgdma_tx_m_read_latency_counter,
                                     sgdma_tx_m_read_readdata,
                                     sgdma_tx_m_read_readdatavalid,
                                     sgdma_tx_m_read_waitrequest
                                  )
;

  output  [ 31: 0] sgdma_tx_m_read_address_to_slave;
  output           sgdma_tx_m_read_latency_counter;
  output  [ 31: 0] sgdma_tx_m_read_readdata;
  output           sgdma_tx_m_read_readdatavalid;
  output           sgdma_tx_m_read_waitrequest;
  input            clk;
  input   [ 31: 0] cpu_ddr_clock_bridge_s1_readdata_from_sa;
  input            cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  input            d1_cpu_ddr_clock_bridge_s1_end_xfer;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_m_read_address;
  input            sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1;
  input            sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1;
  input            sgdma_tx_m_read_read;
  input            sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1;
  input            sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_sgdma_tx_m_read_latency_counter;
  wire             pre_flush_sgdma_tx_m_read_readdatavalid;
  wire             r_0;
  reg     [ 31: 0] sgdma_tx_m_read_address_last_time;
  wire    [ 31: 0] sgdma_tx_m_read_address_to_slave;
  wire             sgdma_tx_m_read_is_granted_some_slave;
  reg              sgdma_tx_m_read_latency_counter;
  reg              sgdma_tx_m_read_read_but_no_slave_selected;
  reg              sgdma_tx_m_read_read_last_time;
  wire    [ 31: 0] sgdma_tx_m_read_readdata;
  wire             sgdma_tx_m_read_readdatavalid;
  wire             sgdma_tx_m_read_run;
  wire             sgdma_tx_m_read_waitrequest;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1 | ~sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1) & (sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1 | ~sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1) & ((~sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1 | ~(sgdma_tx_m_read_read) | (1 & ~cpu_ddr_clock_bridge_s1_waitrequest_from_sa & (sgdma_tx_m_read_read))));

  //cascaded wait assignment, which is an e_assign
  assign sgdma_tx_m_read_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign sgdma_tx_m_read_address_to_slave = {6'b111,
    sgdma_tx_m_read_address[25 : 0]};

  //sgdma_tx_m_read_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_read_but_no_slave_selected <= 0;
      else 
        sgdma_tx_m_read_read_but_no_slave_selected <= sgdma_tx_m_read_read & sgdma_tx_m_read_run & ~sgdma_tx_m_read_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign sgdma_tx_m_read_is_granted_some_slave = sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_sgdma_tx_m_read_readdatavalid = sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign sgdma_tx_m_read_readdatavalid = sgdma_tx_m_read_read_but_no_slave_selected |
    pre_flush_sgdma_tx_m_read_readdatavalid;

  //sgdma_tx/m_read readdata mux, which is an e_mux
  assign sgdma_tx_m_read_readdata = cpu_ddr_clock_bridge_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign sgdma_tx_m_read_waitrequest = ~sgdma_tx_m_read_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_latency_counter <= 0;
      else 
        sgdma_tx_m_read_latency_counter <= p1_sgdma_tx_m_read_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_sgdma_tx_m_read_latency_counter = ((sgdma_tx_m_read_run & sgdma_tx_m_read_read))? latency_load_value :
    (sgdma_tx_m_read_latency_counter)? sgdma_tx_m_read_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sgdma_tx_m_read_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_address_last_time <= 0;
      else 
        sgdma_tx_m_read_address_last_time <= sgdma_tx_m_read_address;
    end


  //sgdma_tx/m_read waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= sgdma_tx_m_read_waitrequest & (sgdma_tx_m_read_read);
    end


  //sgdma_tx_m_read_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_m_read_address != sgdma_tx_m_read_address_last_time))
        begin
          $write("%0d ns: sgdma_tx_m_read_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //sgdma_tx_m_read_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sgdma_tx_m_read_read_last_time <= 0;
      else 
        sgdma_tx_m_read_read_last_time <= sgdma_tx_m_read_read;
    end


  //sgdma_tx_m_read_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (sgdma_tx_m_read_read != sgdma_tx_m_read_read_last_time))
        begin
          $write("%0d ns: sgdma_tx_m_read_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sgdma_tx_out_arbitrator (
                                 // inputs:
                                  clk,
                                  reset_n,
                                  sgdma_tx_out_data,
                                  sgdma_tx_out_empty,
                                  sgdma_tx_out_endofpacket,
                                  sgdma_tx_out_error,
                                  sgdma_tx_out_startofpacket,
                                  sgdma_tx_out_valid,
                                  tse_mac_transmit_ready_from_sa,

                                 // outputs:
                                  sgdma_tx_out_ready
                               )
;

  output           sgdma_tx_out_ready;
  input            clk;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_out_data;
  input   [  1: 0] sgdma_tx_out_empty;
  input            sgdma_tx_out_endofpacket;
  input            sgdma_tx_out_error;
  input            sgdma_tx_out_startofpacket;
  input            sgdma_tx_out_valid;
  input            tse_mac_transmit_ready_from_sa;

  wire             sgdma_tx_out_ready;
  //mux sgdma_tx_out_ready, which is an e_mux
  assign sgdma_tx_out_ready = tse_mac_transmit_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_slow_peripheral_bridge_s1_module (
                                                                          // inputs:
                                                                           clear_fifo,
                                                                           clk,
                                                                           data_in,
                                                                           read,
                                                                           reset_n,
                                                                           sync_reset,
                                                                           write,

                                                                          // outputs:
                                                                           data_out,
                                                                           empty,
                                                                           fifo_contains_ones_n,
                                                                           full
                                                                        )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  reg              full_18;
  reg              full_19;
  reg              full_2;
  reg              full_20;
  reg              full_21;
  reg              full_22;
  reg              full_23;
  reg              full_24;
  reg              full_25;
  reg              full_26;
  reg              full_27;
  reg              full_28;
  reg              full_29;
  reg              full_3;
  reg              full_30;
  reg              full_31;
  reg              full_32;
  wire             full_33;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  6: 0] how_many_ones;
  wire    [  6: 0] one_count_minus_one;
  wire    [  6: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p18_full_18;
  wire             p18_stage_18;
  wire             p19_full_19;
  wire             p19_stage_19;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p20_full_20;
  wire             p20_stage_20;
  wire             p21_full_21;
  wire             p21_stage_21;
  wire             p22_full_22;
  wire             p22_stage_22;
  wire             p23_full_23;
  wire             p23_stage_23;
  wire             p24_full_24;
  wire             p24_stage_24;
  wire             p25_full_25;
  wire             p25_stage_25;
  wire             p26_full_26;
  wire             p26_stage_26;
  wire             p27_full_27;
  wire             p27_stage_27;
  wire             p28_full_28;
  wire             p28_stage_28;
  wire             p29_full_29;
  wire             p29_stage_29;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p30_full_30;
  wire             p30_stage_30;
  wire             p31_full_31;
  wire             p31_stage_31;
  wire             p32_full_32;
  wire             p32_stage_32;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_18;
  reg              stage_19;
  reg              stage_2;
  reg              stage_20;
  reg              stage_21;
  reg              stage_22;
  reg              stage_23;
  reg              stage_24;
  reg              stage_25;
  reg              stage_26;
  reg              stage_27;
  reg              stage_28;
  reg              stage_29;
  reg              stage_3;
  reg              stage_30;
  reg              stage_31;
  reg              stage_32;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  6: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_32;
  assign empty = !full_0;
  assign full_33 = 0;
  //data_32, which is an e_mux
  assign p32_stage_32 = ((full_33 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_32 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_32))
          if (sync_reset & full_32 & !((full_33 == 0) & read & write))
              stage_32 <= 0;
          else 
            stage_32 <= p32_stage_32;
    end


  //control_32, which is an e_mux
  assign p32_full_32 = ((read & !write) == 0)? full_31 :
    0;

  //control_reg_32, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_32 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_32 <= 0;
          else 
            full_32 <= p32_full_32;
    end


  //data_31, which is an e_mux
  assign p31_stage_31 = ((full_32 & ~clear_fifo) == 0)? data_in :
    stage_32;

  //data_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_31 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_31))
          if (sync_reset & full_31 & !((full_32 == 0) & read & write))
              stage_31 <= 0;
          else 
            stage_31 <= p31_stage_31;
    end


  //control_31, which is an e_mux
  assign p31_full_31 = ((read & !write) == 0)? full_30 :
    full_32;

  //control_reg_31, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_31 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_31 <= 0;
          else 
            full_31 <= p31_full_31;
    end


  //data_30, which is an e_mux
  assign p30_stage_30 = ((full_31 & ~clear_fifo) == 0)? data_in :
    stage_31;

  //data_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_30 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_30))
          if (sync_reset & full_30 & !((full_31 == 0) & read & write))
              stage_30 <= 0;
          else 
            stage_30 <= p30_stage_30;
    end


  //control_30, which is an e_mux
  assign p30_full_30 = ((read & !write) == 0)? full_29 :
    full_31;

  //control_reg_30, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_30 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_30 <= 0;
          else 
            full_30 <= p30_full_30;
    end


  //data_29, which is an e_mux
  assign p29_stage_29 = ((full_30 & ~clear_fifo) == 0)? data_in :
    stage_30;

  //data_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_29 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_29))
          if (sync_reset & full_29 & !((full_30 == 0) & read & write))
              stage_29 <= 0;
          else 
            stage_29 <= p29_stage_29;
    end


  //control_29, which is an e_mux
  assign p29_full_29 = ((read & !write) == 0)? full_28 :
    full_30;

  //control_reg_29, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_29 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_29 <= 0;
          else 
            full_29 <= p29_full_29;
    end


  //data_28, which is an e_mux
  assign p28_stage_28 = ((full_29 & ~clear_fifo) == 0)? data_in :
    stage_29;

  //data_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_28 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_28))
          if (sync_reset & full_28 & !((full_29 == 0) & read & write))
              stage_28 <= 0;
          else 
            stage_28 <= p28_stage_28;
    end


  //control_28, which is an e_mux
  assign p28_full_28 = ((read & !write) == 0)? full_27 :
    full_29;

  //control_reg_28, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_28 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_28 <= 0;
          else 
            full_28 <= p28_full_28;
    end


  //data_27, which is an e_mux
  assign p27_stage_27 = ((full_28 & ~clear_fifo) == 0)? data_in :
    stage_28;

  //data_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_27 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_27))
          if (sync_reset & full_27 & !((full_28 == 0) & read & write))
              stage_27 <= 0;
          else 
            stage_27 <= p27_stage_27;
    end


  //control_27, which is an e_mux
  assign p27_full_27 = ((read & !write) == 0)? full_26 :
    full_28;

  //control_reg_27, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_27 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_27 <= 0;
          else 
            full_27 <= p27_full_27;
    end


  //data_26, which is an e_mux
  assign p26_stage_26 = ((full_27 & ~clear_fifo) == 0)? data_in :
    stage_27;

  //data_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_26 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_26))
          if (sync_reset & full_26 & !((full_27 == 0) & read & write))
              stage_26 <= 0;
          else 
            stage_26 <= p26_stage_26;
    end


  //control_26, which is an e_mux
  assign p26_full_26 = ((read & !write) == 0)? full_25 :
    full_27;

  //control_reg_26, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_26 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_26 <= 0;
          else 
            full_26 <= p26_full_26;
    end


  //data_25, which is an e_mux
  assign p25_stage_25 = ((full_26 & ~clear_fifo) == 0)? data_in :
    stage_26;

  //data_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_25 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_25))
          if (sync_reset & full_25 & !((full_26 == 0) & read & write))
              stage_25 <= 0;
          else 
            stage_25 <= p25_stage_25;
    end


  //control_25, which is an e_mux
  assign p25_full_25 = ((read & !write) == 0)? full_24 :
    full_26;

  //control_reg_25, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_25 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_25 <= 0;
          else 
            full_25 <= p25_full_25;
    end


  //data_24, which is an e_mux
  assign p24_stage_24 = ((full_25 & ~clear_fifo) == 0)? data_in :
    stage_25;

  //data_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_24 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_24))
          if (sync_reset & full_24 & !((full_25 == 0) & read & write))
              stage_24 <= 0;
          else 
            stage_24 <= p24_stage_24;
    end


  //control_24, which is an e_mux
  assign p24_full_24 = ((read & !write) == 0)? full_23 :
    full_25;

  //control_reg_24, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_24 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_24 <= 0;
          else 
            full_24 <= p24_full_24;
    end


  //data_23, which is an e_mux
  assign p23_stage_23 = ((full_24 & ~clear_fifo) == 0)? data_in :
    stage_24;

  //data_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_23 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_23))
          if (sync_reset & full_23 & !((full_24 == 0) & read & write))
              stage_23 <= 0;
          else 
            stage_23 <= p23_stage_23;
    end


  //control_23, which is an e_mux
  assign p23_full_23 = ((read & !write) == 0)? full_22 :
    full_24;

  //control_reg_23, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_23 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_23 <= 0;
          else 
            full_23 <= p23_full_23;
    end


  //data_22, which is an e_mux
  assign p22_stage_22 = ((full_23 & ~clear_fifo) == 0)? data_in :
    stage_23;

  //data_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_22 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_22))
          if (sync_reset & full_22 & !((full_23 == 0) & read & write))
              stage_22 <= 0;
          else 
            stage_22 <= p22_stage_22;
    end


  //control_22, which is an e_mux
  assign p22_full_22 = ((read & !write) == 0)? full_21 :
    full_23;

  //control_reg_22, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_22 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_22 <= 0;
          else 
            full_22 <= p22_full_22;
    end


  //data_21, which is an e_mux
  assign p21_stage_21 = ((full_22 & ~clear_fifo) == 0)? data_in :
    stage_22;

  //data_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_21 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_21))
          if (sync_reset & full_21 & !((full_22 == 0) & read & write))
              stage_21 <= 0;
          else 
            stage_21 <= p21_stage_21;
    end


  //control_21, which is an e_mux
  assign p21_full_21 = ((read & !write) == 0)? full_20 :
    full_22;

  //control_reg_21, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_21 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_21 <= 0;
          else 
            full_21 <= p21_full_21;
    end


  //data_20, which is an e_mux
  assign p20_stage_20 = ((full_21 & ~clear_fifo) == 0)? data_in :
    stage_21;

  //data_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_20 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_20))
          if (sync_reset & full_20 & !((full_21 == 0) & read & write))
              stage_20 <= 0;
          else 
            stage_20 <= p20_stage_20;
    end


  //control_20, which is an e_mux
  assign p20_full_20 = ((read & !write) == 0)? full_19 :
    full_21;

  //control_reg_20, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_20 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_20 <= 0;
          else 
            full_20 <= p20_full_20;
    end


  //data_19, which is an e_mux
  assign p19_stage_19 = ((full_20 & ~clear_fifo) == 0)? data_in :
    stage_20;

  //data_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_19 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_19))
          if (sync_reset & full_19 & !((full_20 == 0) & read & write))
              stage_19 <= 0;
          else 
            stage_19 <= p19_stage_19;
    end


  //control_19, which is an e_mux
  assign p19_full_19 = ((read & !write) == 0)? full_18 :
    full_20;

  //control_reg_19, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_19 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_19 <= 0;
          else 
            full_19 <= p19_full_19;
    end


  //data_18, which is an e_mux
  assign p18_stage_18 = ((full_19 & ~clear_fifo) == 0)? data_in :
    stage_19;

  //data_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_18 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_18))
          if (sync_reset & full_18 & !((full_19 == 0) & read & write))
              stage_18 <= 0;
          else 
            stage_18 <= p18_stage_18;
    end


  //control_18, which is an e_mux
  assign p18_full_18 = ((read & !write) == 0)? full_17 :
    full_19;

  //control_reg_18, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_18 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_18 <= 0;
          else 
            full_18 <= p18_full_18;
    end


  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    stage_18;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    full_18;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module slow_peripheral_bridge_s1_arbitrator (
                                              // inputs:
                                               clk,
                                               cpu_data_master_address_to_slave,
                                               cpu_data_master_byteenable,
                                               cpu_data_master_latency_counter,
                                               cpu_data_master_read,
                                               cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                               cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                               cpu_data_master_write,
                                               cpu_data_master_writedata,
                                               reset_n,
                                               slow_peripheral_bridge_s1_endofpacket,
                                               slow_peripheral_bridge_s1_readdata,
                                               slow_peripheral_bridge_s1_readdatavalid,
                                               slow_peripheral_bridge_s1_waitrequest,

                                              // outputs:
                                               cpu_data_master_granted_slow_peripheral_bridge_s1,
                                               cpu_data_master_qualified_request_slow_peripheral_bridge_s1,
                                               cpu_data_master_read_data_valid_slow_peripheral_bridge_s1,
                                               cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register,
                                               cpu_data_master_requests_slow_peripheral_bridge_s1,
                                               d1_slow_peripheral_bridge_s1_end_xfer,
                                               slow_peripheral_bridge_s1_address,
                                               slow_peripheral_bridge_s1_byteenable,
                                               slow_peripheral_bridge_s1_endofpacket_from_sa,
                                               slow_peripheral_bridge_s1_nativeaddress,
                                               slow_peripheral_bridge_s1_read,
                                               slow_peripheral_bridge_s1_readdata_from_sa,
                                               slow_peripheral_bridge_s1_reset_n,
                                               slow_peripheral_bridge_s1_waitrequest_from_sa,
                                               slow_peripheral_bridge_s1_write,
                                               slow_peripheral_bridge_s1_writedata
                                            )
;

  output           cpu_data_master_granted_slow_peripheral_bridge_s1;
  output           cpu_data_master_qualified_request_slow_peripheral_bridge_s1;
  output           cpu_data_master_read_data_valid_slow_peripheral_bridge_s1;
  output           cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  output           cpu_data_master_requests_slow_peripheral_bridge_s1;
  output           d1_slow_peripheral_bridge_s1_end_xfer;
  output  [  5: 0] slow_peripheral_bridge_s1_address;
  output  [  3: 0] slow_peripheral_bridge_s1_byteenable;
  output           slow_peripheral_bridge_s1_endofpacket_from_sa;
  output  [  5: 0] slow_peripheral_bridge_s1_nativeaddress;
  output           slow_peripheral_bridge_s1_read;
  output  [ 31: 0] slow_peripheral_bridge_s1_readdata_from_sa;
  output           slow_peripheral_bridge_s1_reset_n;
  output           slow_peripheral_bridge_s1_waitrequest_from_sa;
  output           slow_peripheral_bridge_s1_write;
  output  [ 31: 0] slow_peripheral_bridge_s1_writedata;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input            slow_peripheral_bridge_s1_endofpacket;
  input   [ 31: 0] slow_peripheral_bridge_s1_readdata;
  input            slow_peripheral_bridge_s1_readdatavalid;
  input            slow_peripheral_bridge_s1_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_slow_peripheral_bridge_s1;
  wire             cpu_data_master_qualified_request_slow_peripheral_bridge_s1;
  wire             cpu_data_master_rdv_fifo_empty_slow_peripheral_bridge_s1;
  wire             cpu_data_master_rdv_fifo_output_from_slow_peripheral_bridge_s1;
  wire             cpu_data_master_read_data_valid_slow_peripheral_bridge_s1;
  wire             cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  wire             cpu_data_master_requests_slow_peripheral_bridge_s1;
  wire             cpu_data_master_saved_grant_slow_peripheral_bridge_s1;
  reg              d1_reasons_to_wait;
  reg              d1_slow_peripheral_bridge_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_slow_peripheral_bridge_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 28: 0] shifted_address_to_slow_peripheral_bridge_s1_from_cpu_data_master;
  wire    [  5: 0] slow_peripheral_bridge_s1_address;
  wire             slow_peripheral_bridge_s1_allgrants;
  wire             slow_peripheral_bridge_s1_allow_new_arb_cycle;
  wire             slow_peripheral_bridge_s1_any_bursting_master_saved_grant;
  wire             slow_peripheral_bridge_s1_any_continuerequest;
  wire             slow_peripheral_bridge_s1_arb_counter_enable;
  reg              slow_peripheral_bridge_s1_arb_share_counter;
  wire             slow_peripheral_bridge_s1_arb_share_counter_next_value;
  wire             slow_peripheral_bridge_s1_arb_share_set_values;
  wire             slow_peripheral_bridge_s1_beginbursttransfer_internal;
  wire             slow_peripheral_bridge_s1_begins_xfer;
  wire    [  3: 0] slow_peripheral_bridge_s1_byteenable;
  wire             slow_peripheral_bridge_s1_end_xfer;
  wire             slow_peripheral_bridge_s1_endofpacket_from_sa;
  wire             slow_peripheral_bridge_s1_firsttransfer;
  wire             slow_peripheral_bridge_s1_grant_vector;
  wire             slow_peripheral_bridge_s1_in_a_read_cycle;
  wire             slow_peripheral_bridge_s1_in_a_write_cycle;
  wire             slow_peripheral_bridge_s1_master_qreq_vector;
  wire             slow_peripheral_bridge_s1_move_on_to_next_transaction;
  wire    [  5: 0] slow_peripheral_bridge_s1_nativeaddress;
  wire             slow_peripheral_bridge_s1_non_bursting_master_requests;
  wire             slow_peripheral_bridge_s1_read;
  wire    [ 31: 0] slow_peripheral_bridge_s1_readdata_from_sa;
  wire             slow_peripheral_bridge_s1_readdatavalid_from_sa;
  reg              slow_peripheral_bridge_s1_reg_firsttransfer;
  wire             slow_peripheral_bridge_s1_reset_n;
  reg              slow_peripheral_bridge_s1_slavearbiterlockenable;
  wire             slow_peripheral_bridge_s1_slavearbiterlockenable2;
  wire             slow_peripheral_bridge_s1_unreg_firsttransfer;
  wire             slow_peripheral_bridge_s1_waitrequest_from_sa;
  wire             slow_peripheral_bridge_s1_waits_for_read;
  wire             slow_peripheral_bridge_s1_waits_for_write;
  wire             slow_peripheral_bridge_s1_write;
  wire    [ 31: 0] slow_peripheral_bridge_s1_writedata;
  wire             wait_for_slow_peripheral_bridge_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~slow_peripheral_bridge_s1_end_xfer;
    end


  assign slow_peripheral_bridge_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_slow_peripheral_bridge_s1));
  //assign slow_peripheral_bridge_s1_readdatavalid_from_sa = slow_peripheral_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign slow_peripheral_bridge_s1_readdatavalid_from_sa = slow_peripheral_bridge_s1_readdatavalid;

  //assign slow_peripheral_bridge_s1_readdata_from_sa = slow_peripheral_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign slow_peripheral_bridge_s1_readdata_from_sa = slow_peripheral_bridge_s1_readdata;

  assign cpu_data_master_requests_slow_peripheral_bridge_s1 = ({cpu_data_master_address_to_slave[28 : 8] , 8'b0} == 29'h0) & (cpu_data_master_read | cpu_data_master_write);
  //assign slow_peripheral_bridge_s1_waitrequest_from_sa = slow_peripheral_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign slow_peripheral_bridge_s1_waitrequest_from_sa = slow_peripheral_bridge_s1_waitrequest;

  //slow_peripheral_bridge_s1_arb_share_counter set values, which is an e_mux
  assign slow_peripheral_bridge_s1_arb_share_set_values = 1;

  //slow_peripheral_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  assign slow_peripheral_bridge_s1_non_bursting_master_requests = cpu_data_master_requests_slow_peripheral_bridge_s1;

  //slow_peripheral_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign slow_peripheral_bridge_s1_any_bursting_master_saved_grant = 0;

  //slow_peripheral_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign slow_peripheral_bridge_s1_arb_share_counter_next_value = slow_peripheral_bridge_s1_firsttransfer ? (slow_peripheral_bridge_s1_arb_share_set_values - 1) : |slow_peripheral_bridge_s1_arb_share_counter ? (slow_peripheral_bridge_s1_arb_share_counter - 1) : 0;

  //slow_peripheral_bridge_s1_allgrants all slave grants, which is an e_mux
  assign slow_peripheral_bridge_s1_allgrants = |slow_peripheral_bridge_s1_grant_vector;

  //slow_peripheral_bridge_s1_end_xfer assignment, which is an e_assign
  assign slow_peripheral_bridge_s1_end_xfer = ~(slow_peripheral_bridge_s1_waits_for_read | slow_peripheral_bridge_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_slow_peripheral_bridge_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_slow_peripheral_bridge_s1 = slow_peripheral_bridge_s1_end_xfer & (~slow_peripheral_bridge_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //slow_peripheral_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign slow_peripheral_bridge_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_slow_peripheral_bridge_s1 & slow_peripheral_bridge_s1_allgrants) | (end_xfer_arb_share_counter_term_slow_peripheral_bridge_s1 & ~slow_peripheral_bridge_s1_non_bursting_master_requests);

  //slow_peripheral_bridge_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_s1_arb_share_counter <= 0;
      else if (slow_peripheral_bridge_s1_arb_counter_enable)
          slow_peripheral_bridge_s1_arb_share_counter <= slow_peripheral_bridge_s1_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_s1_slavearbiterlockenable <= 0;
      else if ((|slow_peripheral_bridge_s1_master_qreq_vector & end_xfer_arb_share_counter_term_slow_peripheral_bridge_s1) | (end_xfer_arb_share_counter_term_slow_peripheral_bridge_s1 & ~slow_peripheral_bridge_s1_non_bursting_master_requests))
          slow_peripheral_bridge_s1_slavearbiterlockenable <= |slow_peripheral_bridge_s1_arb_share_counter_next_value;
    end


  //cpu/data_master slow_peripheral_bridge/s1 arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = slow_peripheral_bridge_s1_slavearbiterlockenable & cpu_data_master_continuerequest;

  //slow_peripheral_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_s1_slavearbiterlockenable2 = |slow_peripheral_bridge_s1_arb_share_counter_next_value;

  //cpu/data_master slow_peripheral_bridge/s1 arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = slow_peripheral_bridge_s1_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //slow_peripheral_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign slow_peripheral_bridge_s1_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_slow_peripheral_bridge_s1 = cpu_data_master_requests_slow_peripheral_bridge_s1 & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register))));
  //unique name for slow_peripheral_bridge_s1_move_on_to_next_transaction, which is an e_assign
  assign slow_peripheral_bridge_s1_move_on_to_next_transaction = slow_peripheral_bridge_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_slow_peripheral_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_slow_peripheral_bridge_s1_module rdv_fifo_for_cpu_data_master_to_slow_peripheral_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_slow_peripheral_bridge_s1),
      .data_out             (cpu_data_master_rdv_fifo_output_from_slow_peripheral_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_slow_peripheral_bridge_s1),
      .full                 (),
      .read                 (slow_peripheral_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~slow_peripheral_bridge_s1_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register = ~cpu_data_master_rdv_fifo_empty_slow_peripheral_bridge_s1;
  //local readdatavalid cpu_data_master_read_data_valid_slow_peripheral_bridge_s1, which is an e_mux
  assign cpu_data_master_read_data_valid_slow_peripheral_bridge_s1 = slow_peripheral_bridge_s1_readdatavalid_from_sa;

  //slow_peripheral_bridge_s1_writedata mux, which is an e_mux
  assign slow_peripheral_bridge_s1_writedata = cpu_data_master_writedata;

  //assign slow_peripheral_bridge_s1_endofpacket_from_sa = slow_peripheral_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign slow_peripheral_bridge_s1_endofpacket_from_sa = slow_peripheral_bridge_s1_endofpacket;

  //master is always granted when requested
  assign cpu_data_master_granted_slow_peripheral_bridge_s1 = cpu_data_master_qualified_request_slow_peripheral_bridge_s1;

  //cpu/data_master saved-grant slow_peripheral_bridge/s1, which is an e_assign
  assign cpu_data_master_saved_grant_slow_peripheral_bridge_s1 = cpu_data_master_requests_slow_peripheral_bridge_s1;

  //allow new arb cycle for slow_peripheral_bridge/s1, which is an e_assign
  assign slow_peripheral_bridge_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign slow_peripheral_bridge_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign slow_peripheral_bridge_s1_master_qreq_vector = 1;

  //slow_peripheral_bridge_s1_reset_n assignment, which is an e_assign
  assign slow_peripheral_bridge_s1_reset_n = reset_n;

  //slow_peripheral_bridge_s1_firsttransfer first transaction, which is an e_assign
  assign slow_peripheral_bridge_s1_firsttransfer = slow_peripheral_bridge_s1_begins_xfer ? slow_peripheral_bridge_s1_unreg_firsttransfer : slow_peripheral_bridge_s1_reg_firsttransfer;

  //slow_peripheral_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign slow_peripheral_bridge_s1_unreg_firsttransfer = ~(slow_peripheral_bridge_s1_slavearbiterlockenable & slow_peripheral_bridge_s1_any_continuerequest);

  //slow_peripheral_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_s1_reg_firsttransfer <= 1'b1;
      else if (slow_peripheral_bridge_s1_begins_xfer)
          slow_peripheral_bridge_s1_reg_firsttransfer <= slow_peripheral_bridge_s1_unreg_firsttransfer;
    end


  //slow_peripheral_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign slow_peripheral_bridge_s1_beginbursttransfer_internal = slow_peripheral_bridge_s1_begins_xfer;

  //slow_peripheral_bridge_s1_read assignment, which is an e_mux
  assign slow_peripheral_bridge_s1_read = cpu_data_master_granted_slow_peripheral_bridge_s1 & cpu_data_master_read;

  //slow_peripheral_bridge_s1_write assignment, which is an e_mux
  assign slow_peripheral_bridge_s1_write = cpu_data_master_granted_slow_peripheral_bridge_s1 & cpu_data_master_write;

  assign shifted_address_to_slow_peripheral_bridge_s1_from_cpu_data_master = cpu_data_master_address_to_slave;
  //slow_peripheral_bridge_s1_address mux, which is an e_mux
  assign slow_peripheral_bridge_s1_address = shifted_address_to_slow_peripheral_bridge_s1_from_cpu_data_master >> 2;

  //slaveid slow_peripheral_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign slow_peripheral_bridge_s1_nativeaddress = cpu_data_master_address_to_slave >> 2;

  //d1_slow_peripheral_bridge_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_slow_peripheral_bridge_s1_end_xfer <= 1;
      else 
        d1_slow_peripheral_bridge_s1_end_xfer <= slow_peripheral_bridge_s1_end_xfer;
    end


  //slow_peripheral_bridge_s1_waits_for_read in a cycle, which is an e_mux
  assign slow_peripheral_bridge_s1_waits_for_read = slow_peripheral_bridge_s1_in_a_read_cycle & slow_peripheral_bridge_s1_waitrequest_from_sa;

  //slow_peripheral_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  assign slow_peripheral_bridge_s1_in_a_read_cycle = cpu_data_master_granted_slow_peripheral_bridge_s1 & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = slow_peripheral_bridge_s1_in_a_read_cycle;

  //slow_peripheral_bridge_s1_waits_for_write in a cycle, which is an e_mux
  assign slow_peripheral_bridge_s1_waits_for_write = slow_peripheral_bridge_s1_in_a_write_cycle & slow_peripheral_bridge_s1_waitrequest_from_sa;

  //slow_peripheral_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  assign slow_peripheral_bridge_s1_in_a_write_cycle = cpu_data_master_granted_slow_peripheral_bridge_s1 & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = slow_peripheral_bridge_s1_in_a_write_cycle;

  assign wait_for_slow_peripheral_bridge_s1_counter = 0;
  //slow_peripheral_bridge_s1_byteenable byte enable port mux, which is an e_mux
  assign slow_peripheral_bridge_s1_byteenable = (cpu_data_master_granted_slow_peripheral_bridge_s1)? cpu_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //slow_peripheral_bridge/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module slow_peripheral_bridge_m1_arbitrator (
                                              // inputs:
                                               button_pio_s1_readdata_from_sa,
                                               clk,
                                               cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa,
                                               cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa,
                                               cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa,
                                               cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa,
                                               cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa,
                                               cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa,
                                               cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa,
                                               cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa,
                                               cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa,
                                               d1_button_pio_s1_end_xfer,
                                               d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer,
                                               d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer,
                                               d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer,
                                               d1_high_res_timer_s1_end_xfer,
                                               d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                               d1_led_pio_s1_end_xfer,
                                               d1_performance_counter_control_slave_end_xfer,
                                               d1_sys_clk_timer_s1_end_xfer,
                                               d1_sysid_control_slave_end_xfer,
                                               high_res_timer_s1_readdata_from_sa,
                                               jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                               jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                               led_pio_s1_readdata_from_sa,
                                               performance_counter_control_slave_readdata_from_sa,
                                               reset_n,
                                               slow_peripheral_bridge_m1_address,
                                               slow_peripheral_bridge_m1_byteenable,
                                               slow_peripheral_bridge_m1_granted_button_pio_s1,
                                               slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in,
                                               slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in,
                                               slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in,
                                               slow_peripheral_bridge_m1_granted_high_res_timer_s1,
                                               slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave,
                                               slow_peripheral_bridge_m1_granted_led_pio_s1,
                                               slow_peripheral_bridge_m1_granted_performance_counter_control_slave,
                                               slow_peripheral_bridge_m1_granted_sys_clk_timer_s1,
                                               slow_peripheral_bridge_m1_granted_sysid_control_slave,
                                               slow_peripheral_bridge_m1_qualified_request_button_pio_s1,
                                               slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in,
                                               slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in,
                                               slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in,
                                               slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1,
                                               slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave,
                                               slow_peripheral_bridge_m1_qualified_request_led_pio_s1,
                                               slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave,
                                               slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1,
                                               slow_peripheral_bridge_m1_qualified_request_sysid_control_slave,
                                               slow_peripheral_bridge_m1_read,
                                               slow_peripheral_bridge_m1_read_data_valid_button_pio_s1,
                                               slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in,
                                               slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in,
                                               slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in,
                                               slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1,
                                               slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
                                               slow_peripheral_bridge_m1_read_data_valid_led_pio_s1,
                                               slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave,
                                               slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1,
                                               slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave,
                                               slow_peripheral_bridge_m1_requests_button_pio_s1,
                                               slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in,
                                               slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in,
                                               slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in,
                                               slow_peripheral_bridge_m1_requests_high_res_timer_s1,
                                               slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave,
                                               slow_peripheral_bridge_m1_requests_led_pio_s1,
                                               slow_peripheral_bridge_m1_requests_performance_counter_control_slave,
                                               slow_peripheral_bridge_m1_requests_sys_clk_timer_s1,
                                               slow_peripheral_bridge_m1_requests_sysid_control_slave,
                                               slow_peripheral_bridge_m1_write,
                                               slow_peripheral_bridge_m1_writedata,
                                               sys_clk_timer_s1_readdata_from_sa,
                                               sysid_control_slave_readdata_from_sa,

                                              // outputs:
                                               slow_peripheral_bridge_m1_address_to_slave,
                                               slow_peripheral_bridge_m1_endofpacket,
                                               slow_peripheral_bridge_m1_latency_counter,
                                               slow_peripheral_bridge_m1_readdata,
                                               slow_peripheral_bridge_m1_readdatavalid,
                                               slow_peripheral_bridge_m1_reset_n,
                                               slow_peripheral_bridge_m1_waitrequest
                                            )
;

  output  [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  output           slow_peripheral_bridge_m1_endofpacket;
  output           slow_peripheral_bridge_m1_latency_counter;
  output  [ 31: 0] slow_peripheral_bridge_m1_readdata;
  output           slow_peripheral_bridge_m1_readdatavalid;
  output           slow_peripheral_bridge_m1_reset_n;
  output           slow_peripheral_bridge_m1_waitrequest;
  input   [ 31: 0] button_pio_s1_readdata_from_sa;
  input            clk;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa;
  input            d1_button_pio_s1_end_xfer;
  input            d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer;
  input            d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer;
  input            d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer;
  input            d1_high_res_timer_s1_end_xfer;
  input            d1_jtag_uart_avalon_jtag_slave_end_xfer;
  input            d1_led_pio_s1_end_xfer;
  input            d1_performance_counter_control_slave_end_xfer;
  input            d1_sys_clk_timer_s1_end_xfer;
  input            d1_sysid_control_slave_end_xfer;
  input   [ 15: 0] high_res_timer_s1_readdata_from_sa;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  input   [ 31: 0] led_pio_s1_readdata_from_sa;
  input   [ 31: 0] performance_counter_control_slave_readdata_from_sa;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address;
  input   [  3: 0] slow_peripheral_bridge_m1_byteenable;
  input            slow_peripheral_bridge_m1_granted_button_pio_s1;
  input            slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  input            slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  input            slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  input            slow_peripheral_bridge_m1_granted_high_res_timer_s1;
  input            slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  input            slow_peripheral_bridge_m1_granted_led_pio_s1;
  input            slow_peripheral_bridge_m1_granted_performance_counter_control_slave;
  input            slow_peripheral_bridge_m1_granted_sys_clk_timer_s1;
  input            slow_peripheral_bridge_m1_granted_sysid_control_slave;
  input            slow_peripheral_bridge_m1_qualified_request_button_pio_s1;
  input            slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  input            slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  input            slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  input            slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1;
  input            slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  input            slow_peripheral_bridge_m1_qualified_request_led_pio_s1;
  input            slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave;
  input            slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1;
  input            slow_peripheral_bridge_m1_qualified_request_sysid_control_slave;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_read_data_valid_button_pio_s1;
  input            slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  input            slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  input            slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  input            slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1;
  input            slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  input            slow_peripheral_bridge_m1_read_data_valid_led_pio_s1;
  input            slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave;
  input            slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1;
  input            slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave;
  input            slow_peripheral_bridge_m1_requests_button_pio_s1;
  input            slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  input            slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  input            slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  input            slow_peripheral_bridge_m1_requests_high_res_timer_s1;
  input            slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  input            slow_peripheral_bridge_m1_requests_led_pio_s1;
  input            slow_peripheral_bridge_m1_requests_performance_counter_control_slave;
  input            slow_peripheral_bridge_m1_requests_sys_clk_timer_s1;
  input            slow_peripheral_bridge_m1_requests_sysid_control_slave;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] slow_peripheral_bridge_m1_writedata;
  input   [ 15: 0] sys_clk_timer_s1_readdata_from_sa;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_slow_peripheral_bridge_m1_latency_counter;
  wire             pre_flush_slow_peripheral_bridge_m1_readdatavalid;
  wire             r_0;
  wire             r_1;
  reg     [  7: 0] slow_peripheral_bridge_m1_address_last_time;
  wire    [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  reg     [  3: 0] slow_peripheral_bridge_m1_byteenable_last_time;
  wire             slow_peripheral_bridge_m1_endofpacket;
  wire             slow_peripheral_bridge_m1_is_granted_some_slave;
  reg              slow_peripheral_bridge_m1_latency_counter;
  reg              slow_peripheral_bridge_m1_read_but_no_slave_selected;
  reg              slow_peripheral_bridge_m1_read_last_time;
  wire    [ 31: 0] slow_peripheral_bridge_m1_readdata;
  wire             slow_peripheral_bridge_m1_readdatavalid;
  wire             slow_peripheral_bridge_m1_reset_n;
  wire             slow_peripheral_bridge_m1_run;
  wire             slow_peripheral_bridge_m1_waitrequest;
  reg              slow_peripheral_bridge_m1_write_last_time;
  reg     [ 31: 0] slow_peripheral_bridge_m1_writedata_last_time;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (slow_peripheral_bridge_m1_qualified_request_button_pio_s1 | ~slow_peripheral_bridge_m1_requests_button_pio_s1) & ((~slow_peripheral_bridge_m1_qualified_request_button_pio_s1 | ~slow_peripheral_bridge_m1_read | (1 & ~d1_button_pio_s1_end_xfer & slow_peripheral_bridge_m1_read))) & ((~slow_peripheral_bridge_m1_qualified_request_button_pio_s1 | ~slow_peripheral_bridge_m1_write | (1 & slow_peripheral_bridge_m1_write))) & 1 & (slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in | ~slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in) & ((~slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in | ~(slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write) | (1 & ~cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)))) & ((~slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in | ~(slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write) | (1 & ~cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)))) & 1 & (slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in | ~slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in) & ((~slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in | ~(slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write) | (1 & ~cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)))) & ((~slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in | ~(slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write) | (1 & ~cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)))) & 1 & (slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in | ~slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in) & ((~slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in | ~(slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write) | (1 & ~cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)))) & ((~slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in | ~(slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write) | (1 & ~cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)))) & 1 & (slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1 | ~slow_peripheral_bridge_m1_requests_high_res_timer_s1) & ((~slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1 | ~slow_peripheral_bridge_m1_read | (1 & ~d1_high_res_timer_s1_end_xfer & slow_peripheral_bridge_m1_read))) & ((~slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1 | ~slow_peripheral_bridge_m1_write | (1 & slow_peripheral_bridge_m1_write)));

  //cascaded wait assignment, which is an e_assign
  assign slow_peripheral_bridge_m1_run = r_0 & r_1;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave) & ((~slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~(slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write) | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)))) & ((~slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~(slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write) | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)))) & 1 & (slow_peripheral_bridge_m1_qualified_request_led_pio_s1 | ~slow_peripheral_bridge_m1_requests_led_pio_s1) & ((~slow_peripheral_bridge_m1_qualified_request_led_pio_s1 | ~slow_peripheral_bridge_m1_read | (1 & ~d1_led_pio_s1_end_xfer & slow_peripheral_bridge_m1_read))) & ((~slow_peripheral_bridge_m1_qualified_request_led_pio_s1 | ~slow_peripheral_bridge_m1_write | (1 & slow_peripheral_bridge_m1_write))) & 1 & (slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave | ~slow_peripheral_bridge_m1_requests_performance_counter_control_slave) & ((~slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave | ~(slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write) | (1 & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)))) & ((~slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave | ~(slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write) | (1 & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)))) & 1 & (slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1 | ~slow_peripheral_bridge_m1_requests_sys_clk_timer_s1) & ((~slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1 | ~slow_peripheral_bridge_m1_read | (1 & ~d1_sys_clk_timer_s1_end_xfer & slow_peripheral_bridge_m1_read))) & ((~slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1 | ~slow_peripheral_bridge_m1_write | (1 & slow_peripheral_bridge_m1_write))) & 1 & (slow_peripheral_bridge_m1_qualified_request_sysid_control_slave | ~slow_peripheral_bridge_m1_requests_sysid_control_slave) & ((~slow_peripheral_bridge_m1_qualified_request_sysid_control_slave | ~slow_peripheral_bridge_m1_read | (1 & ~d1_sysid_control_slave_end_xfer & slow_peripheral_bridge_m1_read))) & ((~slow_peripheral_bridge_m1_qualified_request_sysid_control_slave | ~slow_peripheral_bridge_m1_write | (1 & slow_peripheral_bridge_m1_write)));

  //optimize select-logic by passing only those address bits which matter.
  assign slow_peripheral_bridge_m1_address_to_slave = slow_peripheral_bridge_m1_address[7 : 0];

  //slow_peripheral_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_m1_read_but_no_slave_selected <= 0;
      else 
        slow_peripheral_bridge_m1_read_but_no_slave_selected <= slow_peripheral_bridge_m1_read & slow_peripheral_bridge_m1_run & ~slow_peripheral_bridge_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign slow_peripheral_bridge_m1_is_granted_some_slave = slow_peripheral_bridge_m1_granted_button_pio_s1 |
    slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in |
    slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in |
    slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in |
    slow_peripheral_bridge_m1_granted_high_res_timer_s1 |
    slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave |
    slow_peripheral_bridge_m1_granted_led_pio_s1 |
    slow_peripheral_bridge_m1_granted_performance_counter_control_slave |
    slow_peripheral_bridge_m1_granted_sys_clk_timer_s1 |
    slow_peripheral_bridge_m1_granted_sysid_control_slave;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_slow_peripheral_bridge_m1_readdatavalid = slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign slow_peripheral_bridge_m1_readdatavalid = slow_peripheral_bridge_m1_read_but_no_slave_selected |
    pre_flush_slow_peripheral_bridge_m1_readdatavalid |
    slow_peripheral_bridge_m1_read_data_valid_button_pio_s1 |
    slow_peripheral_bridge_m1_read_but_no_slave_selected |
    pre_flush_slow_peripheral_bridge_m1_readdatavalid |
    slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in |
    slow_peripheral_bridge_m1_read_but_no_slave_selected |
    pre_flush_slow_peripheral_bridge_m1_readdatavalid |
    slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in |
    slow_peripheral_bridge_m1_read_but_no_slave_selected |
    pre_flush_slow_peripheral_bridge_m1_readdatavalid |
    slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in |
    slow_peripheral_bridge_m1_read_but_no_slave_selected |
    pre_flush_slow_peripheral_bridge_m1_readdatavalid |
    slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1 |
    slow_peripheral_bridge_m1_read_but_no_slave_selected |
    pre_flush_slow_peripheral_bridge_m1_readdatavalid |
    slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave |
    slow_peripheral_bridge_m1_read_but_no_slave_selected |
    pre_flush_slow_peripheral_bridge_m1_readdatavalid |
    slow_peripheral_bridge_m1_read_data_valid_led_pio_s1 |
    slow_peripheral_bridge_m1_read_but_no_slave_selected |
    pre_flush_slow_peripheral_bridge_m1_readdatavalid |
    slow_peripheral_bridge_m1_read_but_no_slave_selected |
    pre_flush_slow_peripheral_bridge_m1_readdatavalid |
    slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1 |
    slow_peripheral_bridge_m1_read_but_no_slave_selected |
    pre_flush_slow_peripheral_bridge_m1_readdatavalid |
    slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave;

  //slow_peripheral_bridge/m1 readdata mux, which is an e_mux
  assign slow_peripheral_bridge_m1_readdata = ({32 {~(slow_peripheral_bridge_m1_qualified_request_button_pio_s1 & slow_peripheral_bridge_m1_read)}} | button_pio_s1_readdata_from_sa) &
    ({32 {~(slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in & slow_peripheral_bridge_m1_read)}} | cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa) &
    ({32 {~(slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in & slow_peripheral_bridge_m1_read)}} | cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa) &
    ({32 {~(slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in & slow_peripheral_bridge_m1_read)}} | cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa) &
    ({32 {~(slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1 & slow_peripheral_bridge_m1_read)}} | high_res_timer_s1_readdata_from_sa) &
    ({32 {~(slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave & slow_peripheral_bridge_m1_read)}} | jtag_uart_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~(slow_peripheral_bridge_m1_qualified_request_led_pio_s1 & slow_peripheral_bridge_m1_read)}} | led_pio_s1_readdata_from_sa) &
    ({32 {~slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave}} | performance_counter_control_slave_readdata_from_sa) &
    ({32 {~(slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1 & slow_peripheral_bridge_m1_read)}} | sys_clk_timer_s1_readdata_from_sa) &
    ({32 {~(slow_peripheral_bridge_m1_qualified_request_sysid_control_slave & slow_peripheral_bridge_m1_read)}} | sysid_control_slave_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign slow_peripheral_bridge_m1_waitrequest = ~slow_peripheral_bridge_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_m1_latency_counter <= 0;
      else 
        slow_peripheral_bridge_m1_latency_counter <= p1_slow_peripheral_bridge_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_slow_peripheral_bridge_m1_latency_counter = ((slow_peripheral_bridge_m1_run & slow_peripheral_bridge_m1_read))? latency_load_value :
    (slow_peripheral_bridge_m1_latency_counter)? slow_peripheral_bridge_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {slow_peripheral_bridge_m1_requests_performance_counter_control_slave}} & 1;

  //slow_peripheral_bridge_m1_reset_n assignment, which is an e_assign
  assign slow_peripheral_bridge_m1_reset_n = reset_n;

  //mux slow_peripheral_bridge_m1_endofpacket, which is an e_mux
  assign slow_peripheral_bridge_m1_endofpacket = (slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in)? cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa :
    (slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in)? cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa :
    cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //slow_peripheral_bridge_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_m1_address_last_time <= 0;
      else 
        slow_peripheral_bridge_m1_address_last_time <= slow_peripheral_bridge_m1_address;
    end


  //slow_peripheral_bridge/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= slow_peripheral_bridge_m1_waitrequest & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write);
    end


  //slow_peripheral_bridge_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (slow_peripheral_bridge_m1_address != slow_peripheral_bridge_m1_address_last_time))
        begin
          $write("%0d ns: slow_peripheral_bridge_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //slow_peripheral_bridge_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_m1_byteenable_last_time <= 0;
      else 
        slow_peripheral_bridge_m1_byteenable_last_time <= slow_peripheral_bridge_m1_byteenable;
    end


  //slow_peripheral_bridge_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (slow_peripheral_bridge_m1_byteenable != slow_peripheral_bridge_m1_byteenable_last_time))
        begin
          $write("%0d ns: slow_peripheral_bridge_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //slow_peripheral_bridge_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_m1_read_last_time <= 0;
      else 
        slow_peripheral_bridge_m1_read_last_time <= slow_peripheral_bridge_m1_read;
    end


  //slow_peripheral_bridge_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (slow_peripheral_bridge_m1_read != slow_peripheral_bridge_m1_read_last_time))
        begin
          $write("%0d ns: slow_peripheral_bridge_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //slow_peripheral_bridge_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_m1_write_last_time <= 0;
      else 
        slow_peripheral_bridge_m1_write_last_time <= slow_peripheral_bridge_m1_write;
    end


  //slow_peripheral_bridge_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (slow_peripheral_bridge_m1_write != slow_peripheral_bridge_m1_write_last_time))
        begin
          $write("%0d ns: slow_peripheral_bridge_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //slow_peripheral_bridge_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          slow_peripheral_bridge_m1_writedata_last_time <= 0;
      else 
        slow_peripheral_bridge_m1_writedata_last_time <= slow_peripheral_bridge_m1_writedata;
    end


  //slow_peripheral_bridge_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (slow_peripheral_bridge_m1_writedata != slow_peripheral_bridge_m1_writedata_last_time) & slow_peripheral_bridge_m1_write)
        begin
          $write("%0d ns: slow_peripheral_bridge_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module slow_peripheral_bridge_bridge_arbitrator 
;



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sys_clk_timer_s1_arbitrator (
                                     // inputs:
                                      clk,
                                      reset_n,
                                      slow_peripheral_bridge_m1_address_to_slave,
                                      slow_peripheral_bridge_m1_latency_counter,
                                      slow_peripheral_bridge_m1_nativeaddress,
                                      slow_peripheral_bridge_m1_read,
                                      slow_peripheral_bridge_m1_write,
                                      slow_peripheral_bridge_m1_writedata,
                                      sys_clk_timer_s1_irq,
                                      sys_clk_timer_s1_readdata,

                                     // outputs:
                                      d1_sys_clk_timer_s1_end_xfer,
                                      slow_peripheral_bridge_m1_granted_sys_clk_timer_s1,
                                      slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1,
                                      slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1,
                                      slow_peripheral_bridge_m1_requests_sys_clk_timer_s1,
                                      sys_clk_timer_s1_address,
                                      sys_clk_timer_s1_chipselect,
                                      sys_clk_timer_s1_irq_from_sa,
                                      sys_clk_timer_s1_readdata_from_sa,
                                      sys_clk_timer_s1_reset_n,
                                      sys_clk_timer_s1_write_n,
                                      sys_clk_timer_s1_writedata
                                   )
;

  output           d1_sys_clk_timer_s1_end_xfer;
  output           slow_peripheral_bridge_m1_granted_sys_clk_timer_s1;
  output           slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1;
  output           slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1;
  output           slow_peripheral_bridge_m1_requests_sys_clk_timer_s1;
  output  [  2: 0] sys_clk_timer_s1_address;
  output           sys_clk_timer_s1_chipselect;
  output           sys_clk_timer_s1_irq_from_sa;
  output  [ 15: 0] sys_clk_timer_s1_readdata_from_sa;
  output           sys_clk_timer_s1_reset_n;
  output           sys_clk_timer_s1_write_n;
  output  [ 15: 0] sys_clk_timer_s1_writedata;
  input            clk;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  input            slow_peripheral_bridge_m1_latency_counter;
  input   [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] slow_peripheral_bridge_m1_writedata;
  input            sys_clk_timer_s1_irq;
  input   [ 15: 0] sys_clk_timer_s1_readdata;

  reg              d1_reasons_to_wait;
  reg              d1_sys_clk_timer_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sys_clk_timer_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             slow_peripheral_bridge_m1_arbiterlock;
  wire             slow_peripheral_bridge_m1_arbiterlock2;
  wire             slow_peripheral_bridge_m1_continuerequest;
  wire             slow_peripheral_bridge_m1_granted_sys_clk_timer_s1;
  wire             slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1;
  wire             slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1;
  wire             slow_peripheral_bridge_m1_requests_sys_clk_timer_s1;
  wire             slow_peripheral_bridge_m1_saved_grant_sys_clk_timer_s1;
  wire    [  2: 0] sys_clk_timer_s1_address;
  wire             sys_clk_timer_s1_allgrants;
  wire             sys_clk_timer_s1_allow_new_arb_cycle;
  wire             sys_clk_timer_s1_any_bursting_master_saved_grant;
  wire             sys_clk_timer_s1_any_continuerequest;
  wire             sys_clk_timer_s1_arb_counter_enable;
  reg              sys_clk_timer_s1_arb_share_counter;
  wire             sys_clk_timer_s1_arb_share_counter_next_value;
  wire             sys_clk_timer_s1_arb_share_set_values;
  wire             sys_clk_timer_s1_beginbursttransfer_internal;
  wire             sys_clk_timer_s1_begins_xfer;
  wire             sys_clk_timer_s1_chipselect;
  wire             sys_clk_timer_s1_end_xfer;
  wire             sys_clk_timer_s1_firsttransfer;
  wire             sys_clk_timer_s1_grant_vector;
  wire             sys_clk_timer_s1_in_a_read_cycle;
  wire             sys_clk_timer_s1_in_a_write_cycle;
  wire             sys_clk_timer_s1_irq_from_sa;
  wire             sys_clk_timer_s1_master_qreq_vector;
  wire             sys_clk_timer_s1_non_bursting_master_requests;
  wire    [ 15: 0] sys_clk_timer_s1_readdata_from_sa;
  reg              sys_clk_timer_s1_reg_firsttransfer;
  wire             sys_clk_timer_s1_reset_n;
  reg              sys_clk_timer_s1_slavearbiterlockenable;
  wire             sys_clk_timer_s1_slavearbiterlockenable2;
  wire             sys_clk_timer_s1_unreg_firsttransfer;
  wire             sys_clk_timer_s1_waits_for_read;
  wire             sys_clk_timer_s1_waits_for_write;
  wire             sys_clk_timer_s1_write_n;
  wire    [ 15: 0] sys_clk_timer_s1_writedata;
  wire             wait_for_sys_clk_timer_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sys_clk_timer_s1_end_xfer;
    end


  assign sys_clk_timer_s1_begins_xfer = ~d1_reasons_to_wait & ((slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1));
  //assign sys_clk_timer_s1_readdata_from_sa = sys_clk_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sys_clk_timer_s1_readdata_from_sa = sys_clk_timer_s1_readdata;

  assign slow_peripheral_bridge_m1_requests_sys_clk_timer_s1 = ({slow_peripheral_bridge_m1_address_to_slave[7 : 5] , 5'b0} == 8'ha0) & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write);
  //sys_clk_timer_s1_arb_share_counter set values, which is an e_mux
  assign sys_clk_timer_s1_arb_share_set_values = 1;

  //sys_clk_timer_s1_non_bursting_master_requests mux, which is an e_mux
  assign sys_clk_timer_s1_non_bursting_master_requests = slow_peripheral_bridge_m1_requests_sys_clk_timer_s1;

  //sys_clk_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign sys_clk_timer_s1_any_bursting_master_saved_grant = 0;

  //sys_clk_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign sys_clk_timer_s1_arb_share_counter_next_value = sys_clk_timer_s1_firsttransfer ? (sys_clk_timer_s1_arb_share_set_values - 1) : |sys_clk_timer_s1_arb_share_counter ? (sys_clk_timer_s1_arb_share_counter - 1) : 0;

  //sys_clk_timer_s1_allgrants all slave grants, which is an e_mux
  assign sys_clk_timer_s1_allgrants = |sys_clk_timer_s1_grant_vector;

  //sys_clk_timer_s1_end_xfer assignment, which is an e_assign
  assign sys_clk_timer_s1_end_xfer = ~(sys_clk_timer_s1_waits_for_read | sys_clk_timer_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_sys_clk_timer_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sys_clk_timer_s1 = sys_clk_timer_s1_end_xfer & (~sys_clk_timer_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sys_clk_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign sys_clk_timer_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_sys_clk_timer_s1 & sys_clk_timer_s1_allgrants) | (end_xfer_arb_share_counter_term_sys_clk_timer_s1 & ~sys_clk_timer_s1_non_bursting_master_requests);

  //sys_clk_timer_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_clk_timer_s1_arb_share_counter <= 0;
      else if (sys_clk_timer_s1_arb_counter_enable)
          sys_clk_timer_s1_arb_share_counter <= sys_clk_timer_s1_arb_share_counter_next_value;
    end


  //sys_clk_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_clk_timer_s1_slavearbiterlockenable <= 0;
      else if ((|sys_clk_timer_s1_master_qreq_vector & end_xfer_arb_share_counter_term_sys_clk_timer_s1) | (end_xfer_arb_share_counter_term_sys_clk_timer_s1 & ~sys_clk_timer_s1_non_bursting_master_requests))
          sys_clk_timer_s1_slavearbiterlockenable <= |sys_clk_timer_s1_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge/m1 sys_clk_timer/s1 arbiterlock, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock = sys_clk_timer_s1_slavearbiterlockenable & slow_peripheral_bridge_m1_continuerequest;

  //sys_clk_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sys_clk_timer_s1_slavearbiterlockenable2 = |sys_clk_timer_s1_arb_share_counter_next_value;

  //slow_peripheral_bridge/m1 sys_clk_timer/s1 arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock2 = sys_clk_timer_s1_slavearbiterlockenable2 & slow_peripheral_bridge_m1_continuerequest;

  //sys_clk_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sys_clk_timer_s1_any_continuerequest = 1;

  //slow_peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  assign slow_peripheral_bridge_m1_continuerequest = 1;

  assign slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1 = slow_peripheral_bridge_m1_requests_sys_clk_timer_s1 & ~((slow_peripheral_bridge_m1_read & ((slow_peripheral_bridge_m1_latency_counter != 0))));
  //local readdatavalid slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1 = slow_peripheral_bridge_m1_granted_sys_clk_timer_s1 & slow_peripheral_bridge_m1_read & ~sys_clk_timer_s1_waits_for_read;

  //sys_clk_timer_s1_writedata mux, which is an e_mux
  assign sys_clk_timer_s1_writedata = slow_peripheral_bridge_m1_writedata;

  //master is always granted when requested
  assign slow_peripheral_bridge_m1_granted_sys_clk_timer_s1 = slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1;

  //slow_peripheral_bridge/m1 saved-grant sys_clk_timer/s1, which is an e_assign
  assign slow_peripheral_bridge_m1_saved_grant_sys_clk_timer_s1 = slow_peripheral_bridge_m1_requests_sys_clk_timer_s1;

  //allow new arb cycle for sys_clk_timer/s1, which is an e_assign
  assign sys_clk_timer_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sys_clk_timer_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sys_clk_timer_s1_master_qreq_vector = 1;

  //sys_clk_timer_s1_reset_n assignment, which is an e_assign
  assign sys_clk_timer_s1_reset_n = reset_n;

  assign sys_clk_timer_s1_chipselect = slow_peripheral_bridge_m1_granted_sys_clk_timer_s1;
  //sys_clk_timer_s1_firsttransfer first transaction, which is an e_assign
  assign sys_clk_timer_s1_firsttransfer = sys_clk_timer_s1_begins_xfer ? sys_clk_timer_s1_unreg_firsttransfer : sys_clk_timer_s1_reg_firsttransfer;

  //sys_clk_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign sys_clk_timer_s1_unreg_firsttransfer = ~(sys_clk_timer_s1_slavearbiterlockenable & sys_clk_timer_s1_any_continuerequest);

  //sys_clk_timer_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sys_clk_timer_s1_reg_firsttransfer <= 1'b1;
      else if (sys_clk_timer_s1_begins_xfer)
          sys_clk_timer_s1_reg_firsttransfer <= sys_clk_timer_s1_unreg_firsttransfer;
    end


  //sys_clk_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sys_clk_timer_s1_beginbursttransfer_internal = sys_clk_timer_s1_begins_xfer;

  //~sys_clk_timer_s1_write_n assignment, which is an e_mux
  assign sys_clk_timer_s1_write_n = ~(slow_peripheral_bridge_m1_granted_sys_clk_timer_s1 & slow_peripheral_bridge_m1_write);

  //sys_clk_timer_s1_address mux, which is an e_mux
  assign sys_clk_timer_s1_address = slow_peripheral_bridge_m1_nativeaddress;

  //d1_sys_clk_timer_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sys_clk_timer_s1_end_xfer <= 1;
      else 
        d1_sys_clk_timer_s1_end_xfer <= sys_clk_timer_s1_end_xfer;
    end


  //sys_clk_timer_s1_waits_for_read in a cycle, which is an e_mux
  assign sys_clk_timer_s1_waits_for_read = sys_clk_timer_s1_in_a_read_cycle & sys_clk_timer_s1_begins_xfer;

  //sys_clk_timer_s1_in_a_read_cycle assignment, which is an e_assign
  assign sys_clk_timer_s1_in_a_read_cycle = slow_peripheral_bridge_m1_granted_sys_clk_timer_s1 & slow_peripheral_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sys_clk_timer_s1_in_a_read_cycle;

  //sys_clk_timer_s1_waits_for_write in a cycle, which is an e_mux
  assign sys_clk_timer_s1_waits_for_write = sys_clk_timer_s1_in_a_write_cycle & 0;

  //sys_clk_timer_s1_in_a_write_cycle assignment, which is an e_assign
  assign sys_clk_timer_s1_in_a_write_cycle = slow_peripheral_bridge_m1_granted_sys_clk_timer_s1 & slow_peripheral_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sys_clk_timer_s1_in_a_write_cycle;

  assign wait_for_sys_clk_timer_s1_counter = 0;
  //assign sys_clk_timer_s1_irq_from_sa = sys_clk_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sys_clk_timer_s1_irq_from_sa = sys_clk_timer_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sys_clk_timer/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sysid_control_slave_arbitrator (
                                        // inputs:
                                         clk,
                                         reset_n,
                                         slow_peripheral_bridge_m1_address_to_slave,
                                         slow_peripheral_bridge_m1_latency_counter,
                                         slow_peripheral_bridge_m1_nativeaddress,
                                         slow_peripheral_bridge_m1_read,
                                         slow_peripheral_bridge_m1_write,
                                         sysid_control_slave_readdata,

                                        // outputs:
                                         d1_sysid_control_slave_end_xfer,
                                         slow_peripheral_bridge_m1_granted_sysid_control_slave,
                                         slow_peripheral_bridge_m1_qualified_request_sysid_control_slave,
                                         slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave,
                                         slow_peripheral_bridge_m1_requests_sysid_control_slave,
                                         sysid_control_slave_address,
                                         sysid_control_slave_readdata_from_sa,
                                         sysid_control_slave_reset_n
                                      )
;

  output           d1_sysid_control_slave_end_xfer;
  output           slow_peripheral_bridge_m1_granted_sysid_control_slave;
  output           slow_peripheral_bridge_m1_qualified_request_sysid_control_slave;
  output           slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave;
  output           slow_peripheral_bridge_m1_requests_sysid_control_slave;
  output           sysid_control_slave_address;
  output  [ 31: 0] sysid_control_slave_readdata_from_sa;
  output           sysid_control_slave_reset_n;
  input            clk;
  input            reset_n;
  input   [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  input            slow_peripheral_bridge_m1_latency_counter;
  input   [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  input            slow_peripheral_bridge_m1_read;
  input            slow_peripheral_bridge_m1_write;
  input   [ 31: 0] sysid_control_slave_readdata;

  reg              d1_reasons_to_wait;
  reg              d1_sysid_control_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sysid_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             slow_peripheral_bridge_m1_arbiterlock;
  wire             slow_peripheral_bridge_m1_arbiterlock2;
  wire             slow_peripheral_bridge_m1_continuerequest;
  wire             slow_peripheral_bridge_m1_granted_sysid_control_slave;
  wire             slow_peripheral_bridge_m1_qualified_request_sysid_control_slave;
  wire             slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave;
  wire             slow_peripheral_bridge_m1_requests_sysid_control_slave;
  wire             slow_peripheral_bridge_m1_saved_grant_sysid_control_slave;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_allgrants;
  wire             sysid_control_slave_allow_new_arb_cycle;
  wire             sysid_control_slave_any_bursting_master_saved_grant;
  wire             sysid_control_slave_any_continuerequest;
  wire             sysid_control_slave_arb_counter_enable;
  reg              sysid_control_slave_arb_share_counter;
  wire             sysid_control_slave_arb_share_counter_next_value;
  wire             sysid_control_slave_arb_share_set_values;
  wire             sysid_control_slave_beginbursttransfer_internal;
  wire             sysid_control_slave_begins_xfer;
  wire             sysid_control_slave_end_xfer;
  wire             sysid_control_slave_firsttransfer;
  wire             sysid_control_slave_grant_vector;
  wire             sysid_control_slave_in_a_read_cycle;
  wire             sysid_control_slave_in_a_write_cycle;
  wire             sysid_control_slave_master_qreq_vector;
  wire             sysid_control_slave_non_bursting_master_requests;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  reg              sysid_control_slave_reg_firsttransfer;
  wire             sysid_control_slave_reset_n;
  reg              sysid_control_slave_slavearbiterlockenable;
  wire             sysid_control_slave_slavearbiterlockenable2;
  wire             sysid_control_slave_unreg_firsttransfer;
  wire             sysid_control_slave_waits_for_read;
  wire             sysid_control_slave_waits_for_write;
  wire             wait_for_sysid_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sysid_control_slave_end_xfer;
    end


  assign sysid_control_slave_begins_xfer = ~d1_reasons_to_wait & ((slow_peripheral_bridge_m1_qualified_request_sysid_control_slave));
  //assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata;

  assign slow_peripheral_bridge_m1_requests_sysid_control_slave = (({slow_peripheral_bridge_m1_address_to_slave[7 : 3] , 3'b0} == 8'he8) & (slow_peripheral_bridge_m1_read | slow_peripheral_bridge_m1_write)) & slow_peripheral_bridge_m1_read;
  //sysid_control_slave_arb_share_counter set values, which is an e_mux
  assign sysid_control_slave_arb_share_set_values = 1;

  //sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign sysid_control_slave_non_bursting_master_requests = slow_peripheral_bridge_m1_requests_sysid_control_slave;

  //sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign sysid_control_slave_any_bursting_master_saved_grant = 0;

  //sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign sysid_control_slave_arb_share_counter_next_value = sysid_control_slave_firsttransfer ? (sysid_control_slave_arb_share_set_values - 1) : |sysid_control_slave_arb_share_counter ? (sysid_control_slave_arb_share_counter - 1) : 0;

  //sysid_control_slave_allgrants all slave grants, which is an e_mux
  assign sysid_control_slave_allgrants = |sysid_control_slave_grant_vector;

  //sysid_control_slave_end_xfer assignment, which is an e_assign
  assign sysid_control_slave_end_xfer = ~(sysid_control_slave_waits_for_read | sysid_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sysid_control_slave = sysid_control_slave_end_xfer & (~sysid_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign sysid_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_sysid_control_slave & sysid_control_slave_allgrants) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests);

  //sysid_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_arb_share_counter <= 0;
      else if (sysid_control_slave_arb_counter_enable)
          sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
    end


  //sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_slavearbiterlockenable <= 0;
      else if ((|sysid_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_sysid_control_slave) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests))
          sysid_control_slave_slavearbiterlockenable <= |sysid_control_slave_arb_share_counter_next_value;
    end


  //slow_peripheral_bridge/m1 sysid/control_slave arbiterlock, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock = sysid_control_slave_slavearbiterlockenable & slow_peripheral_bridge_m1_continuerequest;

  //sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sysid_control_slave_slavearbiterlockenable2 = |sysid_control_slave_arb_share_counter_next_value;

  //slow_peripheral_bridge/m1 sysid/control_slave arbiterlock2, which is an e_assign
  assign slow_peripheral_bridge_m1_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & slow_peripheral_bridge_m1_continuerequest;

  //sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sysid_control_slave_any_continuerequest = 1;

  //slow_peripheral_bridge_m1_continuerequest continued request, which is an e_assign
  assign slow_peripheral_bridge_m1_continuerequest = 1;

  assign slow_peripheral_bridge_m1_qualified_request_sysid_control_slave = slow_peripheral_bridge_m1_requests_sysid_control_slave & ~((slow_peripheral_bridge_m1_read & ((slow_peripheral_bridge_m1_latency_counter != 0))));
  //local readdatavalid slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave, which is an e_mux
  assign slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave = slow_peripheral_bridge_m1_granted_sysid_control_slave & slow_peripheral_bridge_m1_read & ~sysid_control_slave_waits_for_read;

  //master is always granted when requested
  assign slow_peripheral_bridge_m1_granted_sysid_control_slave = slow_peripheral_bridge_m1_qualified_request_sysid_control_slave;

  //slow_peripheral_bridge/m1 saved-grant sysid/control_slave, which is an e_assign
  assign slow_peripheral_bridge_m1_saved_grant_sysid_control_slave = slow_peripheral_bridge_m1_requests_sysid_control_slave;

  //allow new arb cycle for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sysid_control_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sysid_control_slave_master_qreq_vector = 1;

  //sysid_control_slave_reset_n assignment, which is an e_assign
  assign sysid_control_slave_reset_n = reset_n;

  //sysid_control_slave_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_firsttransfer = sysid_control_slave_begins_xfer ? sysid_control_slave_unreg_firsttransfer : sysid_control_slave_reg_firsttransfer;

  //sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_unreg_firsttransfer = ~(sysid_control_slave_slavearbiterlockenable & sysid_control_slave_any_continuerequest);

  //sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_reg_firsttransfer <= 1'b1;
      else if (sysid_control_slave_begins_xfer)
          sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
    end


  //sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sysid_control_slave_beginbursttransfer_internal = sysid_control_slave_begins_xfer;

  //sysid_control_slave_address mux, which is an e_mux
  assign sysid_control_slave_address = slow_peripheral_bridge_m1_nativeaddress;

  //d1_sysid_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sysid_control_slave_end_xfer <= 1;
      else 
        d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end


  //sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_read = sysid_control_slave_in_a_read_cycle & sysid_control_slave_begins_xfer;

  //sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_read_cycle = slow_peripheral_bridge_m1_granted_sysid_control_slave & slow_peripheral_bridge_m1_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sysid_control_slave_in_a_read_cycle;

  //sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_write = sysid_control_slave_in_a_write_cycle & 0;

  //sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_write_cycle = slow_peripheral_bridge_m1_granted_sysid_control_slave & slow_peripheral_bridge_m1_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sysid_control_slave_in_a_write_cycle;

  assign wait_for_sysid_control_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sysid/control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_mac_control_port_arbitrator (
                                         // inputs:
                                          clk,
                                          cpu_data_master_address_to_slave,
                                          cpu_data_master_latency_counter,
                                          cpu_data_master_read,
                                          cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register,
                                          cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register,
                                          cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register,
                                          cpu_data_master_write,
                                          cpu_data_master_writedata,
                                          reset_n,
                                          tse_mac_control_port_readdata,
                                          tse_mac_control_port_waitrequest,

                                         // outputs:
                                          cpu_data_master_granted_tse_mac_control_port,
                                          cpu_data_master_qualified_request_tse_mac_control_port,
                                          cpu_data_master_read_data_valid_tse_mac_control_port,
                                          cpu_data_master_requests_tse_mac_control_port,
                                          d1_tse_mac_control_port_end_xfer,
                                          tse_mac_control_port_address,
                                          tse_mac_control_port_read,
                                          tse_mac_control_port_readdata_from_sa,
                                          tse_mac_control_port_reset,
                                          tse_mac_control_port_waitrequest_from_sa,
                                          tse_mac_control_port_write,
                                          tse_mac_control_port_writedata
                                       )
;

  output           cpu_data_master_granted_tse_mac_control_port;
  output           cpu_data_master_qualified_request_tse_mac_control_port;
  output           cpu_data_master_read_data_valid_tse_mac_control_port;
  output           cpu_data_master_requests_tse_mac_control_port;
  output           d1_tse_mac_control_port_end_xfer;
  output  [  7: 0] tse_mac_control_port_address;
  output           tse_mac_control_port_read;
  output  [ 31: 0] tse_mac_control_port_readdata_from_sa;
  output           tse_mac_control_port_reset;
  output           tse_mac_control_port_waitrequest_from_sa;
  output           tse_mac_control_port_write;
  output  [ 31: 0] tse_mac_control_port_writedata;
  input            clk;
  input   [ 28: 0] cpu_data_master_address_to_slave;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  input            cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] tse_mac_control_port_readdata;
  input            tse_mac_control_port_waitrequest;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_tse_mac_control_port;
  wire             cpu_data_master_qualified_request_tse_mac_control_port;
  wire             cpu_data_master_read_data_valid_tse_mac_control_port;
  wire             cpu_data_master_requests_tse_mac_control_port;
  wire             cpu_data_master_saved_grant_tse_mac_control_port;
  reg              d1_reasons_to_wait;
  reg              d1_tse_mac_control_port_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tse_mac_control_port;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 28: 0] shifted_address_to_tse_mac_control_port_from_cpu_data_master;
  wire    [  7: 0] tse_mac_control_port_address;
  wire             tse_mac_control_port_allgrants;
  wire             tse_mac_control_port_allow_new_arb_cycle;
  wire             tse_mac_control_port_any_bursting_master_saved_grant;
  wire             tse_mac_control_port_any_continuerequest;
  wire             tse_mac_control_port_arb_counter_enable;
  reg              tse_mac_control_port_arb_share_counter;
  wire             tse_mac_control_port_arb_share_counter_next_value;
  wire             tse_mac_control_port_arb_share_set_values;
  wire             tse_mac_control_port_beginbursttransfer_internal;
  wire             tse_mac_control_port_begins_xfer;
  wire             tse_mac_control_port_end_xfer;
  wire             tse_mac_control_port_firsttransfer;
  wire             tse_mac_control_port_grant_vector;
  wire             tse_mac_control_port_in_a_read_cycle;
  wire             tse_mac_control_port_in_a_write_cycle;
  wire             tse_mac_control_port_master_qreq_vector;
  wire             tse_mac_control_port_non_bursting_master_requests;
  wire             tse_mac_control_port_read;
  wire    [ 31: 0] tse_mac_control_port_readdata_from_sa;
  reg              tse_mac_control_port_reg_firsttransfer;
  wire             tse_mac_control_port_reset;
  reg              tse_mac_control_port_slavearbiterlockenable;
  wire             tse_mac_control_port_slavearbiterlockenable2;
  wire             tse_mac_control_port_unreg_firsttransfer;
  wire             tse_mac_control_port_waitrequest_from_sa;
  wire             tse_mac_control_port_waits_for_read;
  wire             tse_mac_control_port_waits_for_write;
  wire             tse_mac_control_port_write;
  wire    [ 31: 0] tse_mac_control_port_writedata;
  wire             wait_for_tse_mac_control_port_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tse_mac_control_port_end_xfer;
    end


  assign tse_mac_control_port_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_tse_mac_control_port));
  //assign tse_mac_control_port_readdata_from_sa = tse_mac_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_mac_control_port_readdata_from_sa = tse_mac_control_port_readdata;

  assign cpu_data_master_requests_tse_mac_control_port = ({cpu_data_master_address_to_slave[28 : 10] , 10'b0} == 29'h1002800) & (cpu_data_master_read | cpu_data_master_write);
  //assign tse_mac_control_port_waitrequest_from_sa = tse_mac_control_port_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_mac_control_port_waitrequest_from_sa = tse_mac_control_port_waitrequest;

  //tse_mac_control_port_arb_share_counter set values, which is an e_mux
  assign tse_mac_control_port_arb_share_set_values = 1;

  //tse_mac_control_port_non_bursting_master_requests mux, which is an e_mux
  assign tse_mac_control_port_non_bursting_master_requests = cpu_data_master_requests_tse_mac_control_port;

  //tse_mac_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  assign tse_mac_control_port_any_bursting_master_saved_grant = 0;

  //tse_mac_control_port_arb_share_counter_next_value assignment, which is an e_assign
  assign tse_mac_control_port_arb_share_counter_next_value = tse_mac_control_port_firsttransfer ? (tse_mac_control_port_arb_share_set_values - 1) : |tse_mac_control_port_arb_share_counter ? (tse_mac_control_port_arb_share_counter - 1) : 0;

  //tse_mac_control_port_allgrants all slave grants, which is an e_mux
  assign tse_mac_control_port_allgrants = |tse_mac_control_port_grant_vector;

  //tse_mac_control_port_end_xfer assignment, which is an e_assign
  assign tse_mac_control_port_end_xfer = ~(tse_mac_control_port_waits_for_read | tse_mac_control_port_waits_for_write);

  //end_xfer_arb_share_counter_term_tse_mac_control_port arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tse_mac_control_port = tse_mac_control_port_end_xfer & (~tse_mac_control_port_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tse_mac_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  assign tse_mac_control_port_arb_counter_enable = (end_xfer_arb_share_counter_term_tse_mac_control_port & tse_mac_control_port_allgrants) | (end_xfer_arb_share_counter_term_tse_mac_control_port & ~tse_mac_control_port_non_bursting_master_requests);

  //tse_mac_control_port_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_mac_control_port_arb_share_counter <= 0;
      else if (tse_mac_control_port_arb_counter_enable)
          tse_mac_control_port_arb_share_counter <= tse_mac_control_port_arb_share_counter_next_value;
    end


  //tse_mac_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_mac_control_port_slavearbiterlockenable <= 0;
      else if ((|tse_mac_control_port_master_qreq_vector & end_xfer_arb_share_counter_term_tse_mac_control_port) | (end_xfer_arb_share_counter_term_tse_mac_control_port & ~tse_mac_control_port_non_bursting_master_requests))
          tse_mac_control_port_slavearbiterlockenable <= |tse_mac_control_port_arb_share_counter_next_value;
    end


  //cpu/data_master tse_mac/control_port arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = tse_mac_control_port_slavearbiterlockenable & cpu_data_master_continuerequest;

  //tse_mac_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tse_mac_control_port_slavearbiterlockenable2 = |tse_mac_control_port_arb_share_counter_next_value;

  //cpu/data_master tse_mac/control_port arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = tse_mac_control_port_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //tse_mac_control_port_any_continuerequest at least one master continues requesting, which is an e_assign
  assign tse_mac_control_port_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_tse_mac_control_port = cpu_data_master_requests_tse_mac_control_port & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (|cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register) | (|cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register))));
  //local readdatavalid cpu_data_master_read_data_valid_tse_mac_control_port, which is an e_mux
  assign cpu_data_master_read_data_valid_tse_mac_control_port = cpu_data_master_granted_tse_mac_control_port & cpu_data_master_read & ~tse_mac_control_port_waits_for_read;

  //tse_mac_control_port_writedata mux, which is an e_mux
  assign tse_mac_control_port_writedata = cpu_data_master_writedata;

  //master is always granted when requested
  assign cpu_data_master_granted_tse_mac_control_port = cpu_data_master_qualified_request_tse_mac_control_port;

  //cpu/data_master saved-grant tse_mac/control_port, which is an e_assign
  assign cpu_data_master_saved_grant_tse_mac_control_port = cpu_data_master_requests_tse_mac_control_port;

  //allow new arb cycle for tse_mac/control_port, which is an e_assign
  assign tse_mac_control_port_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign tse_mac_control_port_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign tse_mac_control_port_master_qreq_vector = 1;

  //~tse_mac_control_port_reset assignment, which is an e_assign
  assign tse_mac_control_port_reset = ~reset_n;

  //tse_mac_control_port_firsttransfer first transaction, which is an e_assign
  assign tse_mac_control_port_firsttransfer = tse_mac_control_port_begins_xfer ? tse_mac_control_port_unreg_firsttransfer : tse_mac_control_port_reg_firsttransfer;

  //tse_mac_control_port_unreg_firsttransfer first transaction, which is an e_assign
  assign tse_mac_control_port_unreg_firsttransfer = ~(tse_mac_control_port_slavearbiterlockenable & tse_mac_control_port_any_continuerequest);

  //tse_mac_control_port_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_mac_control_port_reg_firsttransfer <= 1'b1;
      else if (tse_mac_control_port_begins_xfer)
          tse_mac_control_port_reg_firsttransfer <= tse_mac_control_port_unreg_firsttransfer;
    end


  //tse_mac_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tse_mac_control_port_beginbursttransfer_internal = tse_mac_control_port_begins_xfer;

  //tse_mac_control_port_read assignment, which is an e_mux
  assign tse_mac_control_port_read = cpu_data_master_granted_tse_mac_control_port & cpu_data_master_read;

  //tse_mac_control_port_write assignment, which is an e_mux
  assign tse_mac_control_port_write = cpu_data_master_granted_tse_mac_control_port & cpu_data_master_write;

  assign shifted_address_to_tse_mac_control_port_from_cpu_data_master = cpu_data_master_address_to_slave;
  //tse_mac_control_port_address mux, which is an e_mux
  assign tse_mac_control_port_address = shifted_address_to_tse_mac_control_port_from_cpu_data_master >> 2;

  //d1_tse_mac_control_port_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tse_mac_control_port_end_xfer <= 1;
      else 
        d1_tse_mac_control_port_end_xfer <= tse_mac_control_port_end_xfer;
    end


  //tse_mac_control_port_waits_for_read in a cycle, which is an e_mux
  assign tse_mac_control_port_waits_for_read = tse_mac_control_port_in_a_read_cycle & tse_mac_control_port_waitrequest_from_sa;

  //tse_mac_control_port_in_a_read_cycle assignment, which is an e_assign
  assign tse_mac_control_port_in_a_read_cycle = cpu_data_master_granted_tse_mac_control_port & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tse_mac_control_port_in_a_read_cycle;

  //tse_mac_control_port_waits_for_write in a cycle, which is an e_mux
  assign tse_mac_control_port_waits_for_write = tse_mac_control_port_in_a_write_cycle & tse_mac_control_port_waitrequest_from_sa;

  //tse_mac_control_port_in_a_write_cycle assignment, which is an e_assign
  assign tse_mac_control_port_in_a_write_cycle = cpu_data_master_granted_tse_mac_control_port & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tse_mac_control_port_in_a_write_cycle;

  assign wait_for_tse_mac_control_port_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tse_mac/control_port enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_mac_transmit_arbitrator (
                                     // inputs:
                                      clk,
                                      reset_n,
                                      sgdma_tx_out_data,
                                      sgdma_tx_out_empty,
                                      sgdma_tx_out_endofpacket,
                                      sgdma_tx_out_error,
                                      sgdma_tx_out_startofpacket,
                                      sgdma_tx_out_valid,
                                      tse_mac_transmit_ready,

                                     // outputs:
                                      tse_mac_transmit_data,
                                      tse_mac_transmit_empty,
                                      tse_mac_transmit_endofpacket,
                                      tse_mac_transmit_error,
                                      tse_mac_transmit_ready_from_sa,
                                      tse_mac_transmit_startofpacket,
                                      tse_mac_transmit_valid
                                   )
;

  output  [ 31: 0] tse_mac_transmit_data;
  output  [  1: 0] tse_mac_transmit_empty;
  output           tse_mac_transmit_endofpacket;
  output           tse_mac_transmit_error;
  output           tse_mac_transmit_ready_from_sa;
  output           tse_mac_transmit_startofpacket;
  output           tse_mac_transmit_valid;
  input            clk;
  input            reset_n;
  input   [ 31: 0] sgdma_tx_out_data;
  input   [  1: 0] sgdma_tx_out_empty;
  input            sgdma_tx_out_endofpacket;
  input            sgdma_tx_out_error;
  input            sgdma_tx_out_startofpacket;
  input            sgdma_tx_out_valid;
  input            tse_mac_transmit_ready;

  wire    [ 31: 0] tse_mac_transmit_data;
  wire    [  1: 0] tse_mac_transmit_empty;
  wire             tse_mac_transmit_endofpacket;
  wire             tse_mac_transmit_error;
  wire             tse_mac_transmit_ready_from_sa;
  wire             tse_mac_transmit_startofpacket;
  wire             tse_mac_transmit_valid;
  //mux tse_mac_transmit_data, which is an e_mux
  assign tse_mac_transmit_data = sgdma_tx_out_data;

  //mux tse_mac_transmit_endofpacket, which is an e_mux
  assign tse_mac_transmit_endofpacket = sgdma_tx_out_endofpacket;

  //mux tse_mac_transmit_error, which is an e_mux
  assign tse_mac_transmit_error = sgdma_tx_out_error;

  //mux tse_mac_transmit_empty, which is an e_mux
  assign tse_mac_transmit_empty = sgdma_tx_out_empty;

  //assign tse_mac_transmit_ready_from_sa = tse_mac_transmit_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_mac_transmit_ready_from_sa = tse_mac_transmit_ready;

  //mux tse_mac_transmit_startofpacket, which is an e_mux
  assign tse_mac_transmit_startofpacket = sgdma_tx_out_startofpacket;

  //mux tse_mac_transmit_valid, which is an e_mux
  assign tse_mac_transmit_valid = sgdma_tx_out_valid;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_mac_receive_arbitrator (
                                    // inputs:
                                     clk,
                                     reset_n,
                                     sgdma_rx_in_ready_from_sa,
                                     tse_mac_receive_data,
                                     tse_mac_receive_empty,
                                     tse_mac_receive_endofpacket,
                                     tse_mac_receive_error,
                                     tse_mac_receive_startofpacket,
                                     tse_mac_receive_valid,

                                    // outputs:
                                     tse_mac_receive_ready
                                  )
;

  output           tse_mac_receive_ready;
  input            clk;
  input            reset_n;
  input            sgdma_rx_in_ready_from_sa;
  input   [ 31: 0] tse_mac_receive_data;
  input   [  1: 0] tse_mac_receive_empty;
  input            tse_mac_receive_endofpacket;
  input   [  5: 0] tse_mac_receive_error;
  input            tse_mac_receive_startofpacket;
  input            tse_mac_receive_valid;

  wire             tse_mac_receive_ready;
  //mux tse_mac_receive_ready, which is an e_mux
  assign tse_mac_receive_ready = sgdma_rx_in_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_pll_s1_arbitrator (
                               // inputs:
                                clk,
                                cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave,
                                cycloneIII_3c120_niosII_standard_sopc_clock_1_out_nativeaddress,
                                cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read,
                                cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write,
                                cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata,
                                reset_n,
                                tse_pll_s1_readdata,
                                tse_pll_s1_resetrequest,

                               // outputs:
                                cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1,
                                cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1,
                                cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_data_valid_tse_pll_s1,
                                cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1,
                                d1_tse_pll_s1_end_xfer,
                                tse_pll_s1_address,
                                tse_pll_s1_chipselect,
                                tse_pll_s1_read,
                                tse_pll_s1_readdata_from_sa,
                                tse_pll_s1_reset_n,
                                tse_pll_s1_resetrequest_from_sa,
                                tse_pll_s1_write,
                                tse_pll_s1_writedata
                             )
;

  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_data_valid_tse_pll_s1;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1;
  output           d1_tse_pll_s1_end_xfer;
  output  [  2: 0] tse_pll_s1_address;
  output           tse_pll_s1_chipselect;
  output           tse_pll_s1_read;
  output  [ 15: 0] tse_pll_s1_readdata_from_sa;
  output           tse_pll_s1_reset_n;
  output           tse_pll_s1_resetrequest_from_sa;
  output           tse_pll_s1_write;
  output  [ 15: 0] tse_pll_s1_writedata;
  input            clk;
  input   [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave;
  input   [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_nativeaddress;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata;
  input            reset_n;
  input   [ 15: 0] tse_pll_s1_readdata;
  input            tse_pll_s1_resetrequest;

  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_arbiterlock;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_arbiterlock2;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_continuerequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_data_valid_tse_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_saved_grant_tse_pll_s1;
  reg              d1_reasons_to_wait;
  reg              d1_tse_pll_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tse_pll_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  2: 0] tse_pll_s1_address;
  wire             tse_pll_s1_allgrants;
  wire             tse_pll_s1_allow_new_arb_cycle;
  wire             tse_pll_s1_any_bursting_master_saved_grant;
  wire             tse_pll_s1_any_continuerequest;
  wire             tse_pll_s1_arb_counter_enable;
  reg              tse_pll_s1_arb_share_counter;
  wire             tse_pll_s1_arb_share_counter_next_value;
  wire             tse_pll_s1_arb_share_set_values;
  wire             tse_pll_s1_beginbursttransfer_internal;
  wire             tse_pll_s1_begins_xfer;
  wire             tse_pll_s1_chipselect;
  wire             tse_pll_s1_end_xfer;
  wire             tse_pll_s1_firsttransfer;
  wire             tse_pll_s1_grant_vector;
  wire             tse_pll_s1_in_a_read_cycle;
  wire             tse_pll_s1_in_a_write_cycle;
  wire             tse_pll_s1_master_qreq_vector;
  wire             tse_pll_s1_non_bursting_master_requests;
  wire             tse_pll_s1_read;
  wire    [ 15: 0] tse_pll_s1_readdata_from_sa;
  reg              tse_pll_s1_reg_firsttransfer;
  wire             tse_pll_s1_reset_n;
  wire             tse_pll_s1_resetrequest_from_sa;
  reg              tse_pll_s1_slavearbiterlockenable;
  wire             tse_pll_s1_slavearbiterlockenable2;
  wire             tse_pll_s1_unreg_firsttransfer;
  wire             tse_pll_s1_waits_for_read;
  wire             tse_pll_s1_waits_for_write;
  wire             tse_pll_s1_write;
  wire    [ 15: 0] tse_pll_s1_writedata;
  wire             wait_for_tse_pll_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tse_pll_s1_end_xfer;
    end


  assign tse_pll_s1_begins_xfer = ~d1_reasons_to_wait & ((cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1));
  //assign tse_pll_s1_readdata_from_sa = tse_pll_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_pll_s1_readdata_from_sa = tse_pll_s1_readdata;

  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1 = (1) & (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read | cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write);
  //tse_pll_s1_arb_share_counter set values, which is an e_mux
  assign tse_pll_s1_arb_share_set_values = 1;

  //tse_pll_s1_non_bursting_master_requests mux, which is an e_mux
  assign tse_pll_s1_non_bursting_master_requests = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1;

  //tse_pll_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign tse_pll_s1_any_bursting_master_saved_grant = 0;

  //tse_pll_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign tse_pll_s1_arb_share_counter_next_value = tse_pll_s1_firsttransfer ? (tse_pll_s1_arb_share_set_values - 1) : |tse_pll_s1_arb_share_counter ? (tse_pll_s1_arb_share_counter - 1) : 0;

  //tse_pll_s1_allgrants all slave grants, which is an e_mux
  assign tse_pll_s1_allgrants = |tse_pll_s1_grant_vector;

  //tse_pll_s1_end_xfer assignment, which is an e_assign
  assign tse_pll_s1_end_xfer = ~(tse_pll_s1_waits_for_read | tse_pll_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tse_pll_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tse_pll_s1 = tse_pll_s1_end_xfer & (~tse_pll_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tse_pll_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign tse_pll_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_tse_pll_s1 & tse_pll_s1_allgrants) | (end_xfer_arb_share_counter_term_tse_pll_s1 & ~tse_pll_s1_non_bursting_master_requests);

  //tse_pll_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_pll_s1_arb_share_counter <= 0;
      else if (tse_pll_s1_arb_counter_enable)
          tse_pll_s1_arb_share_counter <= tse_pll_s1_arb_share_counter_next_value;
    end


  //tse_pll_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_pll_s1_slavearbiterlockenable <= 0;
      else if ((|tse_pll_s1_master_qreq_vector & end_xfer_arb_share_counter_term_tse_pll_s1) | (end_xfer_arb_share_counter_term_tse_pll_s1 & ~tse_pll_s1_non_bursting_master_requests))
          tse_pll_s1_slavearbiterlockenable <= |tse_pll_s1_arb_share_counter_next_value;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_1/out tse_pll/s1 arbiterlock, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_arbiterlock = tse_pll_s1_slavearbiterlockenable & cycloneIII_3c120_niosII_standard_sopc_clock_1_out_continuerequest;

  //tse_pll_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tse_pll_s1_slavearbiterlockenable2 = |tse_pll_s1_arb_share_counter_next_value;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1/out tse_pll/s1 arbiterlock2, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_arbiterlock2 = tse_pll_s1_slavearbiterlockenable2 & cycloneIII_3c120_niosII_standard_sopc_clock_1_out_continuerequest;

  //tse_pll_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign tse_pll_s1_any_continuerequest = 1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_continuerequest continued request, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_continuerequest = 1;

  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1 = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1;
  //tse_pll_s1_writedata mux, which is an e_mux
  assign tse_pll_s1_writedata = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata;

  //master is always granted when requested
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1 = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1/out saved-grant tse_pll/s1, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_saved_grant_tse_pll_s1 = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1;

  //allow new arb cycle for tse_pll/s1, which is an e_assign
  assign tse_pll_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign tse_pll_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign tse_pll_s1_master_qreq_vector = 1;

  //tse_pll_s1_reset_n assignment, which is an e_assign
  assign tse_pll_s1_reset_n = reset_n;

  //assign tse_pll_s1_resetrequest_from_sa = tse_pll_s1_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_pll_s1_resetrequest_from_sa = tse_pll_s1_resetrequest;

  assign tse_pll_s1_chipselect = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1;
  //tse_pll_s1_firsttransfer first transaction, which is an e_assign
  assign tse_pll_s1_firsttransfer = tse_pll_s1_begins_xfer ? tse_pll_s1_unreg_firsttransfer : tse_pll_s1_reg_firsttransfer;

  //tse_pll_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign tse_pll_s1_unreg_firsttransfer = ~(tse_pll_s1_slavearbiterlockenable & tse_pll_s1_any_continuerequest);

  //tse_pll_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_pll_s1_reg_firsttransfer <= 1'b1;
      else if (tse_pll_s1_begins_xfer)
          tse_pll_s1_reg_firsttransfer <= tse_pll_s1_unreg_firsttransfer;
    end


  //tse_pll_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tse_pll_s1_beginbursttransfer_internal = tse_pll_s1_begins_xfer;

  //tse_pll_s1_read assignment, which is an e_mux
  assign tse_pll_s1_read = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read;

  //tse_pll_s1_write assignment, which is an e_mux
  assign tse_pll_s1_write = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write;

  //tse_pll_s1_address mux, which is an e_mux
  assign tse_pll_s1_address = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_nativeaddress;

  //d1_tse_pll_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tse_pll_s1_end_xfer <= 1;
      else 
        d1_tse_pll_s1_end_xfer <= tse_pll_s1_end_xfer;
    end


  //tse_pll_s1_waits_for_read in a cycle, which is an e_mux
  assign tse_pll_s1_waits_for_read = tse_pll_s1_in_a_read_cycle & tse_pll_s1_begins_xfer;

  //tse_pll_s1_in_a_read_cycle assignment, which is an e_assign
  assign tse_pll_s1_in_a_read_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tse_pll_s1_in_a_read_cycle;

  //tse_pll_s1_waits_for_write in a cycle, which is an e_mux
  assign tse_pll_s1_waits_for_write = tse_pll_s1_in_a_write_cycle & 0;

  //tse_pll_s1_in_a_write_cycle assignment, which is an e_assign
  assign tse_pll_s1_in_a_write_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tse_pll_s1_in_a_write_cycle;

  assign wait_for_tse_pll_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tse_pll/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tse_tx_pll_s1_arbitrator (
                                  // inputs:
                                   clk,
                                   cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave,
                                   cycloneIII_3c120_niosII_standard_sopc_clock_2_out_nativeaddress,
                                   cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read,
                                   cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write,
                                   cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata,
                                   reset_n,
                                   tse_tx_pll_s1_readdata,
                                   tse_tx_pll_s1_resetrequest,

                                  // outputs:
                                   cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1,
                                   cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1,
                                   cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_data_valid_tse_tx_pll_s1,
                                   cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1,
                                   d1_tse_tx_pll_s1_end_xfer,
                                   tse_tx_pll_s1_address,
                                   tse_tx_pll_s1_chipselect,
                                   tse_tx_pll_s1_read,
                                   tse_tx_pll_s1_readdata_from_sa,
                                   tse_tx_pll_s1_reset_n,
                                   tse_tx_pll_s1_resetrequest_from_sa,
                                   tse_tx_pll_s1_write,
                                   tse_tx_pll_s1_writedata
                                )
;

  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_data_valid_tse_tx_pll_s1;
  output           cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1;
  output           d1_tse_tx_pll_s1_end_xfer;
  output  [  2: 0] tse_tx_pll_s1_address;
  output           tse_tx_pll_s1_chipselect;
  output           tse_tx_pll_s1_read;
  output  [ 15: 0] tse_tx_pll_s1_readdata_from_sa;
  output           tse_tx_pll_s1_reset_n;
  output           tse_tx_pll_s1_resetrequest_from_sa;
  output           tse_tx_pll_s1_write;
  output  [ 15: 0] tse_tx_pll_s1_writedata;
  input            clk;
  input   [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave;
  input   [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_nativeaddress;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read;
  input            cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write;
  input   [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata;
  input            reset_n;
  input   [ 15: 0] tse_tx_pll_s1_readdata;
  input            tse_tx_pll_s1_resetrequest;

  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_arbiterlock;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_arbiterlock2;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_continuerequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_data_valid_tse_tx_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_saved_grant_tse_tx_pll_s1;
  reg              d1_reasons_to_wait;
  reg              d1_tse_tx_pll_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tse_tx_pll_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  2: 0] tse_tx_pll_s1_address;
  wire             tse_tx_pll_s1_allgrants;
  wire             tse_tx_pll_s1_allow_new_arb_cycle;
  wire             tse_tx_pll_s1_any_bursting_master_saved_grant;
  wire             tse_tx_pll_s1_any_continuerequest;
  wire             tse_tx_pll_s1_arb_counter_enable;
  reg              tse_tx_pll_s1_arb_share_counter;
  wire             tse_tx_pll_s1_arb_share_counter_next_value;
  wire             tse_tx_pll_s1_arb_share_set_values;
  wire             tse_tx_pll_s1_beginbursttransfer_internal;
  wire             tse_tx_pll_s1_begins_xfer;
  wire             tse_tx_pll_s1_chipselect;
  wire             tse_tx_pll_s1_end_xfer;
  wire             tse_tx_pll_s1_firsttransfer;
  wire             tse_tx_pll_s1_grant_vector;
  wire             tse_tx_pll_s1_in_a_read_cycle;
  wire             tse_tx_pll_s1_in_a_write_cycle;
  wire             tse_tx_pll_s1_master_qreq_vector;
  wire             tse_tx_pll_s1_non_bursting_master_requests;
  wire             tse_tx_pll_s1_read;
  wire    [ 15: 0] tse_tx_pll_s1_readdata_from_sa;
  reg              tse_tx_pll_s1_reg_firsttransfer;
  wire             tse_tx_pll_s1_reset_n;
  wire             tse_tx_pll_s1_resetrequest_from_sa;
  reg              tse_tx_pll_s1_slavearbiterlockenable;
  wire             tse_tx_pll_s1_slavearbiterlockenable2;
  wire             tse_tx_pll_s1_unreg_firsttransfer;
  wire             tse_tx_pll_s1_waits_for_read;
  wire             tse_tx_pll_s1_waits_for_write;
  wire             tse_tx_pll_s1_write;
  wire    [ 15: 0] tse_tx_pll_s1_writedata;
  wire             wait_for_tse_tx_pll_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tse_tx_pll_s1_end_xfer;
    end


  assign tse_tx_pll_s1_begins_xfer = ~d1_reasons_to_wait & ((cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1));
  //assign tse_tx_pll_s1_readdata_from_sa = tse_tx_pll_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_tx_pll_s1_readdata_from_sa = tse_tx_pll_s1_readdata;

  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1 = (1) & (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read | cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write);
  //tse_tx_pll_s1_arb_share_counter set values, which is an e_mux
  assign tse_tx_pll_s1_arb_share_set_values = 1;

  //tse_tx_pll_s1_non_bursting_master_requests mux, which is an e_mux
  assign tse_tx_pll_s1_non_bursting_master_requests = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1;

  //tse_tx_pll_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign tse_tx_pll_s1_any_bursting_master_saved_grant = 0;

  //tse_tx_pll_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign tse_tx_pll_s1_arb_share_counter_next_value = tse_tx_pll_s1_firsttransfer ? (tse_tx_pll_s1_arb_share_set_values - 1) : |tse_tx_pll_s1_arb_share_counter ? (tse_tx_pll_s1_arb_share_counter - 1) : 0;

  //tse_tx_pll_s1_allgrants all slave grants, which is an e_mux
  assign tse_tx_pll_s1_allgrants = |tse_tx_pll_s1_grant_vector;

  //tse_tx_pll_s1_end_xfer assignment, which is an e_assign
  assign tse_tx_pll_s1_end_xfer = ~(tse_tx_pll_s1_waits_for_read | tse_tx_pll_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tse_tx_pll_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tse_tx_pll_s1 = tse_tx_pll_s1_end_xfer & (~tse_tx_pll_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tse_tx_pll_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign tse_tx_pll_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_tse_tx_pll_s1 & tse_tx_pll_s1_allgrants) | (end_xfer_arb_share_counter_term_tse_tx_pll_s1 & ~tse_tx_pll_s1_non_bursting_master_requests);

  //tse_tx_pll_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_tx_pll_s1_arb_share_counter <= 0;
      else if (tse_tx_pll_s1_arb_counter_enable)
          tse_tx_pll_s1_arb_share_counter <= tse_tx_pll_s1_arb_share_counter_next_value;
    end


  //tse_tx_pll_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_tx_pll_s1_slavearbiterlockenable <= 0;
      else if ((|tse_tx_pll_s1_master_qreq_vector & end_xfer_arb_share_counter_term_tse_tx_pll_s1) | (end_xfer_arb_share_counter_term_tse_tx_pll_s1 & ~tse_tx_pll_s1_non_bursting_master_requests))
          tse_tx_pll_s1_slavearbiterlockenable <= |tse_tx_pll_s1_arb_share_counter_next_value;
    end


  //cycloneIII_3c120_niosII_standard_sopc_clock_2/out tse_tx_pll/s1 arbiterlock, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_arbiterlock = tse_tx_pll_s1_slavearbiterlockenable & cycloneIII_3c120_niosII_standard_sopc_clock_2_out_continuerequest;

  //tse_tx_pll_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tse_tx_pll_s1_slavearbiterlockenable2 = |tse_tx_pll_s1_arb_share_counter_next_value;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2/out tse_tx_pll/s1 arbiterlock2, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_arbiterlock2 = tse_tx_pll_s1_slavearbiterlockenable2 & cycloneIII_3c120_niosII_standard_sopc_clock_2_out_continuerequest;

  //tse_tx_pll_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign tse_tx_pll_s1_any_continuerequest = 1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_continuerequest continued request, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_continuerequest = 1;

  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1 = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1;
  //tse_tx_pll_s1_writedata mux, which is an e_mux
  assign tse_tx_pll_s1_writedata = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata;

  //master is always granted when requested
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1 = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2/out saved-grant tse_tx_pll/s1, which is an e_assign
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_saved_grant_tse_tx_pll_s1 = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1;

  //allow new arb cycle for tse_tx_pll/s1, which is an e_assign
  assign tse_tx_pll_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign tse_tx_pll_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign tse_tx_pll_s1_master_qreq_vector = 1;

  //tse_tx_pll_s1_reset_n assignment, which is an e_assign
  assign tse_tx_pll_s1_reset_n = reset_n;

  //assign tse_tx_pll_s1_resetrequest_from_sa = tse_tx_pll_s1_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tse_tx_pll_s1_resetrequest_from_sa = tse_tx_pll_s1_resetrequest;

  assign tse_tx_pll_s1_chipselect = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1;
  //tse_tx_pll_s1_firsttransfer first transaction, which is an e_assign
  assign tse_tx_pll_s1_firsttransfer = tse_tx_pll_s1_begins_xfer ? tse_tx_pll_s1_unreg_firsttransfer : tse_tx_pll_s1_reg_firsttransfer;

  //tse_tx_pll_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign tse_tx_pll_s1_unreg_firsttransfer = ~(tse_tx_pll_s1_slavearbiterlockenable & tse_tx_pll_s1_any_continuerequest);

  //tse_tx_pll_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tse_tx_pll_s1_reg_firsttransfer <= 1'b1;
      else if (tse_tx_pll_s1_begins_xfer)
          tse_tx_pll_s1_reg_firsttransfer <= tse_tx_pll_s1_unreg_firsttransfer;
    end


  //tse_tx_pll_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tse_tx_pll_s1_beginbursttransfer_internal = tse_tx_pll_s1_begins_xfer;

  //tse_tx_pll_s1_read assignment, which is an e_mux
  assign tse_tx_pll_s1_read = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read;

  //tse_tx_pll_s1_write assignment, which is an e_mux
  assign tse_tx_pll_s1_write = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write;

  //tse_tx_pll_s1_address mux, which is an e_mux
  assign tse_tx_pll_s1_address = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_nativeaddress;

  //d1_tse_tx_pll_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tse_tx_pll_s1_end_xfer <= 1;
      else 
        d1_tse_tx_pll_s1_end_xfer <= tse_tx_pll_s1_end_xfer;
    end


  //tse_tx_pll_s1_waits_for_read in a cycle, which is an e_mux
  assign tse_tx_pll_s1_waits_for_read = tse_tx_pll_s1_in_a_read_cycle & tse_tx_pll_s1_begins_xfer;

  //tse_tx_pll_s1_in_a_read_cycle assignment, which is an e_assign
  assign tse_tx_pll_s1_in_a_read_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tse_tx_pll_s1_in_a_read_cycle;

  //tse_tx_pll_s1_waits_for_write in a cycle, which is an e_mux
  assign tse_tx_pll_s1_waits_for_write = tse_tx_pll_s1_in_a_write_cycle & 0;

  //tse_tx_pll_s1_in_a_write_cycle assignment, which is an e_assign
  assign tse_tx_pll_s1_in_a_write_cycle = cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1 & cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tse_tx_pll_s1_in_a_write_cycle;

  assign wait_for_tse_tx_pll_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tse_tx_pll/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_reset_pll_c2_out_domain_synch_module (
                                                                                    // inputs:
                                                                                     clk,
                                                                                     data_in,
                                                                                     reset_n,

                                                                                    // outputs:
                                                                                     data_out
                                                                                  )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_reset_pll_c0_out_domain_synch_module (
                                                                                    // inputs:
                                                                                     clk,
                                                                                     data_in,
                                                                                     reset_n,

                                                                                    // outputs:
                                                                                     data_out
                                                                                  )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_reset_ddr2_sdram_phy_clk_out_domain_synch_module (
                                                                                                // inputs:
                                                                                                 clk,
                                                                                                 data_in,
                                                                                                 reset_n,

                                                                                                // outputs:
                                                                                                 data_out
                                                                                              )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_reset_clk_domain_synch_module (
                                                                             // inputs:
                                                                              clk,
                                                                              data_in,
                                                                              reset_n,

                                                                             // outputs:
                                                                              data_out
                                                                           )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc_reset_clk_to_tse_pll_domain_synch_module (
                                                                                        // inputs:
                                                                                         clk,
                                                                                         data_in,
                                                                                         reset_n,

                                                                                        // outputs:
                                                                                         data_out
                                                                                      )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cycloneIII_3c120_niosII_standard_sopc (
                                               // 1) global signals:
                                                clk,
                                                clk_125,
                                                clk_to_tse_pll,
                                                ddr2_sdram_aux_full_rate_clk_out,
                                                ddr2_sdram_aux_half_rate_clk_out,
                                                ddr2_sdram_phy_clk_out,
                                                pll_c0_out,
                                                pll_c2_out,
                                                pll_c3_out,
                                                pll_c4_out,
                                                reset_n,
                                                tse_pll_c0_out,
                                                tse_tx_pll_c0_out,
                                                tse_tx_pll_c1_out,
                                                tse_tx_pll_c2_out,
                                                tse_tx_pll_c3_out,

                                               // the_button_pio
                                                in_port_to_the_button_pio,

                                               // the_ddr2_sdram
                                                global_reset_n_to_the_ddr2_sdram,
                                                local_init_done_from_the_ddr2_sdram,
                                                local_refresh_ack_from_the_ddr2_sdram,
                                                local_wdata_req_from_the_ddr2_sdram,
                                                mem_addr_from_the_ddr2_sdram,
                                                mem_ba_from_the_ddr2_sdram,
                                                mem_cas_n_from_the_ddr2_sdram,
                                                mem_cke_from_the_ddr2_sdram,
                                                mem_clk_n_to_and_from_the_ddr2_sdram,
                                                mem_clk_to_and_from_the_ddr2_sdram,
                                                mem_cs_n_from_the_ddr2_sdram,
                                                mem_dm_from_the_ddr2_sdram,
                                                mem_dq_to_and_from_the_ddr2_sdram,
                                                mem_dqs_to_and_from_the_ddr2_sdram,
                                                mem_odt_from_the_ddr2_sdram,
                                                mem_ras_n_from_the_ddr2_sdram,
                                                mem_we_n_from_the_ddr2_sdram,
                                                reset_phy_clk_n_from_the_ddr2_sdram,

                                               // the_flash_tristate_bridge_avalon_slave
                                                cs_n_to_the_max2,
                                                flash_tristate_bridge_address,
                                                flash_tristate_bridge_data,
                                                oe_n_to_the_max2,
                                                read_n_to_the_ext_flash,
                                                select_n_to_the_ext_flash,
                                                we_n_to_the_max2,
                                                write_n_to_the_ext_flash,

                                               // the_led_pio
                                                out_port_from_the_led_pio,

                                               // the_pll
                                                locked_from_the_pll,

                                               // the_tse_mac
                                                ena_10_from_the_tse_mac,
                                                eth_mode_from_the_tse_mac,
                                                mdc_from_the_tse_mac,
                                                mdio_in_to_the_tse_mac,
                                                mdio_oen_from_the_tse_mac,
                                                mdio_out_from_the_tse_mac,
                                                rgmii_in_to_the_tse_mac,
                                                rgmii_out_from_the_tse_mac,
                                                rx_clk_to_the_tse_mac,
                                                rx_control_to_the_tse_mac,
                                                set_1000_to_the_tse_mac,
                                                set_10_to_the_tse_mac,
                                                tx_clk_to_the_tse_mac,
                                                tx_control_from_the_tse_mac,

                                               // the_tse_pll
                                                locked_from_the_tse_pll,

                                               // the_tse_tx_pll
                                                locked_from_the_tse_tx_pll
                                             )
;

  output           cs_n_to_the_max2;
  output           ddr2_sdram_aux_full_rate_clk_out;
  output           ddr2_sdram_aux_half_rate_clk_out;
  output           ddr2_sdram_phy_clk_out;
  output           ena_10_from_the_tse_mac;
  output           eth_mode_from_the_tse_mac;
  output  [ 25: 0] flash_tristate_bridge_address;
  inout   [ 31: 0] flash_tristate_bridge_data;
  output           local_init_done_from_the_ddr2_sdram;
  output           local_refresh_ack_from_the_ddr2_sdram;
  output           local_wdata_req_from_the_ddr2_sdram;
  output           locked_from_the_pll;
  output           locked_from_the_tse_pll;
  output           locked_from_the_tse_tx_pll;
  output           mdc_from_the_tse_mac;
  output           mdio_oen_from_the_tse_mac;
  output           mdio_out_from_the_tse_mac;
  output  [ 12: 0] mem_addr_from_the_ddr2_sdram;
  output  [  1: 0] mem_ba_from_the_ddr2_sdram;
  output           mem_cas_n_from_the_ddr2_sdram;
  output           mem_cke_from_the_ddr2_sdram;
  inout            mem_clk_n_to_and_from_the_ddr2_sdram;
  inout            mem_clk_to_and_from_the_ddr2_sdram;
  output           mem_cs_n_from_the_ddr2_sdram;
  output  [  1: 0] mem_dm_from_the_ddr2_sdram;
  inout   [ 15: 0] mem_dq_to_and_from_the_ddr2_sdram;
  inout   [  1: 0] mem_dqs_to_and_from_the_ddr2_sdram;
  output           mem_odt_from_the_ddr2_sdram;
  output           mem_ras_n_from_the_ddr2_sdram;
  output           mem_we_n_from_the_ddr2_sdram;
  output           oe_n_to_the_max2;
  output  [  7: 0] out_port_from_the_led_pio;
  output           pll_c0_out;
  output           pll_c2_out;
  output           pll_c3_out;
  output           pll_c4_out;
  output           read_n_to_the_ext_flash;
  output           reset_phy_clk_n_from_the_ddr2_sdram;
  output  [  3: 0] rgmii_out_from_the_tse_mac;
  output           select_n_to_the_ext_flash;
  output           tse_pll_c0_out;
  output           tse_tx_pll_c0_out;
  output           tse_tx_pll_c1_out;
  output           tse_tx_pll_c2_out;
  output           tse_tx_pll_c3_out;
  output           tx_control_from_the_tse_mac;
  output           we_n_to_the_max2;
  output           write_n_to_the_ext_flash;
  input            clk;
  input            clk_125;
  input            clk_to_tse_pll;
  input            global_reset_n_to_the_ddr2_sdram;
  input   [  3: 0] in_port_to_the_button_pio;
  input            mdio_in_to_the_tse_mac;
  input            reset_n;
  input   [  3: 0] rgmii_in_to_the_tse_mac;
  input            rx_clk_to_the_tse_mac;
  input            rx_control_to_the_tse_mac;
  input            set_1000_to_the_tse_mac;
  input            set_10_to_the_tse_mac;
  input            tx_clk_to_the_tse_mac;

  wire    [  1: 0] button_pio_s1_address;
  wire             button_pio_s1_chipselect;
  wire             button_pio_s1_irq;
  wire             button_pio_s1_irq_from_sa;
  wire    [ 31: 0] button_pio_s1_readdata;
  wire    [ 31: 0] button_pio_s1_readdata_from_sa;
  wire             button_pio_s1_reset_n;
  wire             button_pio_s1_write_n;
  wire    [ 31: 0] button_pio_s1_writedata;
  wire             clk_125_reset_n;
  wire             clk_reset_n;
  wire             clk_to_tse_pll_reset_n;
  wire    [ 28: 0] cpu_data_master_address;
  wire    [ 28: 0] cpu_data_master_address_to_slave;
  wire    [  3: 0] cpu_data_master_byteenable;
  wire             cpu_data_master_debugaccess;
  wire             cpu_data_master_granted_cpu_ddr_clock_bridge_s1;
  wire             cpu_data_master_granted_cpu_jtag_debug_module;
  wire             cpu_data_master_granted_descriptor_memory_s1;
  wire             cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_data_master_granted_sgdma_rx_csr;
  wire             cpu_data_master_granted_sgdma_tx_csr;
  wire             cpu_data_master_granted_slow_peripheral_bridge_s1;
  wire             cpu_data_master_granted_tse_mac_control_port;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_latency_counter;
  wire             cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1;
  wire             cpu_data_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_data_master_qualified_request_descriptor_memory_s1;
  wire             cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_data_master_qualified_request_sgdma_rx_csr;
  wire             cpu_data_master_qualified_request_sgdma_tx_csr;
  wire             cpu_data_master_qualified_request_slow_peripheral_bridge_s1;
  wire             cpu_data_master_qualified_request_tse_mac_control_port;
  wire             cpu_data_master_read;
  wire             cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1;
  wire             cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  wire             cpu_data_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_data_master_read_data_valid_descriptor_memory_s1;
  wire             cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  wire             cpu_data_master_read_data_valid_sgdma_rx_csr;
  wire             cpu_data_master_read_data_valid_sgdma_tx_csr;
  wire             cpu_data_master_read_data_valid_slow_peripheral_bridge_s1;
  wire             cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register;
  wire             cpu_data_master_read_data_valid_tse_mac_control_port;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_requests_cpu_ddr_clock_bridge_s1;
  wire             cpu_data_master_requests_cpu_jtag_debug_module;
  wire             cpu_data_master_requests_descriptor_memory_s1;
  wire             cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_data_master_requests_sgdma_rx_csr;
  wire             cpu_data_master_requests_sgdma_tx_csr;
  wire             cpu_data_master_requests_slow_peripheral_bridge_s1;
  wire             cpu_data_master_requests_tse_mac_control_port;
  wire             cpu_data_master_waitrequest;
  wire             cpu_data_master_write;
  wire    [ 31: 0] cpu_data_master_writedata;
  wire    [ 25: 0] cpu_ddr_clock_bridge_m1_address;
  wire    [ 25: 0] cpu_ddr_clock_bridge_m1_address_to_slave;
  wire    [  3: 0] cpu_ddr_clock_bridge_m1_byteenable;
  wire             cpu_ddr_clock_bridge_m1_endofpacket;
  wire             cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1;
  wire             cpu_ddr_clock_bridge_m1_latency_counter;
  wire    [ 23: 0] cpu_ddr_clock_bridge_m1_nativeaddress;
  wire             cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1;
  wire             cpu_ddr_clock_bridge_m1_read;
  wire             cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1;
  wire             cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register;
  wire    [ 31: 0] cpu_ddr_clock_bridge_m1_readdata;
  wire             cpu_ddr_clock_bridge_m1_readdatavalid;
  wire             cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1;
  wire             cpu_ddr_clock_bridge_m1_reset_n;
  wire             cpu_ddr_clock_bridge_m1_waitrequest;
  wire             cpu_ddr_clock_bridge_m1_write;
  wire    [ 31: 0] cpu_ddr_clock_bridge_m1_writedata;
  wire    [ 23: 0] cpu_ddr_clock_bridge_s1_address;
  wire    [  3: 0] cpu_ddr_clock_bridge_s1_byteenable;
  wire             cpu_ddr_clock_bridge_s1_endofpacket;
  wire             cpu_ddr_clock_bridge_s1_endofpacket_from_sa;
  wire    [ 23: 0] cpu_ddr_clock_bridge_s1_nativeaddress;
  wire             cpu_ddr_clock_bridge_s1_read;
  wire    [ 31: 0] cpu_ddr_clock_bridge_s1_readdata;
  wire    [ 31: 0] cpu_ddr_clock_bridge_s1_readdata_from_sa;
  wire             cpu_ddr_clock_bridge_s1_readdatavalid;
  wire             cpu_ddr_clock_bridge_s1_reset_n;
  wire             cpu_ddr_clock_bridge_s1_waitrequest;
  wire             cpu_ddr_clock_bridge_s1_waitrequest_from_sa;
  wire             cpu_ddr_clock_bridge_s1_write;
  wire    [ 31: 0] cpu_ddr_clock_bridge_s1_writedata;
  wire    [ 28: 0] cpu_instruction_master_address;
  wire    [ 28: 0] cpu_instruction_master_address_to_slave;
  wire             cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1;
  wire             cpu_instruction_master_granted_cpu_jtag_debug_module;
  wire             cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_latency_counter;
  wire             cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1;
  wire             cpu_instruction_master_qualified_request_cpu_jtag_debug_module;
  wire             cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_read;
  wire             cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1;
  wire             cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  wire             cpu_instruction_master_read_data_valid_cpu_jtag_debug_module;
  wire             cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1;
  wire             cpu_instruction_master_requests_cpu_jtag_debug_module;
  wire             cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1;
  wire             cpu_instruction_master_waitrequest;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire             cpu_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  wire             cs_n_to_the_max2;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_address;
  wire    [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_byteenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa;
  wire    [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_nativeaddress;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_read;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reset_n;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_in_write;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_in_writedata;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave;
  wire    [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_endofpacket;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1;
  wire    [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_nativeaddress;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_data_valid_pll_s1;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_readdata;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_reset_n;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_waitrequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_address;
  wire    [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_byteenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa;
  wire    [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_nativeaddress;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_read;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reset_n;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_in_write;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_in_writedata;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave;
  wire    [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_endofpacket;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1;
  wire    [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_nativeaddress;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_data_valid_tse_pll_s1;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_readdata;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_reset_n;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_waitrequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_address;
  wire    [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_byteenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa;
  wire    [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_nativeaddress;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_read;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reset_n;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_in_write;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_in_writedata;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address;
  wire    [  3: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave;
  wire    [  1: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_endofpacket;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1;
  wire    [  2: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_nativeaddress;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_data_valid_tse_tx_pll_s1;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_readdata;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_reset_n;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_waitrequest;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write;
  wire    [ 15: 0] cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata;
  wire             d1_button_pio_s1_end_xfer;
  wire             d1_cpu_ddr_clock_bridge_s1_end_xfer;
  wire             d1_cpu_jtag_debug_module_end_xfer;
  wire             d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer;
  wire             d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer;
  wire             d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer;
  wire             d1_ddr2_sdram_s1_end_xfer;
  wire             d1_descriptor_memory_s1_end_xfer;
  wire             d1_flash_tristate_bridge_avalon_slave_end_xfer;
  wire             d1_high_res_timer_s1_end_xfer;
  wire             d1_jtag_uart_avalon_jtag_slave_end_xfer;
  wire             d1_led_pio_s1_end_xfer;
  wire             d1_performance_counter_control_slave_end_xfer;
  wire             d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer;
  wire             d1_pll_s1_end_xfer;
  wire             d1_sgdma_rx_csr_end_xfer;
  wire             d1_sgdma_tx_csr_end_xfer;
  wire             d1_slow_peripheral_bridge_s1_end_xfer;
  wire             d1_sys_clk_timer_s1_end_xfer;
  wire             d1_sysid_control_slave_end_xfer;
  wire             d1_tse_mac_control_port_end_xfer;
  wire             d1_tse_pll_s1_end_xfer;
  wire             d1_tse_tx_pll_s1_end_xfer;
  wire             ddr2_sdram_aux_full_rate_clk_out;
  wire             ddr2_sdram_aux_half_rate_clk_out;
  wire             ddr2_sdram_phy_clk_out;
  wire             ddr2_sdram_phy_clk_out_reset_n;
  wire    [ 23: 0] ddr2_sdram_s1_address;
  wire             ddr2_sdram_s1_beginbursttransfer;
  wire    [  2: 0] ddr2_sdram_s1_burstcount;
  wire    [  3: 0] ddr2_sdram_s1_byteenable;
  wire             ddr2_sdram_s1_read;
  wire    [ 31: 0] ddr2_sdram_s1_readdata;
  wire    [ 31: 0] ddr2_sdram_s1_readdata_from_sa;
  wire             ddr2_sdram_s1_readdatavalid;
  wire             ddr2_sdram_s1_resetrequest_n;
  wire             ddr2_sdram_s1_resetrequest_n_from_sa;
  wire             ddr2_sdram_s1_waitrequest_n;
  wire             ddr2_sdram_s1_waitrequest_n_from_sa;
  wire             ddr2_sdram_s1_write;
  wire    [ 31: 0] ddr2_sdram_s1_writedata;
  wire    [  9: 0] descriptor_memory_s1_address;
  wire    [  3: 0] descriptor_memory_s1_byteenable;
  wire             descriptor_memory_s1_chipselect;
  wire             descriptor_memory_s1_clken;
  wire    [ 31: 0] descriptor_memory_s1_readdata;
  wire    [ 31: 0] descriptor_memory_s1_readdata_from_sa;
  wire             descriptor_memory_s1_reset;
  wire             descriptor_memory_s1_write;
  wire    [ 31: 0] descriptor_memory_s1_writedata;
  wire             ena_10_from_the_tse_mac;
  wire             eth_mode_from_the_tse_mac;
  wire             ext_flash_s1_wait_counter_eq_0;
  wire    [ 25: 0] flash_tristate_bridge_address;
  wire    [ 31: 0] flash_tristate_bridge_data;
  wire    [  2: 0] high_res_timer_s1_address;
  wire             high_res_timer_s1_chipselect;
  wire             high_res_timer_s1_irq;
  wire             high_res_timer_s1_irq_from_sa;
  wire    [ 15: 0] high_res_timer_s1_readdata;
  wire    [ 15: 0] high_res_timer_s1_readdata_from_sa;
  wire             high_res_timer_s1_reset_n;
  wire             high_res_timer_s1_write_n;
  wire    [ 15: 0] high_res_timer_s1_writedata;
  wire    [ 31: 0] incoming_flash_tristate_bridge_data;
  wire    [ 15: 0] incoming_flash_tristate_bridge_data_with_Xs_converted_to_0;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_irq;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  wire             jtag_uart_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire    [  1: 0] led_pio_s1_address;
  wire             led_pio_s1_chipselect;
  wire    [ 31: 0] led_pio_s1_readdata;
  wire    [ 31: 0] led_pio_s1_readdata_from_sa;
  wire             led_pio_s1_reset_n;
  wire             led_pio_s1_write_n;
  wire    [ 31: 0] led_pio_s1_writedata;
  wire             local_init_done_from_the_ddr2_sdram;
  wire             local_refresh_ack_from_the_ddr2_sdram;
  wire             local_wdata_req_from_the_ddr2_sdram;
  wire             locked_from_the_pll;
  wire             locked_from_the_tse_pll;
  wire             locked_from_the_tse_tx_pll;
  wire             max2_s1_wait_counter_eq_0;
  wire             mdc_from_the_tse_mac;
  wire             mdio_oen_from_the_tse_mac;
  wire             mdio_out_from_the_tse_mac;
  wire    [ 12: 0] mem_addr_from_the_ddr2_sdram;
  wire    [  1: 0] mem_ba_from_the_ddr2_sdram;
  wire             mem_cas_n_from_the_ddr2_sdram;
  wire             mem_cke_from_the_ddr2_sdram;
  wire             mem_clk_n_to_and_from_the_ddr2_sdram;
  wire             mem_clk_to_and_from_the_ddr2_sdram;
  wire             mem_cs_n_from_the_ddr2_sdram;
  wire    [  1: 0] mem_dm_from_the_ddr2_sdram;
  wire    [ 15: 0] mem_dq_to_and_from_the_ddr2_sdram;
  wire    [  1: 0] mem_dqs_to_and_from_the_ddr2_sdram;
  wire             mem_odt_from_the_ddr2_sdram;
  wire             mem_ras_n_from_the_ddr2_sdram;
  wire             mem_we_n_from_the_ddr2_sdram;
  wire             oe_n_to_the_max2;
  wire             out_clk_ddr2_sdram_aux_full_rate_clk;
  wire             out_clk_ddr2_sdram_aux_half_rate_clk;
  wire             out_clk_ddr2_sdram_phy_clk;
  wire             out_clk_pll_c0;
  wire             out_clk_pll_c2;
  wire             out_clk_pll_c3;
  wire             out_clk_pll_c4;
  wire             out_clk_tse_pll_c0;
  wire             out_clk_tse_tx_pll_c0;
  wire             out_clk_tse_tx_pll_c1;
  wire             out_clk_tse_tx_pll_c2;
  wire             out_clk_tse_tx_pll_c3;
  wire    [  7: 0] out_port_from_the_led_pio;
  wire    [  2: 0] performance_counter_control_slave_address;
  wire             performance_counter_control_slave_begintransfer;
  wire    [ 31: 0] performance_counter_control_slave_readdata;
  wire    [ 31: 0] performance_counter_control_slave_readdata_from_sa;
  wire             performance_counter_control_slave_reset_n;
  wire             performance_counter_control_slave_write;
  wire    [ 31: 0] performance_counter_control_slave_writedata;
  wire    [ 26: 0] pipeline_bridge_before_tristate_bridge_m1_address;
  wire    [ 26: 0] pipeline_bridge_before_tristate_bridge_m1_address_to_slave;
  wire             pipeline_bridge_before_tristate_bridge_m1_burstcount;
  wire    [  3: 0] pipeline_bridge_before_tristate_bridge_m1_byteenable;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_chipselect;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_address;
  wire    [ 15: 0] pipeline_bridge_before_tristate_bridge_m1_dbs_write_16;
  wire             pipeline_bridge_before_tristate_bridge_m1_debugaccess;
  wire             pipeline_bridge_before_tristate_bridge_m1_endofpacket;
  wire             pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1;
  wire    [  1: 0] pipeline_bridge_before_tristate_bridge_m1_latency_counter;
  wire             pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_read;
  wire             pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1;
  wire    [ 31: 0] pipeline_bridge_before_tristate_bridge_m1_readdata;
  wire             pipeline_bridge_before_tristate_bridge_m1_readdatavalid;
  wire             pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1;
  wire             pipeline_bridge_before_tristate_bridge_m1_waitrequest;
  wire             pipeline_bridge_before_tristate_bridge_m1_write;
  wire    [ 31: 0] pipeline_bridge_before_tristate_bridge_m1_writedata;
  wire    [ 24: 0] pipeline_bridge_before_tristate_bridge_s1_address;
  wire             pipeline_bridge_before_tristate_bridge_s1_arbiterlock;
  wire             pipeline_bridge_before_tristate_bridge_s1_arbiterlock2;
  wire             pipeline_bridge_before_tristate_bridge_s1_burstcount;
  wire    [  3: 0] pipeline_bridge_before_tristate_bridge_s1_byteenable;
  wire             pipeline_bridge_before_tristate_bridge_s1_chipselect;
  wire             pipeline_bridge_before_tristate_bridge_s1_debugaccess;
  wire             pipeline_bridge_before_tristate_bridge_s1_endofpacket;
  wire             pipeline_bridge_before_tristate_bridge_s1_endofpacket_from_sa;
  wire    [ 24: 0] pipeline_bridge_before_tristate_bridge_s1_nativeaddress;
  wire             pipeline_bridge_before_tristate_bridge_s1_read;
  wire    [ 31: 0] pipeline_bridge_before_tristate_bridge_s1_readdata;
  wire    [ 31: 0] pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa;
  wire             pipeline_bridge_before_tristate_bridge_s1_readdatavalid;
  wire             pipeline_bridge_before_tristate_bridge_s1_reset_n;
  wire             pipeline_bridge_before_tristate_bridge_s1_waitrequest;
  wire             pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa;
  wire             pipeline_bridge_before_tristate_bridge_s1_write;
  wire    [ 31: 0] pipeline_bridge_before_tristate_bridge_s1_writedata;
  wire             pll_c0_out;
  wire             pll_c0_out_reset_n;
  wire             pll_c2_out;
  wire             pll_c2_out_reset_n;
  wire             pll_c3_out;
  wire             pll_c4_out;
  wire    [  2: 0] pll_s1_address;
  wire             pll_s1_chipselect;
  wire             pll_s1_read;
  wire    [ 15: 0] pll_s1_readdata;
  wire    [ 15: 0] pll_s1_readdata_from_sa;
  wire             pll_s1_reset_n;
  wire             pll_s1_resetrequest;
  wire             pll_s1_resetrequest_from_sa;
  wire             pll_s1_write;
  wire    [ 15: 0] pll_s1_writedata;
  wire             read_n_to_the_ext_flash;
  wire             reset_n_sources;
  wire             reset_phy_clk_n_from_the_ddr2_sdram;
  wire    [  3: 0] rgmii_out_from_the_tse_mac;
  wire             select_n_to_the_ext_flash;
  wire    [  3: 0] sgdma_rx_csr_address;
  wire             sgdma_rx_csr_chipselect;
  wire             sgdma_rx_csr_irq;
  wire             sgdma_rx_csr_irq_from_sa;
  wire             sgdma_rx_csr_read;
  wire    [ 31: 0] sgdma_rx_csr_readdata;
  wire    [ 31: 0] sgdma_rx_csr_readdata_from_sa;
  wire             sgdma_rx_csr_reset_n;
  wire             sgdma_rx_csr_write;
  wire    [ 31: 0] sgdma_rx_csr_writedata;
  wire    [ 31: 0] sgdma_rx_descriptor_read_address;
  wire    [ 31: 0] sgdma_rx_descriptor_read_address_to_slave;
  wire             sgdma_rx_descriptor_read_granted_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_latency_counter;
  wire             sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_read;
  wire             sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;
  wire    [ 31: 0] sgdma_rx_descriptor_read_readdata;
  wire             sgdma_rx_descriptor_read_readdatavalid;
  wire             sgdma_rx_descriptor_read_requests_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_read_waitrequest;
  wire    [ 31: 0] sgdma_rx_descriptor_write_address;
  wire    [ 31: 0] sgdma_rx_descriptor_write_address_to_slave;
  wire             sgdma_rx_descriptor_write_granted_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_requests_descriptor_memory_s1;
  wire             sgdma_rx_descriptor_write_waitrequest;
  wire             sgdma_rx_descriptor_write_write;
  wire    [ 31: 0] sgdma_rx_descriptor_write_writedata;
  wire    [ 31: 0] sgdma_rx_in_data;
  wire    [  1: 0] sgdma_rx_in_empty;
  wire             sgdma_rx_in_endofpacket;
  wire    [  5: 0] sgdma_rx_in_error;
  wire             sgdma_rx_in_ready;
  wire             sgdma_rx_in_ready_from_sa;
  wire             sgdma_rx_in_startofpacket;
  wire             sgdma_rx_in_valid;
  wire    [ 31: 0] sgdma_rx_m_write_address;
  wire    [ 31: 0] sgdma_rx_m_write_address_to_slave;
  wire    [  3: 0] sgdma_rx_m_write_byteenable;
  wire             sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1;
  wire             sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1;
  wire             sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1;
  wire             sgdma_rx_m_write_waitrequest;
  wire             sgdma_rx_m_write_write;
  wire    [ 31: 0] sgdma_rx_m_write_writedata;
  wire    [  3: 0] sgdma_tx_csr_address;
  wire             sgdma_tx_csr_chipselect;
  wire             sgdma_tx_csr_irq;
  wire             sgdma_tx_csr_irq_from_sa;
  wire             sgdma_tx_csr_read;
  wire    [ 31: 0] sgdma_tx_csr_readdata;
  wire    [ 31: 0] sgdma_tx_csr_readdata_from_sa;
  wire             sgdma_tx_csr_reset_n;
  wire             sgdma_tx_csr_write;
  wire    [ 31: 0] sgdma_tx_csr_writedata;
  wire    [ 31: 0] sgdma_tx_descriptor_read_address;
  wire    [ 31: 0] sgdma_tx_descriptor_read_address_to_slave;
  wire             sgdma_tx_descriptor_read_granted_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_latency_counter;
  wire             sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_read;
  wire             sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;
  wire    [ 31: 0] sgdma_tx_descriptor_read_readdata;
  wire             sgdma_tx_descriptor_read_readdatavalid;
  wire             sgdma_tx_descriptor_read_requests_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_read_waitrequest;
  wire    [ 31: 0] sgdma_tx_descriptor_write_address;
  wire    [ 31: 0] sgdma_tx_descriptor_write_address_to_slave;
  wire             sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
  wire             sgdma_tx_descriptor_write_waitrequest;
  wire             sgdma_tx_descriptor_write_write;
  wire    [ 31: 0] sgdma_tx_descriptor_write_writedata;
  wire    [ 31: 0] sgdma_tx_m_read_address;
  wire    [ 31: 0] sgdma_tx_m_read_address_to_slave;
  wire             sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_latency_counter;
  wire             sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_read;
  wire             sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register;
  wire    [ 31: 0] sgdma_tx_m_read_readdata;
  wire             sgdma_tx_m_read_readdatavalid;
  wire             sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1;
  wire             sgdma_tx_m_read_waitrequest;
  wire    [ 31: 0] sgdma_tx_out_data;
  wire    [  1: 0] sgdma_tx_out_empty;
  wire             sgdma_tx_out_endofpacket;
  wire             sgdma_tx_out_error;
  wire             sgdma_tx_out_ready;
  wire             sgdma_tx_out_startofpacket;
  wire             sgdma_tx_out_valid;
  wire    [  7: 0] slow_peripheral_bridge_m1_address;
  wire    [  7: 0] slow_peripheral_bridge_m1_address_to_slave;
  wire    [  3: 0] slow_peripheral_bridge_m1_byteenable;
  wire             slow_peripheral_bridge_m1_endofpacket;
  wire             slow_peripheral_bridge_m1_granted_button_pio_s1;
  wire             slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  wire             slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  wire             slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  wire             slow_peripheral_bridge_m1_granted_high_res_timer_s1;
  wire             slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  wire             slow_peripheral_bridge_m1_granted_led_pio_s1;
  wire             slow_peripheral_bridge_m1_granted_performance_counter_control_slave;
  wire             slow_peripheral_bridge_m1_granted_sys_clk_timer_s1;
  wire             slow_peripheral_bridge_m1_granted_sysid_control_slave;
  wire             slow_peripheral_bridge_m1_latency_counter;
  wire    [  5: 0] slow_peripheral_bridge_m1_nativeaddress;
  wire             slow_peripheral_bridge_m1_qualified_request_button_pio_s1;
  wire             slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  wire             slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  wire             slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  wire             slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1;
  wire             slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             slow_peripheral_bridge_m1_qualified_request_led_pio_s1;
  wire             slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave;
  wire             slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1;
  wire             slow_peripheral_bridge_m1_qualified_request_sysid_control_slave;
  wire             slow_peripheral_bridge_m1_read;
  wire             slow_peripheral_bridge_m1_read_data_valid_button_pio_s1;
  wire             slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  wire             slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  wire             slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  wire             slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1;
  wire             slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             slow_peripheral_bridge_m1_read_data_valid_led_pio_s1;
  wire             slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave;
  wire             slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1;
  wire             slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave;
  wire    [ 31: 0] slow_peripheral_bridge_m1_readdata;
  wire             slow_peripheral_bridge_m1_readdatavalid;
  wire             slow_peripheral_bridge_m1_requests_button_pio_s1;
  wire             slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in;
  wire             slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in;
  wire             slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in;
  wire             slow_peripheral_bridge_m1_requests_high_res_timer_s1;
  wire             slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  wire             slow_peripheral_bridge_m1_requests_led_pio_s1;
  wire             slow_peripheral_bridge_m1_requests_performance_counter_control_slave;
  wire             slow_peripheral_bridge_m1_requests_sys_clk_timer_s1;
  wire             slow_peripheral_bridge_m1_requests_sysid_control_slave;
  wire             slow_peripheral_bridge_m1_reset_n;
  wire             slow_peripheral_bridge_m1_waitrequest;
  wire             slow_peripheral_bridge_m1_write;
  wire    [ 31: 0] slow_peripheral_bridge_m1_writedata;
  wire    [  5: 0] slow_peripheral_bridge_s1_address;
  wire    [  3: 0] slow_peripheral_bridge_s1_byteenable;
  wire             slow_peripheral_bridge_s1_endofpacket;
  wire             slow_peripheral_bridge_s1_endofpacket_from_sa;
  wire    [  5: 0] slow_peripheral_bridge_s1_nativeaddress;
  wire             slow_peripheral_bridge_s1_read;
  wire    [ 31: 0] slow_peripheral_bridge_s1_readdata;
  wire    [ 31: 0] slow_peripheral_bridge_s1_readdata_from_sa;
  wire             slow_peripheral_bridge_s1_readdatavalid;
  wire             slow_peripheral_bridge_s1_reset_n;
  wire             slow_peripheral_bridge_s1_waitrequest;
  wire             slow_peripheral_bridge_s1_waitrequest_from_sa;
  wire             slow_peripheral_bridge_s1_write;
  wire    [ 31: 0] slow_peripheral_bridge_s1_writedata;
  wire    [  2: 0] sys_clk_timer_s1_address;
  wire             sys_clk_timer_s1_chipselect;
  wire             sys_clk_timer_s1_irq;
  wire             sys_clk_timer_s1_irq_from_sa;
  wire    [ 15: 0] sys_clk_timer_s1_readdata;
  wire    [ 15: 0] sys_clk_timer_s1_readdata_from_sa;
  wire             sys_clk_timer_s1_reset_n;
  wire             sys_clk_timer_s1_write_n;
  wire    [ 15: 0] sys_clk_timer_s1_writedata;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_clock;
  wire    [ 31: 0] sysid_control_slave_readdata;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  wire             sysid_control_slave_reset_n;
  wire    [  7: 0] tse_mac_control_port_address;
  wire             tse_mac_control_port_read;
  wire    [ 31: 0] tse_mac_control_port_readdata;
  wire    [ 31: 0] tse_mac_control_port_readdata_from_sa;
  wire             tse_mac_control_port_reset;
  wire             tse_mac_control_port_waitrequest;
  wire             tse_mac_control_port_waitrequest_from_sa;
  wire             tse_mac_control_port_write;
  wire    [ 31: 0] tse_mac_control_port_writedata;
  wire    [ 31: 0] tse_mac_receive_data;
  wire    [  1: 0] tse_mac_receive_empty;
  wire             tse_mac_receive_endofpacket;
  wire    [  5: 0] tse_mac_receive_error;
  wire             tse_mac_receive_ready;
  wire             tse_mac_receive_startofpacket;
  wire             tse_mac_receive_valid;
  wire    [ 31: 0] tse_mac_transmit_data;
  wire    [  1: 0] tse_mac_transmit_empty;
  wire             tse_mac_transmit_endofpacket;
  wire             tse_mac_transmit_error;
  wire             tse_mac_transmit_ready;
  wire             tse_mac_transmit_ready_from_sa;
  wire             tse_mac_transmit_startofpacket;
  wire             tse_mac_transmit_valid;
  wire             tse_pll_c0_out;
  wire    [  2: 0] tse_pll_s1_address;
  wire             tse_pll_s1_chipselect;
  wire             tse_pll_s1_read;
  wire    [ 15: 0] tse_pll_s1_readdata;
  wire    [ 15: 0] tse_pll_s1_readdata_from_sa;
  wire             tse_pll_s1_reset_n;
  wire             tse_pll_s1_resetrequest;
  wire             tse_pll_s1_resetrequest_from_sa;
  wire             tse_pll_s1_write;
  wire    [ 15: 0] tse_pll_s1_writedata;
  wire             tse_tx_pll_c0_out;
  wire             tse_tx_pll_c1_out;
  wire             tse_tx_pll_c2_out;
  wire             tse_tx_pll_c3_out;
  wire    [  2: 0] tse_tx_pll_s1_address;
  wire             tse_tx_pll_s1_chipselect;
  wire             tse_tx_pll_s1_read;
  wire    [ 15: 0] tse_tx_pll_s1_readdata;
  wire    [ 15: 0] tse_tx_pll_s1_readdata_from_sa;
  wire             tse_tx_pll_s1_reset_n;
  wire             tse_tx_pll_s1_resetrequest;
  wire             tse_tx_pll_s1_resetrequest_from_sa;
  wire             tse_tx_pll_s1_write;
  wire    [ 15: 0] tse_tx_pll_s1_writedata;
  wire             tx_control_from_the_tse_mac;
  wire             we_n_to_the_max2;
  wire             write_n_to_the_ext_flash;
  button_pio_s1_arbitrator the_button_pio_s1
    (
      .button_pio_s1_address                                     (button_pio_s1_address),
      .button_pio_s1_chipselect                                  (button_pio_s1_chipselect),
      .button_pio_s1_irq                                         (button_pio_s1_irq),
      .button_pio_s1_irq_from_sa                                 (button_pio_s1_irq_from_sa),
      .button_pio_s1_readdata                                    (button_pio_s1_readdata),
      .button_pio_s1_readdata_from_sa                            (button_pio_s1_readdata_from_sa),
      .button_pio_s1_reset_n                                     (button_pio_s1_reset_n),
      .button_pio_s1_write_n                                     (button_pio_s1_write_n),
      .button_pio_s1_writedata                                   (button_pio_s1_writedata),
      .clk                                                       (pll_c2_out),
      .d1_button_pio_s1_end_xfer                                 (d1_button_pio_s1_end_xfer),
      .reset_n                                                   (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address_to_slave                (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_granted_button_pio_s1           (slow_peripheral_bridge_m1_granted_button_pio_s1),
      .slow_peripheral_bridge_m1_latency_counter                 (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_nativeaddress                   (slow_peripheral_bridge_m1_nativeaddress),
      .slow_peripheral_bridge_m1_qualified_request_button_pio_s1 (slow_peripheral_bridge_m1_qualified_request_button_pio_s1),
      .slow_peripheral_bridge_m1_read                            (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_button_pio_s1   (slow_peripheral_bridge_m1_read_data_valid_button_pio_s1),
      .slow_peripheral_bridge_m1_requests_button_pio_s1          (slow_peripheral_bridge_m1_requests_button_pio_s1),
      .slow_peripheral_bridge_m1_write                           (slow_peripheral_bridge_m1_write),
      .slow_peripheral_bridge_m1_writedata                       (slow_peripheral_bridge_m1_writedata)
    );

  button_pio the_button_pio
    (
      .address    (button_pio_s1_address),
      .chipselect (button_pio_s1_chipselect),
      .clk        (pll_c2_out),
      .in_port    (in_port_to_the_button_pio),
      .irq        (button_pio_s1_irq),
      .readdata   (button_pio_s1_readdata),
      .reset_n    (button_pio_s1_reset_n),
      .write_n    (button_pio_s1_write_n),
      .writedata  (button_pio_s1_writedata)
    );

  cpu_jtag_debug_module_arbitrator the_cpu_jtag_debug_module
    (
      .clk                                                                                             (pll_c0_out),
      .cpu_data_master_address_to_slave                                                                (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                                      (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                                                     (cpu_data_master_debugaccess),
      .cpu_data_master_granted_cpu_jtag_debug_module                                                   (cpu_data_master_granted_cpu_jtag_debug_module),
      .cpu_data_master_latency_counter                                                                 (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_cpu_jtag_debug_module                                         (cpu_data_master_qualified_request_cpu_jtag_debug_module),
      .cpu_data_master_read                                                                            (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                          (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_cpu_jtag_debug_module                                           (cpu_data_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register        (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register                        (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register),
      .cpu_data_master_requests_cpu_jtag_debug_module                                                  (cpu_data_master_requests_cpu_jtag_debug_module),
      .cpu_data_master_write                                                                           (cpu_data_master_write),
      .cpu_data_master_writedata                                                                       (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                                                         (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_cpu_jtag_debug_module                                            (cpu_instruction_master_granted_cpu_jtag_debug_module),
      .cpu_instruction_master_latency_counter                                                          (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_cpu_jtag_debug_module                                  (cpu_instruction_master_qualified_request_cpu_jtag_debug_module),
      .cpu_instruction_master_read                                                                     (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                   (cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_instruction_master_read_data_valid_cpu_jtag_debug_module                                    (cpu_instruction_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register (cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_instruction_master_requests_cpu_jtag_debug_module                                           (cpu_instruction_master_requests_cpu_jtag_debug_module),
      .cpu_jtag_debug_module_address                                                                   (cpu_jtag_debug_module_address),
      .cpu_jtag_debug_module_begintransfer                                                             (cpu_jtag_debug_module_begintransfer),
      .cpu_jtag_debug_module_byteenable                                                                (cpu_jtag_debug_module_byteenable),
      .cpu_jtag_debug_module_chipselect                                                                (cpu_jtag_debug_module_chipselect),
      .cpu_jtag_debug_module_debugaccess                                                               (cpu_jtag_debug_module_debugaccess),
      .cpu_jtag_debug_module_readdata                                                                  (cpu_jtag_debug_module_readdata),
      .cpu_jtag_debug_module_readdata_from_sa                                                          (cpu_jtag_debug_module_readdata_from_sa),
      .cpu_jtag_debug_module_reset_n                                                                   (cpu_jtag_debug_module_reset_n),
      .cpu_jtag_debug_module_resetrequest                                                              (cpu_jtag_debug_module_resetrequest),
      .cpu_jtag_debug_module_resetrequest_from_sa                                                      (cpu_jtag_debug_module_resetrequest_from_sa),
      .cpu_jtag_debug_module_write                                                                     (cpu_jtag_debug_module_write),
      .cpu_jtag_debug_module_writedata                                                                 (cpu_jtag_debug_module_writedata),
      .d1_cpu_jtag_debug_module_end_xfer                                                               (d1_cpu_jtag_debug_module_end_xfer),
      .reset_n                                                                                         (pll_c0_out_reset_n)
    );

  cpu_data_master_arbitrator the_cpu_data_master
    (
      .button_pio_s1_irq_from_sa                                                                (button_pio_s1_irq_from_sa),
      .clk                                                                                      (pll_c0_out),
      .cpu_data_master_address                                                                  (cpu_data_master_address),
      .cpu_data_master_address_to_slave                                                         (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                               (cpu_data_master_byteenable),
      .cpu_data_master_granted_cpu_ddr_clock_bridge_s1                                          (cpu_data_master_granted_cpu_ddr_clock_bridge_s1),
      .cpu_data_master_granted_cpu_jtag_debug_module                                            (cpu_data_master_granted_cpu_jtag_debug_module),
      .cpu_data_master_granted_descriptor_memory_s1                                             (cpu_data_master_granted_descriptor_memory_s1),
      .cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1                        (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_data_master_granted_sgdma_rx_csr                                                     (cpu_data_master_granted_sgdma_rx_csr),
      .cpu_data_master_granted_sgdma_tx_csr                                                     (cpu_data_master_granted_sgdma_tx_csr),
      .cpu_data_master_granted_slow_peripheral_bridge_s1                                        (cpu_data_master_granted_slow_peripheral_bridge_s1),
      .cpu_data_master_granted_tse_mac_control_port                                             (cpu_data_master_granted_tse_mac_control_port),
      .cpu_data_master_irq                                                                      (cpu_data_master_irq),
      .cpu_data_master_latency_counter                                                          (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1                                (cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1),
      .cpu_data_master_qualified_request_cpu_jtag_debug_module                                  (cpu_data_master_qualified_request_cpu_jtag_debug_module),
      .cpu_data_master_qualified_request_descriptor_memory_s1                                   (cpu_data_master_qualified_request_descriptor_memory_s1),
      .cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1              (cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_data_master_qualified_request_sgdma_rx_csr                                           (cpu_data_master_qualified_request_sgdma_rx_csr),
      .cpu_data_master_qualified_request_sgdma_tx_csr                                           (cpu_data_master_qualified_request_sgdma_tx_csr),
      .cpu_data_master_qualified_request_slow_peripheral_bridge_s1                              (cpu_data_master_qualified_request_slow_peripheral_bridge_s1),
      .cpu_data_master_qualified_request_tse_mac_control_port                                   (cpu_data_master_qualified_request_tse_mac_control_port),
      .cpu_data_master_read                                                                     (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1                                  (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                   (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_cpu_jtag_debug_module                                    (cpu_data_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_data_master_read_data_valid_descriptor_memory_s1                                     (cpu_data_master_read_data_valid_descriptor_memory_s1),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1                (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_sgdma_rx_csr                                             (cpu_data_master_read_data_valid_sgdma_rx_csr),
      .cpu_data_master_read_data_valid_sgdma_tx_csr                                             (cpu_data_master_read_data_valid_sgdma_tx_csr),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1                                (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register                 (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_tse_mac_control_port                                     (cpu_data_master_read_data_valid_tse_mac_control_port),
      .cpu_data_master_readdata                                                                 (cpu_data_master_readdata),
      .cpu_data_master_readdatavalid                                                            (cpu_data_master_readdatavalid),
      .cpu_data_master_requests_cpu_ddr_clock_bridge_s1                                         (cpu_data_master_requests_cpu_ddr_clock_bridge_s1),
      .cpu_data_master_requests_cpu_jtag_debug_module                                           (cpu_data_master_requests_cpu_jtag_debug_module),
      .cpu_data_master_requests_descriptor_memory_s1                                            (cpu_data_master_requests_descriptor_memory_s1),
      .cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1                       (cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_data_master_requests_sgdma_rx_csr                                                    (cpu_data_master_requests_sgdma_rx_csr),
      .cpu_data_master_requests_sgdma_tx_csr                                                    (cpu_data_master_requests_sgdma_tx_csr),
      .cpu_data_master_requests_slow_peripheral_bridge_s1                                       (cpu_data_master_requests_slow_peripheral_bridge_s1),
      .cpu_data_master_requests_tse_mac_control_port                                            (cpu_data_master_requests_tse_mac_control_port),
      .cpu_data_master_waitrequest                                                              (cpu_data_master_waitrequest),
      .cpu_data_master_write                                                                    (cpu_data_master_write),
      .cpu_data_master_writedata                                                                (cpu_data_master_writedata),
      .cpu_ddr_clock_bridge_s1_readdata_from_sa                                                 (cpu_ddr_clock_bridge_s1_readdata_from_sa),
      .cpu_ddr_clock_bridge_s1_waitrequest_from_sa                                              (cpu_ddr_clock_bridge_s1_waitrequest_from_sa),
      .cpu_jtag_debug_module_readdata_from_sa                                                   (cpu_jtag_debug_module_readdata_from_sa),
      .d1_cpu_ddr_clock_bridge_s1_end_xfer                                                      (d1_cpu_ddr_clock_bridge_s1_end_xfer),
      .d1_cpu_jtag_debug_module_end_xfer                                                        (d1_cpu_jtag_debug_module_end_xfer),
      .d1_descriptor_memory_s1_end_xfer                                                         (d1_descriptor_memory_s1_end_xfer),
      .d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer                                    (d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer),
      .d1_sgdma_rx_csr_end_xfer                                                                 (d1_sgdma_rx_csr_end_xfer),
      .d1_sgdma_tx_csr_end_xfer                                                                 (d1_sgdma_tx_csr_end_xfer),
      .d1_slow_peripheral_bridge_s1_end_xfer                                                    (d1_slow_peripheral_bridge_s1_end_xfer),
      .d1_tse_mac_control_port_end_xfer                                                         (d1_tse_mac_control_port_end_xfer),
      .descriptor_memory_s1_readdata_from_sa                                                    (descriptor_memory_s1_readdata_from_sa),
      .high_res_timer_s1_irq_from_sa                                                            (high_res_timer_s1_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                                                  (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa                               (pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa),
      .pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa                            (pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa),
      .pll_c0_out                                                                               (pll_c0_out),
      .pll_c0_out_reset_n                                                                       (pll_c0_out_reset_n),
      .reset_n                                                                                  (pll_c0_out_reset_n),
      .sgdma_rx_csr_irq_from_sa                                                                 (sgdma_rx_csr_irq_from_sa),
      .sgdma_rx_csr_readdata_from_sa                                                            (sgdma_rx_csr_readdata_from_sa),
      .sgdma_tx_csr_irq_from_sa                                                                 (sgdma_tx_csr_irq_from_sa),
      .sgdma_tx_csr_readdata_from_sa                                                            (sgdma_tx_csr_readdata_from_sa),
      .slow_peripheral_bridge_s1_readdata_from_sa                                               (slow_peripheral_bridge_s1_readdata_from_sa),
      .slow_peripheral_bridge_s1_waitrequest_from_sa                                            (slow_peripheral_bridge_s1_waitrequest_from_sa),
      .sys_clk_timer_s1_irq_from_sa                                                             (sys_clk_timer_s1_irq_from_sa),
      .tse_mac_control_port_readdata_from_sa                                                    (tse_mac_control_port_readdata_from_sa),
      .tse_mac_control_port_waitrequest_from_sa                                                 (tse_mac_control_port_waitrequest_from_sa)
    );

  cpu_instruction_master_arbitrator the_cpu_instruction_master
    (
      .clk                                                                                             (pll_c0_out),
      .cpu_ddr_clock_bridge_s1_readdata_from_sa                                                        (cpu_ddr_clock_bridge_s1_readdata_from_sa),
      .cpu_ddr_clock_bridge_s1_waitrequest_from_sa                                                     (cpu_ddr_clock_bridge_s1_waitrequest_from_sa),
      .cpu_instruction_master_address                                                                  (cpu_instruction_master_address),
      .cpu_instruction_master_address_to_slave                                                         (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1                                          (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1),
      .cpu_instruction_master_granted_cpu_jtag_debug_module                                            (cpu_instruction_master_granted_cpu_jtag_debug_module),
      .cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1                        (cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_instruction_master_latency_counter                                                          (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1                                (cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1),
      .cpu_instruction_master_qualified_request_cpu_jtag_debug_module                                  (cpu_instruction_master_qualified_request_cpu_jtag_debug_module),
      .cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1              (cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_instruction_master_read                                                                     (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1                                  (cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1),
      .cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                   (cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_instruction_master_read_data_valid_cpu_jtag_debug_module                                    (cpu_instruction_master_read_data_valid_cpu_jtag_debug_module),
      .cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1                (cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register (cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_instruction_master_readdata                                                                 (cpu_instruction_master_readdata),
      .cpu_instruction_master_readdatavalid                                                            (cpu_instruction_master_readdatavalid),
      .cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1                                         (cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1),
      .cpu_instruction_master_requests_cpu_jtag_debug_module                                           (cpu_instruction_master_requests_cpu_jtag_debug_module),
      .cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1                       (cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_instruction_master_waitrequest                                                              (cpu_instruction_master_waitrequest),
      .cpu_jtag_debug_module_readdata_from_sa                                                          (cpu_jtag_debug_module_readdata_from_sa),
      .d1_cpu_ddr_clock_bridge_s1_end_xfer                                                             (d1_cpu_ddr_clock_bridge_s1_end_xfer),
      .d1_cpu_jtag_debug_module_end_xfer                                                               (d1_cpu_jtag_debug_module_end_xfer),
      .d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer                                           (d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer),
      .pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa                                      (pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa),
      .pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa                                   (pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa),
      .reset_n                                                                                         (pll_c0_out_reset_n)
    );

  cpu the_cpu
    (
      .clk                                   (pll_c0_out),
      .d_address                             (cpu_data_master_address),
      .d_byteenable                          (cpu_data_master_byteenable),
      .d_irq                                 (cpu_data_master_irq),
      .d_read                                (cpu_data_master_read),
      .d_readdata                            (cpu_data_master_readdata),
      .d_readdatavalid                       (cpu_data_master_readdatavalid),
      .d_waitrequest                         (cpu_data_master_waitrequest),
      .d_write                               (cpu_data_master_write),
      .d_writedata                           (cpu_data_master_writedata),
      .i_address                             (cpu_instruction_master_address),
      .i_read                                (cpu_instruction_master_read),
      .i_readdata                            (cpu_instruction_master_readdata),
      .i_readdatavalid                       (cpu_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_jtag_debug_module_writedata),
      .reset_n                               (cpu_jtag_debug_module_reset_n)
    );

  cpu_ddr_clock_bridge_s1_arbitrator the_cpu_ddr_clock_bridge_s1
    (
      .clk                                                                                             (pll_c0_out),
      .cpu_data_master_address_to_slave                                                                (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                                      (cpu_data_master_byteenable),
      .cpu_data_master_granted_cpu_ddr_clock_bridge_s1                                                 (cpu_data_master_granted_cpu_ddr_clock_bridge_s1),
      .cpu_data_master_latency_counter                                                                 (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1                                       (cpu_data_master_qualified_request_cpu_ddr_clock_bridge_s1),
      .cpu_data_master_read                                                                            (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1                                         (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                          (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register        (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register                        (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register),
      .cpu_data_master_requests_cpu_ddr_clock_bridge_s1                                                (cpu_data_master_requests_cpu_ddr_clock_bridge_s1),
      .cpu_data_master_write                                                                           (cpu_data_master_write),
      .cpu_data_master_writedata                                                                       (cpu_data_master_writedata),
      .cpu_ddr_clock_bridge_s1_address                                                                 (cpu_ddr_clock_bridge_s1_address),
      .cpu_ddr_clock_bridge_s1_byteenable                                                              (cpu_ddr_clock_bridge_s1_byteenable),
      .cpu_ddr_clock_bridge_s1_endofpacket                                                             (cpu_ddr_clock_bridge_s1_endofpacket),
      .cpu_ddr_clock_bridge_s1_endofpacket_from_sa                                                     (cpu_ddr_clock_bridge_s1_endofpacket_from_sa),
      .cpu_ddr_clock_bridge_s1_nativeaddress                                                           (cpu_ddr_clock_bridge_s1_nativeaddress),
      .cpu_ddr_clock_bridge_s1_read                                                                    (cpu_ddr_clock_bridge_s1_read),
      .cpu_ddr_clock_bridge_s1_readdata                                                                (cpu_ddr_clock_bridge_s1_readdata),
      .cpu_ddr_clock_bridge_s1_readdata_from_sa                                                        (cpu_ddr_clock_bridge_s1_readdata_from_sa),
      .cpu_ddr_clock_bridge_s1_readdatavalid                                                           (cpu_ddr_clock_bridge_s1_readdatavalid),
      .cpu_ddr_clock_bridge_s1_reset_n                                                                 (cpu_ddr_clock_bridge_s1_reset_n),
      .cpu_ddr_clock_bridge_s1_waitrequest                                                             (cpu_ddr_clock_bridge_s1_waitrequest),
      .cpu_ddr_clock_bridge_s1_waitrequest_from_sa                                                     (cpu_ddr_clock_bridge_s1_waitrequest_from_sa),
      .cpu_ddr_clock_bridge_s1_write                                                                   (cpu_ddr_clock_bridge_s1_write),
      .cpu_ddr_clock_bridge_s1_writedata                                                               (cpu_ddr_clock_bridge_s1_writedata),
      .cpu_instruction_master_address_to_slave                                                         (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1                                          (cpu_instruction_master_granted_cpu_ddr_clock_bridge_s1),
      .cpu_instruction_master_latency_counter                                                          (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1                                (cpu_instruction_master_qualified_request_cpu_ddr_clock_bridge_s1),
      .cpu_instruction_master_read                                                                     (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1                                  (cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1),
      .cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                   (cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register (cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1                                         (cpu_instruction_master_requests_cpu_ddr_clock_bridge_s1),
      .d1_cpu_ddr_clock_bridge_s1_end_xfer                                                             (d1_cpu_ddr_clock_bridge_s1_end_xfer),
      .reset_n                                                                                         (pll_c0_out_reset_n),
      .sgdma_rx_m_write_address_to_slave                                                               (sgdma_rx_m_write_address_to_slave),
      .sgdma_rx_m_write_byteenable                                                                     (sgdma_rx_m_write_byteenable),
      .sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1                                                (sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1),
      .sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1                                      (sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1),
      .sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1                                               (sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1),
      .sgdma_rx_m_write_write                                                                          (sgdma_rx_m_write_write),
      .sgdma_rx_m_write_writedata                                                                      (sgdma_rx_m_write_writedata),
      .sgdma_tx_m_read_address_to_slave                                                                (sgdma_tx_m_read_address_to_slave),
      .sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1                                                 (sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1),
      .sgdma_tx_m_read_latency_counter                                                                 (sgdma_tx_m_read_latency_counter),
      .sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1                                       (sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1),
      .sgdma_tx_m_read_read                                                                            (sgdma_tx_m_read_read),
      .sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1                                         (sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1),
      .sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                          (sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1                                                (sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1)
    );

  cpu_ddr_clock_bridge_m1_arbitrator the_cpu_ddr_clock_bridge_m1
    (
      .clk                                                                  (ddr2_sdram_phy_clk_out),
      .cpu_ddr_clock_bridge_m1_address                                      (cpu_ddr_clock_bridge_m1_address),
      .cpu_ddr_clock_bridge_m1_address_to_slave                             (cpu_ddr_clock_bridge_m1_address_to_slave),
      .cpu_ddr_clock_bridge_m1_byteenable                                   (cpu_ddr_clock_bridge_m1_byteenable),
      .cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1                        (cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1),
      .cpu_ddr_clock_bridge_m1_latency_counter                              (cpu_ddr_clock_bridge_m1_latency_counter),
      .cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1              (cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1),
      .cpu_ddr_clock_bridge_m1_read                                         (cpu_ddr_clock_bridge_m1_read),
      .cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1                (cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1),
      .cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register (cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register),
      .cpu_ddr_clock_bridge_m1_readdata                                     (cpu_ddr_clock_bridge_m1_readdata),
      .cpu_ddr_clock_bridge_m1_readdatavalid                                (cpu_ddr_clock_bridge_m1_readdatavalid),
      .cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1                       (cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1),
      .cpu_ddr_clock_bridge_m1_reset_n                                      (cpu_ddr_clock_bridge_m1_reset_n),
      .cpu_ddr_clock_bridge_m1_waitrequest                                  (cpu_ddr_clock_bridge_m1_waitrequest),
      .cpu_ddr_clock_bridge_m1_write                                        (cpu_ddr_clock_bridge_m1_write),
      .cpu_ddr_clock_bridge_m1_writedata                                    (cpu_ddr_clock_bridge_m1_writedata),
      .d1_ddr2_sdram_s1_end_xfer                                            (d1_ddr2_sdram_s1_end_xfer),
      .ddr2_sdram_s1_readdata_from_sa                                       (ddr2_sdram_s1_readdata_from_sa),
      .ddr2_sdram_s1_waitrequest_n_from_sa                                  (ddr2_sdram_s1_waitrequest_n_from_sa),
      .reset_n                                                              (ddr2_sdram_phy_clk_out_reset_n)
    );

  cpu_ddr_clock_bridge the_cpu_ddr_clock_bridge
    (
      .master_address       (cpu_ddr_clock_bridge_m1_address),
      .master_byteenable    (cpu_ddr_clock_bridge_m1_byteenable),
      .master_clk           (ddr2_sdram_phy_clk_out),
      .master_endofpacket   (cpu_ddr_clock_bridge_m1_endofpacket),
      .master_nativeaddress (cpu_ddr_clock_bridge_m1_nativeaddress),
      .master_read          (cpu_ddr_clock_bridge_m1_read),
      .master_readdata      (cpu_ddr_clock_bridge_m1_readdata),
      .master_readdatavalid (cpu_ddr_clock_bridge_m1_readdatavalid),
      .master_reset_n       (cpu_ddr_clock_bridge_m1_reset_n),
      .master_waitrequest   (cpu_ddr_clock_bridge_m1_waitrequest),
      .master_write         (cpu_ddr_clock_bridge_m1_write),
      .master_writedata     (cpu_ddr_clock_bridge_m1_writedata),
      .slave_address        (cpu_ddr_clock_bridge_s1_address),
      .slave_byteenable     (cpu_ddr_clock_bridge_s1_byteenable),
      .slave_clk            (pll_c0_out),
      .slave_endofpacket    (cpu_ddr_clock_bridge_s1_endofpacket),
      .slave_nativeaddress  (cpu_ddr_clock_bridge_s1_nativeaddress),
      .slave_read           (cpu_ddr_clock_bridge_s1_read),
      .slave_readdata       (cpu_ddr_clock_bridge_s1_readdata),
      .slave_readdatavalid  (cpu_ddr_clock_bridge_s1_readdatavalid),
      .slave_reset_n        (cpu_ddr_clock_bridge_s1_reset_n),
      .slave_waitrequest    (cpu_ddr_clock_bridge_s1_waitrequest),
      .slave_write          (cpu_ddr_clock_bridge_s1_write),
      .slave_writedata      (cpu_ddr_clock_bridge_s1_writedata)
    );

  cycloneIII_3c120_niosII_standard_sopc_clock_0_in_arbitrator the_cycloneIII_3c120_niosII_standard_sopc_clock_0_in
    (
      .clk                                                                                          (pll_c2_out),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_address                                     (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_address),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_byteenable                                  (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_byteenable),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket                                 (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_nativeaddress                               (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_nativeaddress),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_read                                        (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_read),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata                                    (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa                            (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reset_n                                     (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reset_n),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest                                 (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_write                                       (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_write),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_writedata                                   (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_writedata),
      .d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer                                 (d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer),
      .reset_n                                                                                      (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address_to_slave                                                   (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_byteenable                                                         (slow_peripheral_bridge_m1_byteenable),
      .slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in           (slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in),
      .slow_peripheral_bridge_m1_latency_counter                                                    (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_nativeaddress                                                      (slow_peripheral_bridge_m1_nativeaddress),
      .slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in (slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in),
      .slow_peripheral_bridge_m1_read                                                               (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in   (slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in),
      .slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in          (slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in),
      .slow_peripheral_bridge_m1_write                                                              (slow_peripheral_bridge_m1_write),
      .slow_peripheral_bridge_m1_writedata                                                          (slow_peripheral_bridge_m1_writedata)
    );

  cycloneIII_3c120_niosII_standard_sopc_clock_0_out_arbitrator the_cycloneIII_3c120_niosII_standard_sopc_clock_0_out
    (
      .clk                                                                        (clk),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address                  (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave         (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable               (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1           (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1 (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read                     (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_data_valid_pll_s1   (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_data_valid_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_readdata                 (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_readdata),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1          (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_reset_n                  (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_reset_n),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_waitrequest              (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_waitrequest),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write                    (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata                (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata),
      .d1_pll_s1_end_xfer                                                         (d1_pll_s1_end_xfer),
      .pll_s1_readdata_from_sa                                                    (pll_s1_readdata_from_sa),
      .reset_n                                                                    (clk_reset_n)
    );

  cycloneIII_3c120_niosII_standard_sopc_clock_0 the_cycloneIII_3c120_niosII_standard_sopc_clock_0
    (
      .master_address       (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address),
      .master_byteenable    (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_byteenable),
      .master_clk           (clk),
      .master_endofpacket   (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_endofpacket),
      .master_nativeaddress (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_nativeaddress),
      .master_read          (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read),
      .master_readdata      (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_readdata),
      .master_reset_n       (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_reset_n),
      .master_waitrequest   (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_waitrequest),
      .master_write         (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write),
      .master_writedata     (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata),
      .slave_address        (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_address),
      .slave_byteenable     (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_byteenable),
      .slave_clk            (pll_c2_out),
      .slave_endofpacket    (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket),
      .slave_nativeaddress  (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_nativeaddress),
      .slave_read           (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_read),
      .slave_readdata       (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata),
      .slave_reset_n        (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_reset_n),
      .slave_waitrequest    (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest),
      .slave_write          (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_write),
      .slave_writedata      (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_writedata)
    );

  cycloneIII_3c120_niosII_standard_sopc_clock_1_in_arbitrator the_cycloneIII_3c120_niosII_standard_sopc_clock_1_in
    (
      .clk                                                                                          (pll_c2_out),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_address                                     (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_address),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_byteenable                                  (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_byteenable),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket                                 (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_nativeaddress                               (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_nativeaddress),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_read                                        (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_read),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata                                    (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa                            (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reset_n                                     (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reset_n),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest                                 (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_write                                       (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_write),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_writedata                                   (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_writedata),
      .d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer                                 (d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer),
      .reset_n                                                                                      (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address_to_slave                                                   (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_byteenable                                                         (slow_peripheral_bridge_m1_byteenable),
      .slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in           (slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in),
      .slow_peripheral_bridge_m1_latency_counter                                                    (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_nativeaddress                                                      (slow_peripheral_bridge_m1_nativeaddress),
      .slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in (slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in),
      .slow_peripheral_bridge_m1_read                                                               (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in   (slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in),
      .slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in          (slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in),
      .slow_peripheral_bridge_m1_write                                                              (slow_peripheral_bridge_m1_write),
      .slow_peripheral_bridge_m1_writedata                                                          (slow_peripheral_bridge_m1_writedata)
    );

  cycloneIII_3c120_niosII_standard_sopc_clock_1_out_arbitrator the_cycloneIII_3c120_niosII_standard_sopc_clock_1_out
    (
      .clk                                                                            (clk_to_tse_pll),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address                      (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave             (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable                   (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1           (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1 (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read                         (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_data_valid_tse_pll_s1   (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_data_valid_tse_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_readdata                     (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_readdata),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1          (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_reset_n                      (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_reset_n),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_waitrequest                  (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_waitrequest),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write                        (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata                    (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata),
      .d1_tse_pll_s1_end_xfer                                                         (d1_tse_pll_s1_end_xfer),
      .reset_n                                                                        (clk_to_tse_pll_reset_n),
      .tse_pll_s1_readdata_from_sa                                                    (tse_pll_s1_readdata_from_sa)
    );

  cycloneIII_3c120_niosII_standard_sopc_clock_1 the_cycloneIII_3c120_niosII_standard_sopc_clock_1
    (
      .master_address       (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address),
      .master_byteenable    (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_byteenable),
      .master_clk           (clk_to_tse_pll),
      .master_endofpacket   (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_endofpacket),
      .master_nativeaddress (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_nativeaddress),
      .master_read          (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read),
      .master_readdata      (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_readdata),
      .master_reset_n       (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_reset_n),
      .master_waitrequest   (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_waitrequest),
      .master_write         (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write),
      .master_writedata     (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata),
      .slave_address        (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_address),
      .slave_byteenable     (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_byteenable),
      .slave_clk            (pll_c2_out),
      .slave_endofpacket    (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket),
      .slave_nativeaddress  (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_nativeaddress),
      .slave_read           (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_read),
      .slave_readdata       (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata),
      .slave_reset_n        (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_reset_n),
      .slave_waitrequest    (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest),
      .slave_write          (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_write),
      .slave_writedata      (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_writedata)
    );

  cycloneIII_3c120_niosII_standard_sopc_clock_2_in_arbitrator the_cycloneIII_3c120_niosII_standard_sopc_clock_2_in
    (
      .clk                                                                                          (pll_c2_out),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_address                                     (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_address),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_byteenable                                  (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_byteenable),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket                                 (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_nativeaddress                               (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_nativeaddress),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_read                                        (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_read),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata                                    (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa                            (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reset_n                                     (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reset_n),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest                                 (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_write                                       (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_write),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_writedata                                   (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_writedata),
      .d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer                                 (d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer),
      .reset_n                                                                                      (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address_to_slave                                                   (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_byteenable                                                         (slow_peripheral_bridge_m1_byteenable),
      .slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in           (slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in),
      .slow_peripheral_bridge_m1_latency_counter                                                    (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_nativeaddress                                                      (slow_peripheral_bridge_m1_nativeaddress),
      .slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in (slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in),
      .slow_peripheral_bridge_m1_read                                                               (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in   (slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in),
      .slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in          (slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in),
      .slow_peripheral_bridge_m1_write                                                              (slow_peripheral_bridge_m1_write),
      .slow_peripheral_bridge_m1_writedata                                                          (slow_peripheral_bridge_m1_writedata)
    );

  cycloneIII_3c120_niosII_standard_sopc_clock_2_out_arbitrator the_cycloneIII_3c120_niosII_standard_sopc_clock_2_out
    (
      .clk                                                                               (clk),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address                         (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave                (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable                      (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1           (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1 (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read                            (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_data_valid_tse_tx_pll_s1   (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_data_valid_tse_tx_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_readdata                        (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_readdata),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1          (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_reset_n                         (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_reset_n),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_waitrequest                     (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_waitrequest),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write                           (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata                       (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata),
      .d1_tse_tx_pll_s1_end_xfer                                                         (d1_tse_tx_pll_s1_end_xfer),
      .reset_n                                                                           (clk_reset_n),
      .tse_tx_pll_s1_readdata_from_sa                                                    (tse_tx_pll_s1_readdata_from_sa)
    );

  cycloneIII_3c120_niosII_standard_sopc_clock_2 the_cycloneIII_3c120_niosII_standard_sopc_clock_2
    (
      .master_address       (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address),
      .master_byteenable    (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_byteenable),
      .master_clk           (clk),
      .master_endofpacket   (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_endofpacket),
      .master_nativeaddress (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_nativeaddress),
      .master_read          (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read),
      .master_readdata      (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_readdata),
      .master_reset_n       (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_reset_n),
      .master_waitrequest   (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_waitrequest),
      .master_write         (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write),
      .master_writedata     (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata),
      .slave_address        (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_address),
      .slave_byteenable     (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_byteenable),
      .slave_clk            (pll_c2_out),
      .slave_endofpacket    (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket),
      .slave_nativeaddress  (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_nativeaddress),
      .slave_read           (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_read),
      .slave_readdata       (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata),
      .slave_reset_n        (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_reset_n),
      .slave_waitrequest    (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest),
      .slave_write          (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_write),
      .slave_writedata      (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_writedata)
    );

  ddr2_sdram_s1_arbitrator the_ddr2_sdram_s1
    (
      .clk                                                                  (ddr2_sdram_phy_clk_out),
      .cpu_ddr_clock_bridge_m1_address_to_slave                             (cpu_ddr_clock_bridge_m1_address_to_slave),
      .cpu_ddr_clock_bridge_m1_byteenable                                   (cpu_ddr_clock_bridge_m1_byteenable),
      .cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1                        (cpu_ddr_clock_bridge_m1_granted_ddr2_sdram_s1),
      .cpu_ddr_clock_bridge_m1_latency_counter                              (cpu_ddr_clock_bridge_m1_latency_counter),
      .cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1              (cpu_ddr_clock_bridge_m1_qualified_request_ddr2_sdram_s1),
      .cpu_ddr_clock_bridge_m1_read                                         (cpu_ddr_clock_bridge_m1_read),
      .cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1                (cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1),
      .cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register (cpu_ddr_clock_bridge_m1_read_data_valid_ddr2_sdram_s1_shift_register),
      .cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1                       (cpu_ddr_clock_bridge_m1_requests_ddr2_sdram_s1),
      .cpu_ddr_clock_bridge_m1_write                                        (cpu_ddr_clock_bridge_m1_write),
      .cpu_ddr_clock_bridge_m1_writedata                                    (cpu_ddr_clock_bridge_m1_writedata),
      .d1_ddr2_sdram_s1_end_xfer                                            (d1_ddr2_sdram_s1_end_xfer),
      .ddr2_sdram_s1_address                                                (ddr2_sdram_s1_address),
      .ddr2_sdram_s1_beginbursttransfer                                     (ddr2_sdram_s1_beginbursttransfer),
      .ddr2_sdram_s1_burstcount                                             (ddr2_sdram_s1_burstcount),
      .ddr2_sdram_s1_byteenable                                             (ddr2_sdram_s1_byteenable),
      .ddr2_sdram_s1_read                                                   (ddr2_sdram_s1_read),
      .ddr2_sdram_s1_readdata                                               (ddr2_sdram_s1_readdata),
      .ddr2_sdram_s1_readdata_from_sa                                       (ddr2_sdram_s1_readdata_from_sa),
      .ddr2_sdram_s1_readdatavalid                                          (ddr2_sdram_s1_readdatavalid),
      .ddr2_sdram_s1_resetrequest_n                                         (ddr2_sdram_s1_resetrequest_n),
      .ddr2_sdram_s1_resetrequest_n_from_sa                                 (ddr2_sdram_s1_resetrequest_n_from_sa),
      .ddr2_sdram_s1_waitrequest_n                                          (ddr2_sdram_s1_waitrequest_n),
      .ddr2_sdram_s1_waitrequest_n_from_sa                                  (ddr2_sdram_s1_waitrequest_n_from_sa),
      .ddr2_sdram_s1_write                                                  (ddr2_sdram_s1_write),
      .ddr2_sdram_s1_writedata                                              (ddr2_sdram_s1_writedata),
      .reset_n                                                              (ddr2_sdram_phy_clk_out_reset_n)
    );

  //ddr2_sdram_aux_full_rate_clk_out out_clk assignment, which is an e_assign
  assign ddr2_sdram_aux_full_rate_clk_out = out_clk_ddr2_sdram_aux_full_rate_clk;

  //ddr2_sdram_aux_half_rate_clk_out out_clk assignment, which is an e_assign
  assign ddr2_sdram_aux_half_rate_clk_out = out_clk_ddr2_sdram_aux_half_rate_clk;

  //ddr2_sdram_phy_clk_out out_clk assignment, which is an e_assign
  assign ddr2_sdram_phy_clk_out = out_clk_ddr2_sdram_phy_clk;

  //reset is asserted asynchronously and deasserted synchronously
  cycloneIII_3c120_niosII_standard_sopc_reset_clk_125_domain_synch_module cycloneIII_3c120_niosII_standard_sopc_reset_clk_125_domain_synch
    (
      .clk      (clk_125),
      .data_in  (1'b1),
      .data_out (clk_125_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset sources mux, which is an e_mux
  assign reset_n_sources = ~(~reset_n |
    0 |
    0 |
    0 |
    cpu_jtag_debug_module_resetrequest_from_sa |
    cpu_jtag_debug_module_resetrequest_from_sa |
    0 |
    ~ddr2_sdram_s1_resetrequest_n_from_sa |
    ~ddr2_sdram_s1_resetrequest_n_from_sa |
    0 |
    pll_s1_resetrequest_from_sa |
    pll_s1_resetrequest_from_sa |
    0 |
    tse_pll_s1_resetrequest_from_sa |
    tse_pll_s1_resetrequest_from_sa |
    tse_tx_pll_s1_resetrequest_from_sa |
    tse_tx_pll_s1_resetrequest_from_sa);

  ddr2_sdram the_ddr2_sdram
    (
      .aux_full_rate_clk (out_clk_ddr2_sdram_aux_full_rate_clk),
      .aux_half_rate_clk (out_clk_ddr2_sdram_aux_half_rate_clk),
      .global_reset_n    (global_reset_n_to_the_ddr2_sdram),
      .local_address     (ddr2_sdram_s1_address),
      .local_be          (ddr2_sdram_s1_byteenable),
      .local_burstbegin  (ddr2_sdram_s1_beginbursttransfer),
      .local_init_done   (local_init_done_from_the_ddr2_sdram),
      .local_rdata       (ddr2_sdram_s1_readdata),
      .local_rdata_valid (ddr2_sdram_s1_readdatavalid),
      .local_read_req    (ddr2_sdram_s1_read),
      .local_ready       (ddr2_sdram_s1_waitrequest_n),
      .local_refresh_ack (local_refresh_ack_from_the_ddr2_sdram),
      .local_size        (ddr2_sdram_s1_burstcount),
      .local_wdata       (ddr2_sdram_s1_writedata),
      .local_wdata_req   (local_wdata_req_from_the_ddr2_sdram),
      .local_write_req   (ddr2_sdram_s1_write),
      .mem_addr          (mem_addr_from_the_ddr2_sdram),
      .mem_ba            (mem_ba_from_the_ddr2_sdram),
      .mem_cas_n         (mem_cas_n_from_the_ddr2_sdram),
      .mem_cke           (mem_cke_from_the_ddr2_sdram),
      .mem_clk           (mem_clk_to_and_from_the_ddr2_sdram),
      .mem_clk_n         (mem_clk_n_to_and_from_the_ddr2_sdram),
      .mem_cs_n          (mem_cs_n_from_the_ddr2_sdram),
      .mem_dm            (mem_dm_from_the_ddr2_sdram),
      .mem_dq            (mem_dq_to_and_from_the_ddr2_sdram),
      .mem_dqs           (mem_dqs_to_and_from_the_ddr2_sdram),
      .mem_odt           (mem_odt_from_the_ddr2_sdram),
      .mem_ras_n         (mem_ras_n_from_the_ddr2_sdram),
      .mem_we_n          (mem_we_n_from_the_ddr2_sdram),
      .phy_clk           (out_clk_ddr2_sdram_phy_clk),
      .pll_ref_clk       (clk_125),
      .reset_phy_clk_n   (reset_phy_clk_n_from_the_ddr2_sdram),
      .reset_request_n   (ddr2_sdram_s1_resetrequest_n),
      .soft_reset_n      (clk_125_reset_n)
    );

  descriptor_memory_s1_arbitrator the_descriptor_memory_s1
    (
      .clk                                                                                      (pll_c0_out),
      .cpu_data_master_address_to_slave                                                         (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                               (cpu_data_master_byteenable),
      .cpu_data_master_granted_descriptor_memory_s1                                             (cpu_data_master_granted_descriptor_memory_s1),
      .cpu_data_master_latency_counter                                                          (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_descriptor_memory_s1                                   (cpu_data_master_qualified_request_descriptor_memory_s1),
      .cpu_data_master_read                                                                     (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                   (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_descriptor_memory_s1                                     (cpu_data_master_read_data_valid_descriptor_memory_s1),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register                 (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register),
      .cpu_data_master_requests_descriptor_memory_s1                                            (cpu_data_master_requests_descriptor_memory_s1),
      .cpu_data_master_write                                                                    (cpu_data_master_write),
      .cpu_data_master_writedata                                                                (cpu_data_master_writedata),
      .d1_descriptor_memory_s1_end_xfer                                                         (d1_descriptor_memory_s1_end_xfer),
      .descriptor_memory_s1_address                                                             (descriptor_memory_s1_address),
      .descriptor_memory_s1_byteenable                                                          (descriptor_memory_s1_byteenable),
      .descriptor_memory_s1_chipselect                                                          (descriptor_memory_s1_chipselect),
      .descriptor_memory_s1_clken                                                               (descriptor_memory_s1_clken),
      .descriptor_memory_s1_readdata                                                            (descriptor_memory_s1_readdata),
      .descriptor_memory_s1_readdata_from_sa                                                    (descriptor_memory_s1_readdata_from_sa),
      .descriptor_memory_s1_reset                                                               (descriptor_memory_s1_reset),
      .descriptor_memory_s1_write                                                               (descriptor_memory_s1_write),
      .descriptor_memory_s1_writedata                                                           (descriptor_memory_s1_writedata),
      .reset_n                                                                                  (pll_c0_out_reset_n),
      .sgdma_rx_descriptor_read_address_to_slave                                                (sgdma_rx_descriptor_read_address_to_slave),
      .sgdma_rx_descriptor_read_granted_descriptor_memory_s1                                    (sgdma_rx_descriptor_read_granted_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_latency_counter                                                 (sgdma_rx_descriptor_read_latency_counter),
      .sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1                          (sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_read                                                            (sgdma_rx_descriptor_read_read),
      .sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1                            (sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_requests_descriptor_memory_s1                                   (sgdma_rx_descriptor_read_requests_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_address_to_slave                                               (sgdma_rx_descriptor_write_address_to_slave),
      .sgdma_rx_descriptor_write_granted_descriptor_memory_s1                                   (sgdma_rx_descriptor_write_granted_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1                         (sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_requests_descriptor_memory_s1                                  (sgdma_rx_descriptor_write_requests_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_write                                                          (sgdma_rx_descriptor_write_write),
      .sgdma_rx_descriptor_write_writedata                                                      (sgdma_rx_descriptor_write_writedata),
      .sgdma_tx_descriptor_read_address_to_slave                                                (sgdma_tx_descriptor_read_address_to_slave),
      .sgdma_tx_descriptor_read_granted_descriptor_memory_s1                                    (sgdma_tx_descriptor_read_granted_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_latency_counter                                                 (sgdma_tx_descriptor_read_latency_counter),
      .sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1                          (sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_read                                                            (sgdma_tx_descriptor_read_read),
      .sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1                            (sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_requests_descriptor_memory_s1                                   (sgdma_tx_descriptor_read_requests_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_address_to_slave                                               (sgdma_tx_descriptor_write_address_to_slave),
      .sgdma_tx_descriptor_write_granted_descriptor_memory_s1                                   (sgdma_tx_descriptor_write_granted_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1                         (sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_requests_descriptor_memory_s1                                  (sgdma_tx_descriptor_write_requests_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_write                                                          (sgdma_tx_descriptor_write_write),
      .sgdma_tx_descriptor_write_writedata                                                      (sgdma_tx_descriptor_write_writedata)
    );

  descriptor_memory the_descriptor_memory
    (
      .address    (descriptor_memory_s1_address),
      .byteenable (descriptor_memory_s1_byteenable),
      .chipselect (descriptor_memory_s1_chipselect),
      .clk        (pll_c0_out),
      .clken      (descriptor_memory_s1_clken),
      .readdata   (descriptor_memory_s1_readdata),
      .reset      (descriptor_memory_s1_reset),
      .write      (descriptor_memory_s1_write),
      .writedata  (descriptor_memory_s1_writedata)
    );

  flash_tristate_bridge_avalon_slave_arbitrator the_flash_tristate_bridge_avalon_slave
    (
      .clk                                                                      (pll_c0_out),
      .cs_n_to_the_max2                                                         (cs_n_to_the_max2),
      .d1_flash_tristate_bridge_avalon_slave_end_xfer                           (d1_flash_tristate_bridge_avalon_slave_end_xfer),
      .ext_flash_s1_wait_counter_eq_0                                           (ext_flash_s1_wait_counter_eq_0),
      .flash_tristate_bridge_address                                            (flash_tristate_bridge_address),
      .flash_tristate_bridge_data                                               (flash_tristate_bridge_data),
      .incoming_flash_tristate_bridge_data                                      (incoming_flash_tristate_bridge_data),
      .incoming_flash_tristate_bridge_data_with_Xs_converted_to_0               (incoming_flash_tristate_bridge_data_with_Xs_converted_to_0),
      .max2_s1_wait_counter_eq_0                                                (max2_s1_wait_counter_eq_0),
      .oe_n_to_the_max2                                                         (oe_n_to_the_max2),
      .pipeline_bridge_before_tristate_bridge_m1_address_to_slave               (pipeline_bridge_before_tristate_bridge_m1_address_to_slave),
      .pipeline_bridge_before_tristate_bridge_m1_burstcount                     (pipeline_bridge_before_tristate_bridge_m1_burstcount),
      .pipeline_bridge_before_tristate_bridge_m1_byteenable                     (pipeline_bridge_before_tristate_bridge_m1_byteenable),
      .pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1        (pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1),
      .pipeline_bridge_before_tristate_bridge_m1_chipselect                     (pipeline_bridge_before_tristate_bridge_m1_chipselect),
      .pipeline_bridge_before_tristate_bridge_m1_dbs_address                    (pipeline_bridge_before_tristate_bridge_m1_dbs_address),
      .pipeline_bridge_before_tristate_bridge_m1_dbs_write_16                   (pipeline_bridge_before_tristate_bridge_m1_dbs_write_16),
      .pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1           (pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1),
      .pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1                (pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1),
      .pipeline_bridge_before_tristate_bridge_m1_latency_counter                (pipeline_bridge_before_tristate_bridge_m1_latency_counter),
      .pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1 (pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1),
      .pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1      (pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1),
      .pipeline_bridge_before_tristate_bridge_m1_read                           (pipeline_bridge_before_tristate_bridge_m1_read),
      .pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1   (pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1),
      .pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1        (pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1),
      .pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1          (pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1),
      .pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1               (pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1),
      .pipeline_bridge_before_tristate_bridge_m1_write                          (pipeline_bridge_before_tristate_bridge_m1_write),
      .pipeline_bridge_before_tristate_bridge_m1_writedata                      (pipeline_bridge_before_tristate_bridge_m1_writedata),
      .read_n_to_the_ext_flash                                                  (read_n_to_the_ext_flash),
      .reset_n                                                                  (pll_c0_out_reset_n),
      .select_n_to_the_ext_flash                                                (select_n_to_the_ext_flash),
      .we_n_to_the_max2                                                         (we_n_to_the_max2),
      .write_n_to_the_ext_flash                                                 (write_n_to_the_ext_flash)
    );

  high_res_timer_s1_arbitrator the_high_res_timer_s1
    (
      .clk                                                           (pll_c2_out),
      .d1_high_res_timer_s1_end_xfer                                 (d1_high_res_timer_s1_end_xfer),
      .high_res_timer_s1_address                                     (high_res_timer_s1_address),
      .high_res_timer_s1_chipselect                                  (high_res_timer_s1_chipselect),
      .high_res_timer_s1_irq                                         (high_res_timer_s1_irq),
      .high_res_timer_s1_irq_from_sa                                 (high_res_timer_s1_irq_from_sa),
      .high_res_timer_s1_readdata                                    (high_res_timer_s1_readdata),
      .high_res_timer_s1_readdata_from_sa                            (high_res_timer_s1_readdata_from_sa),
      .high_res_timer_s1_reset_n                                     (high_res_timer_s1_reset_n),
      .high_res_timer_s1_write_n                                     (high_res_timer_s1_write_n),
      .high_res_timer_s1_writedata                                   (high_res_timer_s1_writedata),
      .reset_n                                                       (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address_to_slave                    (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_granted_high_res_timer_s1           (slow_peripheral_bridge_m1_granted_high_res_timer_s1),
      .slow_peripheral_bridge_m1_latency_counter                     (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_nativeaddress                       (slow_peripheral_bridge_m1_nativeaddress),
      .slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1 (slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1),
      .slow_peripheral_bridge_m1_read                                (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1   (slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1),
      .slow_peripheral_bridge_m1_requests_high_res_timer_s1          (slow_peripheral_bridge_m1_requests_high_res_timer_s1),
      .slow_peripheral_bridge_m1_write                               (slow_peripheral_bridge_m1_write),
      .slow_peripheral_bridge_m1_writedata                           (slow_peripheral_bridge_m1_writedata)
    );

  high_res_timer the_high_res_timer
    (
      .address    (high_res_timer_s1_address),
      .chipselect (high_res_timer_s1_chipselect),
      .clk        (pll_c2_out),
      .irq        (high_res_timer_s1_irq),
      .readdata   (high_res_timer_s1_readdata),
      .reset_n    (high_res_timer_s1_reset_n),
      .write_n    (high_res_timer_s1_write_n),
      .writedata  (high_res_timer_s1_writedata)
    );

  jtag_uart_avalon_jtag_slave_arbitrator the_jtag_uart_avalon_jtag_slave
    (
      .clk                                                                     (pll_c2_out),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                                 (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .jtag_uart_avalon_jtag_slave_address                                     (jtag_uart_avalon_jtag_slave_address),
      .jtag_uart_avalon_jtag_slave_chipselect                                  (jtag_uart_avalon_jtag_slave_chipselect),
      .jtag_uart_avalon_jtag_slave_dataavailable                               (jtag_uart_avalon_jtag_slave_dataavailable),
      .jtag_uart_avalon_jtag_slave_dataavailable_from_sa                       (jtag_uart_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_avalon_jtag_slave_irq                                         (jtag_uart_avalon_jtag_slave_irq),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                                 (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_read_n                                      (jtag_uart_avalon_jtag_slave_read_n),
      .jtag_uart_avalon_jtag_slave_readdata                                    (jtag_uart_avalon_jtag_slave_readdata),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                            (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_readyfordata                                (jtag_uart_avalon_jtag_slave_readyfordata),
      .jtag_uart_avalon_jtag_slave_readyfordata_from_sa                        (jtag_uart_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_avalon_jtag_slave_reset_n                                     (jtag_uart_avalon_jtag_slave_reset_n),
      .jtag_uart_avalon_jtag_slave_waitrequest                                 (jtag_uart_avalon_jtag_slave_waitrequest),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa                         (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_avalon_jtag_slave_write_n                                     (jtag_uart_avalon_jtag_slave_write_n),
      .jtag_uart_avalon_jtag_slave_writedata                                   (jtag_uart_avalon_jtag_slave_writedata),
      .reset_n                                                                 (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address_to_slave                              (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave           (slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave),
      .slow_peripheral_bridge_m1_latency_counter                               (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_nativeaddress                                 (slow_peripheral_bridge_m1_nativeaddress),
      .slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave (slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave),
      .slow_peripheral_bridge_m1_read                                          (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave   (slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave),
      .slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave          (slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave),
      .slow_peripheral_bridge_m1_write                                         (slow_peripheral_bridge_m1_write),
      .slow_peripheral_bridge_m1_writedata                                     (slow_peripheral_bridge_m1_writedata)
    );

  jtag_uart the_jtag_uart
    (
      .av_address     (jtag_uart_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_avalon_jtag_slave_writedata),
      .clk            (pll_c2_out),
      .dataavailable  (jtag_uart_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_avalon_jtag_slave_reset_n)
    );

  led_pio_s1_arbitrator the_led_pio_s1
    (
      .clk                                                    (pll_c2_out),
      .d1_led_pio_s1_end_xfer                                 (d1_led_pio_s1_end_xfer),
      .led_pio_s1_address                                     (led_pio_s1_address),
      .led_pio_s1_chipselect                                  (led_pio_s1_chipselect),
      .led_pio_s1_readdata                                    (led_pio_s1_readdata),
      .led_pio_s1_readdata_from_sa                            (led_pio_s1_readdata_from_sa),
      .led_pio_s1_reset_n                                     (led_pio_s1_reset_n),
      .led_pio_s1_write_n                                     (led_pio_s1_write_n),
      .led_pio_s1_writedata                                   (led_pio_s1_writedata),
      .reset_n                                                (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address_to_slave             (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_granted_led_pio_s1           (slow_peripheral_bridge_m1_granted_led_pio_s1),
      .slow_peripheral_bridge_m1_latency_counter              (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_nativeaddress                (slow_peripheral_bridge_m1_nativeaddress),
      .slow_peripheral_bridge_m1_qualified_request_led_pio_s1 (slow_peripheral_bridge_m1_qualified_request_led_pio_s1),
      .slow_peripheral_bridge_m1_read                         (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_led_pio_s1   (slow_peripheral_bridge_m1_read_data_valid_led_pio_s1),
      .slow_peripheral_bridge_m1_requests_led_pio_s1          (slow_peripheral_bridge_m1_requests_led_pio_s1),
      .slow_peripheral_bridge_m1_write                        (slow_peripheral_bridge_m1_write),
      .slow_peripheral_bridge_m1_writedata                    (slow_peripheral_bridge_m1_writedata)
    );

  led_pio the_led_pio
    (
      .address    (led_pio_s1_address),
      .chipselect (led_pio_s1_chipselect),
      .clk        (pll_c2_out),
      .out_port   (out_port_from_the_led_pio),
      .readdata   (led_pio_s1_readdata),
      .reset_n    (led_pio_s1_reset_n),
      .write_n    (led_pio_s1_write_n),
      .writedata  (led_pio_s1_writedata)
    );

  performance_counter_control_slave_arbitrator the_performance_counter_control_slave
    (
      .clk                                                                           (pll_c2_out),
      .d1_performance_counter_control_slave_end_xfer                                 (d1_performance_counter_control_slave_end_xfer),
      .performance_counter_control_slave_address                                     (performance_counter_control_slave_address),
      .performance_counter_control_slave_begintransfer                               (performance_counter_control_slave_begintransfer),
      .performance_counter_control_slave_readdata                                    (performance_counter_control_slave_readdata),
      .performance_counter_control_slave_readdata_from_sa                            (performance_counter_control_slave_readdata_from_sa),
      .performance_counter_control_slave_reset_n                                     (performance_counter_control_slave_reset_n),
      .performance_counter_control_slave_write                                       (performance_counter_control_slave_write),
      .performance_counter_control_slave_writedata                                   (performance_counter_control_slave_writedata),
      .reset_n                                                                       (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address_to_slave                                    (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_granted_performance_counter_control_slave           (slow_peripheral_bridge_m1_granted_performance_counter_control_slave),
      .slow_peripheral_bridge_m1_latency_counter                                     (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_nativeaddress                                       (slow_peripheral_bridge_m1_nativeaddress),
      .slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave (slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave),
      .slow_peripheral_bridge_m1_read                                                (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave   (slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave),
      .slow_peripheral_bridge_m1_requests_performance_counter_control_slave          (slow_peripheral_bridge_m1_requests_performance_counter_control_slave),
      .slow_peripheral_bridge_m1_write                                               (slow_peripheral_bridge_m1_write),
      .slow_peripheral_bridge_m1_writedata                                           (slow_peripheral_bridge_m1_writedata)
    );

  performance_counter the_performance_counter
    (
      .address       (performance_counter_control_slave_address),
      .begintransfer (performance_counter_control_slave_begintransfer),
      .clk           (pll_c2_out),
      .readdata      (performance_counter_control_slave_readdata),
      .reset_n       (performance_counter_control_slave_reset_n),
      .write         (performance_counter_control_slave_write),
      .writedata     (performance_counter_control_slave_writedata)
    );

  pipeline_bridge_before_tristate_bridge_s1_arbitrator the_pipeline_bridge_before_tristate_bridge_s1
    (
      .clk                                                                                             (pll_c0_out),
      .cpu_data_master_address_to_slave                                                                (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                                      (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                                                     (cpu_data_master_debugaccess),
      .cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1                               (cpu_data_master_granted_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_data_master_latency_counter                                                                 (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1                     (cpu_data_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_data_master_read                                                                            (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                          (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1                       (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register        (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register                        (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register),
      .cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1                              (cpu_data_master_requests_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_data_master_write                                                                           (cpu_data_master_write),
      .cpu_data_master_writedata                                                                       (cpu_data_master_writedata),
      .cpu_instruction_master_address_to_slave                                                         (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1                        (cpu_instruction_master_granted_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_instruction_master_latency_counter                                                          (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1              (cpu_instruction_master_qualified_request_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_instruction_master_read                                                                     (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                   (cpu_instruction_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1                (cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1),
      .cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register (cpu_instruction_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1                       (cpu_instruction_master_requests_pipeline_bridge_before_tristate_bridge_s1),
      .d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer                                           (d1_pipeline_bridge_before_tristate_bridge_s1_end_xfer),
      .pipeline_bridge_before_tristate_bridge_s1_address                                               (pipeline_bridge_before_tristate_bridge_s1_address),
      .pipeline_bridge_before_tristate_bridge_s1_arbiterlock                                           (pipeline_bridge_before_tristate_bridge_s1_arbiterlock),
      .pipeline_bridge_before_tristate_bridge_s1_arbiterlock2                                          (pipeline_bridge_before_tristate_bridge_s1_arbiterlock2),
      .pipeline_bridge_before_tristate_bridge_s1_burstcount                                            (pipeline_bridge_before_tristate_bridge_s1_burstcount),
      .pipeline_bridge_before_tristate_bridge_s1_byteenable                                            (pipeline_bridge_before_tristate_bridge_s1_byteenable),
      .pipeline_bridge_before_tristate_bridge_s1_chipselect                                            (pipeline_bridge_before_tristate_bridge_s1_chipselect),
      .pipeline_bridge_before_tristate_bridge_s1_debugaccess                                           (pipeline_bridge_before_tristate_bridge_s1_debugaccess),
      .pipeline_bridge_before_tristate_bridge_s1_endofpacket                                           (pipeline_bridge_before_tristate_bridge_s1_endofpacket),
      .pipeline_bridge_before_tristate_bridge_s1_endofpacket_from_sa                                   (pipeline_bridge_before_tristate_bridge_s1_endofpacket_from_sa),
      .pipeline_bridge_before_tristate_bridge_s1_nativeaddress                                         (pipeline_bridge_before_tristate_bridge_s1_nativeaddress),
      .pipeline_bridge_before_tristate_bridge_s1_read                                                  (pipeline_bridge_before_tristate_bridge_s1_read),
      .pipeline_bridge_before_tristate_bridge_s1_readdata                                              (pipeline_bridge_before_tristate_bridge_s1_readdata),
      .pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa                                      (pipeline_bridge_before_tristate_bridge_s1_readdata_from_sa),
      .pipeline_bridge_before_tristate_bridge_s1_readdatavalid                                         (pipeline_bridge_before_tristate_bridge_s1_readdatavalid),
      .pipeline_bridge_before_tristate_bridge_s1_reset_n                                               (pipeline_bridge_before_tristate_bridge_s1_reset_n),
      .pipeline_bridge_before_tristate_bridge_s1_waitrequest                                           (pipeline_bridge_before_tristate_bridge_s1_waitrequest),
      .pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa                                   (pipeline_bridge_before_tristate_bridge_s1_waitrequest_from_sa),
      .pipeline_bridge_before_tristate_bridge_s1_write                                                 (pipeline_bridge_before_tristate_bridge_s1_write),
      .pipeline_bridge_before_tristate_bridge_s1_writedata                                             (pipeline_bridge_before_tristate_bridge_s1_writedata),
      .reset_n                                                                                         (pll_c0_out_reset_n)
    );

  pipeline_bridge_before_tristate_bridge_m1_arbitrator the_pipeline_bridge_before_tristate_bridge_m1
    (
      .clk                                                                      (pll_c0_out),
      .d1_flash_tristate_bridge_avalon_slave_end_xfer                           (d1_flash_tristate_bridge_avalon_slave_end_xfer),
      .ext_flash_s1_wait_counter_eq_0                                           (ext_flash_s1_wait_counter_eq_0),
      .incoming_flash_tristate_bridge_data                                      (incoming_flash_tristate_bridge_data),
      .incoming_flash_tristate_bridge_data_with_Xs_converted_to_0               (incoming_flash_tristate_bridge_data_with_Xs_converted_to_0),
      .max2_s1_wait_counter_eq_0                                                (max2_s1_wait_counter_eq_0),
      .pipeline_bridge_before_tristate_bridge_m1_address                        (pipeline_bridge_before_tristate_bridge_m1_address),
      .pipeline_bridge_before_tristate_bridge_m1_address_to_slave               (pipeline_bridge_before_tristate_bridge_m1_address_to_slave),
      .pipeline_bridge_before_tristate_bridge_m1_burstcount                     (pipeline_bridge_before_tristate_bridge_m1_burstcount),
      .pipeline_bridge_before_tristate_bridge_m1_byteenable                     (pipeline_bridge_before_tristate_bridge_m1_byteenable),
      .pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1        (pipeline_bridge_before_tristate_bridge_m1_byteenable_ext_flash_s1),
      .pipeline_bridge_before_tristate_bridge_m1_chipselect                     (pipeline_bridge_before_tristate_bridge_m1_chipselect),
      .pipeline_bridge_before_tristate_bridge_m1_dbs_address                    (pipeline_bridge_before_tristate_bridge_m1_dbs_address),
      .pipeline_bridge_before_tristate_bridge_m1_dbs_write_16                   (pipeline_bridge_before_tristate_bridge_m1_dbs_write_16),
      .pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1           (pipeline_bridge_before_tristate_bridge_m1_granted_ext_flash_s1),
      .pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1                (pipeline_bridge_before_tristate_bridge_m1_granted_max2_s1),
      .pipeline_bridge_before_tristate_bridge_m1_latency_counter                (pipeline_bridge_before_tristate_bridge_m1_latency_counter),
      .pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1 (pipeline_bridge_before_tristate_bridge_m1_qualified_request_ext_flash_s1),
      .pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1      (pipeline_bridge_before_tristate_bridge_m1_qualified_request_max2_s1),
      .pipeline_bridge_before_tristate_bridge_m1_read                           (pipeline_bridge_before_tristate_bridge_m1_read),
      .pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1   (pipeline_bridge_before_tristate_bridge_m1_read_data_valid_ext_flash_s1),
      .pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1        (pipeline_bridge_before_tristate_bridge_m1_read_data_valid_max2_s1),
      .pipeline_bridge_before_tristate_bridge_m1_readdata                       (pipeline_bridge_before_tristate_bridge_m1_readdata),
      .pipeline_bridge_before_tristate_bridge_m1_readdatavalid                  (pipeline_bridge_before_tristate_bridge_m1_readdatavalid),
      .pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1          (pipeline_bridge_before_tristate_bridge_m1_requests_ext_flash_s1),
      .pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1               (pipeline_bridge_before_tristate_bridge_m1_requests_max2_s1),
      .pipeline_bridge_before_tristate_bridge_m1_waitrequest                    (pipeline_bridge_before_tristate_bridge_m1_waitrequest),
      .pipeline_bridge_before_tristate_bridge_m1_write                          (pipeline_bridge_before_tristate_bridge_m1_write),
      .pipeline_bridge_before_tristate_bridge_m1_writedata                      (pipeline_bridge_before_tristate_bridge_m1_writedata),
      .reset_n                                                                  (pll_c0_out_reset_n)
    );

  pipeline_bridge_before_tristate_bridge the_pipeline_bridge_before_tristate_bridge
    (
      .clk              (pll_c0_out),
      .m1_address       (pipeline_bridge_before_tristate_bridge_m1_address),
      .m1_burstcount    (pipeline_bridge_before_tristate_bridge_m1_burstcount),
      .m1_byteenable    (pipeline_bridge_before_tristate_bridge_m1_byteenable),
      .m1_chipselect    (pipeline_bridge_before_tristate_bridge_m1_chipselect),
      .m1_debugaccess   (pipeline_bridge_before_tristate_bridge_m1_debugaccess),
      .m1_endofpacket   (pipeline_bridge_before_tristate_bridge_m1_endofpacket),
      .m1_read          (pipeline_bridge_before_tristate_bridge_m1_read),
      .m1_readdata      (pipeline_bridge_before_tristate_bridge_m1_readdata),
      .m1_readdatavalid (pipeline_bridge_before_tristate_bridge_m1_readdatavalid),
      .m1_waitrequest   (pipeline_bridge_before_tristate_bridge_m1_waitrequest),
      .m1_write         (pipeline_bridge_before_tristate_bridge_m1_write),
      .m1_writedata     (pipeline_bridge_before_tristate_bridge_m1_writedata),
      .reset_n          (pipeline_bridge_before_tristate_bridge_s1_reset_n),
      .s1_address       (pipeline_bridge_before_tristate_bridge_s1_address),
      .s1_arbiterlock   (pipeline_bridge_before_tristate_bridge_s1_arbiterlock),
      .s1_arbiterlock2  (pipeline_bridge_before_tristate_bridge_s1_arbiterlock2),
      .s1_burstcount    (pipeline_bridge_before_tristate_bridge_s1_burstcount),
      .s1_byteenable    (pipeline_bridge_before_tristate_bridge_s1_byteenable),
      .s1_chipselect    (pipeline_bridge_before_tristate_bridge_s1_chipselect),
      .s1_debugaccess   (pipeline_bridge_before_tristate_bridge_s1_debugaccess),
      .s1_endofpacket   (pipeline_bridge_before_tristate_bridge_s1_endofpacket),
      .s1_nativeaddress (pipeline_bridge_before_tristate_bridge_s1_nativeaddress),
      .s1_read          (pipeline_bridge_before_tristate_bridge_s1_read),
      .s1_readdata      (pipeline_bridge_before_tristate_bridge_s1_readdata),
      .s1_readdatavalid (pipeline_bridge_before_tristate_bridge_s1_readdatavalid),
      .s1_waitrequest   (pipeline_bridge_before_tristate_bridge_s1_waitrequest),
      .s1_write         (pipeline_bridge_before_tristate_bridge_s1_write),
      .s1_writedata     (pipeline_bridge_before_tristate_bridge_s1_writedata)
    );

  pll_s1_arbitrator the_pll_s1
    (
      .clk                                                                        (clk),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave         (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_address_to_slave),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1           (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_granted_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_nativeaddress            (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_nativeaddress),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1 (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_qualified_request_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read                     (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_data_valid_pll_s1   (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_read_data_valid_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1          (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_requests_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write                    (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_write),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata                (cycloneIII_3c120_niosII_standard_sopc_clock_0_out_writedata),
      .d1_pll_s1_end_xfer                                                         (d1_pll_s1_end_xfer),
      .pll_s1_address                                                             (pll_s1_address),
      .pll_s1_chipselect                                                          (pll_s1_chipselect),
      .pll_s1_read                                                                (pll_s1_read),
      .pll_s1_readdata                                                            (pll_s1_readdata),
      .pll_s1_readdata_from_sa                                                    (pll_s1_readdata_from_sa),
      .pll_s1_reset_n                                                             (pll_s1_reset_n),
      .pll_s1_resetrequest                                                        (pll_s1_resetrequest),
      .pll_s1_resetrequest_from_sa                                                (pll_s1_resetrequest_from_sa),
      .pll_s1_write                                                               (pll_s1_write),
      .pll_s1_writedata                                                           (pll_s1_writedata),
      .reset_n                                                                    (clk_reset_n)
    );

  //pll_c0_out out_clk assignment, which is an e_assign
  assign pll_c0_out = out_clk_pll_c0;

  //pll_c2_out out_clk assignment, which is an e_assign
  assign pll_c2_out = out_clk_pll_c2;

  //pll_c3_out out_clk assignment, which is an e_assign
  assign pll_c3_out = out_clk_pll_c3;

  //pll_c4_out out_clk assignment, which is an e_assign
  assign pll_c4_out = out_clk_pll_c4;

  pll the_pll
    (
      .address      (pll_s1_address),
      .c0           (out_clk_pll_c0),
      .c2           (out_clk_pll_c2),
      .c3           (out_clk_pll_c3),
      .c4           (out_clk_pll_c4),
      .chipselect   (pll_s1_chipselect),
      .clk          (clk),
      .locked       (locked_from_the_pll),
      .read         (pll_s1_read),
      .readdata     (pll_s1_readdata),
      .reset_n      (pll_s1_reset_n),
      .resetrequest (pll_s1_resetrequest),
      .write        (pll_s1_write),
      .writedata    (pll_s1_writedata)
    );

  sgdma_rx_csr_arbitrator the_sgdma_rx_csr
    (
      .clk                                                                                      (pll_c0_out),
      .cpu_data_master_address_to_slave                                                         (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_sgdma_rx_csr                                                     (cpu_data_master_granted_sgdma_rx_csr),
      .cpu_data_master_latency_counter                                                          (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_sgdma_rx_csr                                           (cpu_data_master_qualified_request_sgdma_rx_csr),
      .cpu_data_master_read                                                                     (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                   (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_sgdma_rx_csr                                             (cpu_data_master_read_data_valid_sgdma_rx_csr),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register                 (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register),
      .cpu_data_master_requests_sgdma_rx_csr                                                    (cpu_data_master_requests_sgdma_rx_csr),
      .cpu_data_master_write                                                                    (cpu_data_master_write),
      .cpu_data_master_writedata                                                                (cpu_data_master_writedata),
      .d1_sgdma_rx_csr_end_xfer                                                                 (d1_sgdma_rx_csr_end_xfer),
      .reset_n                                                                                  (pll_c0_out_reset_n),
      .sgdma_rx_csr_address                                                                     (sgdma_rx_csr_address),
      .sgdma_rx_csr_chipselect                                                                  (sgdma_rx_csr_chipselect),
      .sgdma_rx_csr_irq                                                                         (sgdma_rx_csr_irq),
      .sgdma_rx_csr_irq_from_sa                                                                 (sgdma_rx_csr_irq_from_sa),
      .sgdma_rx_csr_read                                                                        (sgdma_rx_csr_read),
      .sgdma_rx_csr_readdata                                                                    (sgdma_rx_csr_readdata),
      .sgdma_rx_csr_readdata_from_sa                                                            (sgdma_rx_csr_readdata_from_sa),
      .sgdma_rx_csr_reset_n                                                                     (sgdma_rx_csr_reset_n),
      .sgdma_rx_csr_write                                                                       (sgdma_rx_csr_write),
      .sgdma_rx_csr_writedata                                                                   (sgdma_rx_csr_writedata)
    );

  sgdma_rx_in_arbitrator the_sgdma_rx_in
    (
      .clk                           (pll_c0_out),
      .reset_n                       (pll_c0_out_reset_n),
      .sgdma_rx_in_data              (sgdma_rx_in_data),
      .sgdma_rx_in_empty             (sgdma_rx_in_empty),
      .sgdma_rx_in_endofpacket       (sgdma_rx_in_endofpacket),
      .sgdma_rx_in_error             (sgdma_rx_in_error),
      .sgdma_rx_in_ready             (sgdma_rx_in_ready),
      .sgdma_rx_in_ready_from_sa     (sgdma_rx_in_ready_from_sa),
      .sgdma_rx_in_startofpacket     (sgdma_rx_in_startofpacket),
      .sgdma_rx_in_valid             (sgdma_rx_in_valid),
      .tse_mac_receive_data          (tse_mac_receive_data),
      .tse_mac_receive_empty         (tse_mac_receive_empty),
      .tse_mac_receive_endofpacket   (tse_mac_receive_endofpacket),
      .tse_mac_receive_error         (tse_mac_receive_error),
      .tse_mac_receive_startofpacket (tse_mac_receive_startofpacket),
      .tse_mac_receive_valid         (tse_mac_receive_valid)
    );

  sgdma_rx_descriptor_read_arbitrator the_sgdma_rx_descriptor_read
    (
      .clk                                                             (pll_c0_out),
      .d1_descriptor_memory_s1_end_xfer                                (d1_descriptor_memory_s1_end_xfer),
      .descriptor_memory_s1_readdata_from_sa                           (descriptor_memory_s1_readdata_from_sa),
      .reset_n                                                         (pll_c0_out_reset_n),
      .sgdma_rx_descriptor_read_address                                (sgdma_rx_descriptor_read_address),
      .sgdma_rx_descriptor_read_address_to_slave                       (sgdma_rx_descriptor_read_address_to_slave),
      .sgdma_rx_descriptor_read_granted_descriptor_memory_s1           (sgdma_rx_descriptor_read_granted_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_latency_counter                        (sgdma_rx_descriptor_read_latency_counter),
      .sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 (sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_read                                   (sgdma_rx_descriptor_read_read),
      .sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1   (sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_readdata                               (sgdma_rx_descriptor_read_readdata),
      .sgdma_rx_descriptor_read_readdatavalid                          (sgdma_rx_descriptor_read_readdatavalid),
      .sgdma_rx_descriptor_read_requests_descriptor_memory_s1          (sgdma_rx_descriptor_read_requests_descriptor_memory_s1),
      .sgdma_rx_descriptor_read_waitrequest                            (sgdma_rx_descriptor_read_waitrequest)
    );

  sgdma_rx_descriptor_write_arbitrator the_sgdma_rx_descriptor_write
    (
      .clk                                                              (pll_c0_out),
      .d1_descriptor_memory_s1_end_xfer                                 (d1_descriptor_memory_s1_end_xfer),
      .reset_n                                                          (pll_c0_out_reset_n),
      .sgdma_rx_descriptor_write_address                                (sgdma_rx_descriptor_write_address),
      .sgdma_rx_descriptor_write_address_to_slave                       (sgdma_rx_descriptor_write_address_to_slave),
      .sgdma_rx_descriptor_write_granted_descriptor_memory_s1           (sgdma_rx_descriptor_write_granted_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 (sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_requests_descriptor_memory_s1          (sgdma_rx_descriptor_write_requests_descriptor_memory_s1),
      .sgdma_rx_descriptor_write_waitrequest                            (sgdma_rx_descriptor_write_waitrequest),
      .sgdma_rx_descriptor_write_write                                  (sgdma_rx_descriptor_write_write),
      .sgdma_rx_descriptor_write_writedata                              (sgdma_rx_descriptor_write_writedata)
    );

  sgdma_rx_m_write_arbitrator the_sgdma_rx_m_write
    (
      .clk                                                        (pll_c0_out),
      .cpu_ddr_clock_bridge_s1_waitrequest_from_sa                (cpu_ddr_clock_bridge_s1_waitrequest_from_sa),
      .d1_cpu_ddr_clock_bridge_s1_end_xfer                        (d1_cpu_ddr_clock_bridge_s1_end_xfer),
      .reset_n                                                    (pll_c0_out_reset_n),
      .sgdma_rx_m_write_address                                   (sgdma_rx_m_write_address),
      .sgdma_rx_m_write_address_to_slave                          (sgdma_rx_m_write_address_to_slave),
      .sgdma_rx_m_write_byteenable                                (sgdma_rx_m_write_byteenable),
      .sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1           (sgdma_rx_m_write_granted_cpu_ddr_clock_bridge_s1),
      .sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1 (sgdma_rx_m_write_qualified_request_cpu_ddr_clock_bridge_s1),
      .sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1          (sgdma_rx_m_write_requests_cpu_ddr_clock_bridge_s1),
      .sgdma_rx_m_write_waitrequest                               (sgdma_rx_m_write_waitrequest),
      .sgdma_rx_m_write_write                                     (sgdma_rx_m_write_write),
      .sgdma_rx_m_write_writedata                                 (sgdma_rx_m_write_writedata)
    );

  sgdma_rx the_sgdma_rx
    (
      .clk                           (pll_c0_out),
      .csr_address                   (sgdma_rx_csr_address),
      .csr_chipselect                (sgdma_rx_csr_chipselect),
      .csr_irq                       (sgdma_rx_csr_irq),
      .csr_read                      (sgdma_rx_csr_read),
      .csr_readdata                  (sgdma_rx_csr_readdata),
      .csr_write                     (sgdma_rx_csr_write),
      .csr_writedata                 (sgdma_rx_csr_writedata),
      .descriptor_read_address       (sgdma_rx_descriptor_read_address),
      .descriptor_read_read          (sgdma_rx_descriptor_read_read),
      .descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),
      .descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),
      .descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),
      .descriptor_write_address      (sgdma_rx_descriptor_write_address),
      .descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),
      .descriptor_write_write        (sgdma_rx_descriptor_write_write),
      .descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),
      .in_data                       (sgdma_rx_in_data),
      .in_empty                      (sgdma_rx_in_empty),
      .in_endofpacket                (sgdma_rx_in_endofpacket),
      .in_error                      (sgdma_rx_in_error),
      .in_ready                      (sgdma_rx_in_ready),
      .in_startofpacket              (sgdma_rx_in_startofpacket),
      .in_valid                      (sgdma_rx_in_valid),
      .m_write_address               (sgdma_rx_m_write_address),
      .m_write_byteenable            (sgdma_rx_m_write_byteenable),
      .m_write_waitrequest           (sgdma_rx_m_write_waitrequest),
      .m_write_write                 (sgdma_rx_m_write_write),
      .m_write_writedata             (sgdma_rx_m_write_writedata),
      .system_reset_n                (sgdma_rx_csr_reset_n)
    );

  sgdma_tx_csr_arbitrator the_sgdma_tx_csr
    (
      .clk                                                                                      (pll_c0_out),
      .cpu_data_master_address_to_slave                                                         (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_sgdma_tx_csr                                                     (cpu_data_master_granted_sgdma_tx_csr),
      .cpu_data_master_latency_counter                                                          (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_sgdma_tx_csr                                           (cpu_data_master_qualified_request_sgdma_tx_csr),
      .cpu_data_master_read                                                                     (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                   (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_sgdma_tx_csr                                             (cpu_data_master_read_data_valid_sgdma_tx_csr),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register                 (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register),
      .cpu_data_master_requests_sgdma_tx_csr                                                    (cpu_data_master_requests_sgdma_tx_csr),
      .cpu_data_master_write                                                                    (cpu_data_master_write),
      .cpu_data_master_writedata                                                                (cpu_data_master_writedata),
      .d1_sgdma_tx_csr_end_xfer                                                                 (d1_sgdma_tx_csr_end_xfer),
      .reset_n                                                                                  (pll_c0_out_reset_n),
      .sgdma_tx_csr_address                                                                     (sgdma_tx_csr_address),
      .sgdma_tx_csr_chipselect                                                                  (sgdma_tx_csr_chipselect),
      .sgdma_tx_csr_irq                                                                         (sgdma_tx_csr_irq),
      .sgdma_tx_csr_irq_from_sa                                                                 (sgdma_tx_csr_irq_from_sa),
      .sgdma_tx_csr_read                                                                        (sgdma_tx_csr_read),
      .sgdma_tx_csr_readdata                                                                    (sgdma_tx_csr_readdata),
      .sgdma_tx_csr_readdata_from_sa                                                            (sgdma_tx_csr_readdata_from_sa),
      .sgdma_tx_csr_reset_n                                                                     (sgdma_tx_csr_reset_n),
      .sgdma_tx_csr_write                                                                       (sgdma_tx_csr_write),
      .sgdma_tx_csr_writedata                                                                   (sgdma_tx_csr_writedata)
    );

  sgdma_tx_descriptor_read_arbitrator the_sgdma_tx_descriptor_read
    (
      .clk                                                             (pll_c0_out),
      .d1_descriptor_memory_s1_end_xfer                                (d1_descriptor_memory_s1_end_xfer),
      .descriptor_memory_s1_readdata_from_sa                           (descriptor_memory_s1_readdata_from_sa),
      .reset_n                                                         (pll_c0_out_reset_n),
      .sgdma_tx_descriptor_read_address                                (sgdma_tx_descriptor_read_address),
      .sgdma_tx_descriptor_read_address_to_slave                       (sgdma_tx_descriptor_read_address_to_slave),
      .sgdma_tx_descriptor_read_granted_descriptor_memory_s1           (sgdma_tx_descriptor_read_granted_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_latency_counter                        (sgdma_tx_descriptor_read_latency_counter),
      .sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 (sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_read                                   (sgdma_tx_descriptor_read_read),
      .sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1   (sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_readdata                               (sgdma_tx_descriptor_read_readdata),
      .sgdma_tx_descriptor_read_readdatavalid                          (sgdma_tx_descriptor_read_readdatavalid),
      .sgdma_tx_descriptor_read_requests_descriptor_memory_s1          (sgdma_tx_descriptor_read_requests_descriptor_memory_s1),
      .sgdma_tx_descriptor_read_waitrequest                            (sgdma_tx_descriptor_read_waitrequest)
    );

  sgdma_tx_descriptor_write_arbitrator the_sgdma_tx_descriptor_write
    (
      .clk                                                              (pll_c0_out),
      .d1_descriptor_memory_s1_end_xfer                                 (d1_descriptor_memory_s1_end_xfer),
      .reset_n                                                          (pll_c0_out_reset_n),
      .sgdma_tx_descriptor_write_address                                (sgdma_tx_descriptor_write_address),
      .sgdma_tx_descriptor_write_address_to_slave                       (sgdma_tx_descriptor_write_address_to_slave),
      .sgdma_tx_descriptor_write_granted_descriptor_memory_s1           (sgdma_tx_descriptor_write_granted_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 (sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_requests_descriptor_memory_s1          (sgdma_tx_descriptor_write_requests_descriptor_memory_s1),
      .sgdma_tx_descriptor_write_waitrequest                            (sgdma_tx_descriptor_write_waitrequest),
      .sgdma_tx_descriptor_write_write                                  (sgdma_tx_descriptor_write_write),
      .sgdma_tx_descriptor_write_writedata                              (sgdma_tx_descriptor_write_writedata)
    );

  sgdma_tx_m_read_arbitrator the_sgdma_tx_m_read
    (
      .clk                                                                    (pll_c0_out),
      .cpu_ddr_clock_bridge_s1_readdata_from_sa                               (cpu_ddr_clock_bridge_s1_readdata_from_sa),
      .cpu_ddr_clock_bridge_s1_waitrequest_from_sa                            (cpu_ddr_clock_bridge_s1_waitrequest_from_sa),
      .d1_cpu_ddr_clock_bridge_s1_end_xfer                                    (d1_cpu_ddr_clock_bridge_s1_end_xfer),
      .reset_n                                                                (pll_c0_out_reset_n),
      .sgdma_tx_m_read_address                                                (sgdma_tx_m_read_address),
      .sgdma_tx_m_read_address_to_slave                                       (sgdma_tx_m_read_address_to_slave),
      .sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1                        (sgdma_tx_m_read_granted_cpu_ddr_clock_bridge_s1),
      .sgdma_tx_m_read_latency_counter                                        (sgdma_tx_m_read_latency_counter),
      .sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1              (sgdma_tx_m_read_qualified_request_cpu_ddr_clock_bridge_s1),
      .sgdma_tx_m_read_read                                                   (sgdma_tx_m_read_read),
      .sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1                (sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1),
      .sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register (sgdma_tx_m_read_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .sgdma_tx_m_read_readdata                                               (sgdma_tx_m_read_readdata),
      .sgdma_tx_m_read_readdatavalid                                          (sgdma_tx_m_read_readdatavalid),
      .sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1                       (sgdma_tx_m_read_requests_cpu_ddr_clock_bridge_s1),
      .sgdma_tx_m_read_waitrequest                                            (sgdma_tx_m_read_waitrequest)
    );

  sgdma_tx_out_arbitrator the_sgdma_tx_out
    (
      .clk                            (pll_c0_out),
      .reset_n                        (pll_c0_out_reset_n),
      .sgdma_tx_out_data              (sgdma_tx_out_data),
      .sgdma_tx_out_empty             (sgdma_tx_out_empty),
      .sgdma_tx_out_endofpacket       (sgdma_tx_out_endofpacket),
      .sgdma_tx_out_error             (sgdma_tx_out_error),
      .sgdma_tx_out_ready             (sgdma_tx_out_ready),
      .sgdma_tx_out_startofpacket     (sgdma_tx_out_startofpacket),
      .sgdma_tx_out_valid             (sgdma_tx_out_valid),
      .tse_mac_transmit_ready_from_sa (tse_mac_transmit_ready_from_sa)
    );

  sgdma_tx the_sgdma_tx
    (
      .clk                           (pll_c0_out),
      .csr_address                   (sgdma_tx_csr_address),
      .csr_chipselect                (sgdma_tx_csr_chipselect),
      .csr_irq                       (sgdma_tx_csr_irq),
      .csr_read                      (sgdma_tx_csr_read),
      .csr_readdata                  (sgdma_tx_csr_readdata),
      .csr_write                     (sgdma_tx_csr_write),
      .csr_writedata                 (sgdma_tx_csr_writedata),
      .descriptor_read_address       (sgdma_tx_descriptor_read_address),
      .descriptor_read_read          (sgdma_tx_descriptor_read_read),
      .descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),
      .descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),
      .descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),
      .descriptor_write_address      (sgdma_tx_descriptor_write_address),
      .descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),
      .descriptor_write_write        (sgdma_tx_descriptor_write_write),
      .descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),
      .m_read_address                (sgdma_tx_m_read_address),
      .m_read_read                   (sgdma_tx_m_read_read),
      .m_read_readdata               (sgdma_tx_m_read_readdata),
      .m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),
      .m_read_waitrequest            (sgdma_tx_m_read_waitrequest),
      .out_data                      (sgdma_tx_out_data),
      .out_empty                     (sgdma_tx_out_empty),
      .out_endofpacket               (sgdma_tx_out_endofpacket),
      .out_error                     (sgdma_tx_out_error),
      .out_ready                     (sgdma_tx_out_ready),
      .out_startofpacket             (sgdma_tx_out_startofpacket),
      .out_valid                     (sgdma_tx_out_valid),
      .system_reset_n                (sgdma_tx_csr_reset_n)
    );

  slow_peripheral_bridge_s1_arbitrator the_slow_peripheral_bridge_s1
    (
      .clk                                                                                      (pll_c0_out),
      .cpu_data_master_address_to_slave                                                         (cpu_data_master_address_to_slave),
      .cpu_data_master_byteenable                                                               (cpu_data_master_byteenable),
      .cpu_data_master_granted_slow_peripheral_bridge_s1                                        (cpu_data_master_granted_slow_peripheral_bridge_s1),
      .cpu_data_master_latency_counter                                                          (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_slow_peripheral_bridge_s1                              (cpu_data_master_qualified_request_slow_peripheral_bridge_s1),
      .cpu_data_master_read                                                                     (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                   (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1                                (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register                 (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register),
      .cpu_data_master_requests_slow_peripheral_bridge_s1                                       (cpu_data_master_requests_slow_peripheral_bridge_s1),
      .cpu_data_master_write                                                                    (cpu_data_master_write),
      .cpu_data_master_writedata                                                                (cpu_data_master_writedata),
      .d1_slow_peripheral_bridge_s1_end_xfer                                                    (d1_slow_peripheral_bridge_s1_end_xfer),
      .reset_n                                                                                  (pll_c0_out_reset_n),
      .slow_peripheral_bridge_s1_address                                                        (slow_peripheral_bridge_s1_address),
      .slow_peripheral_bridge_s1_byteenable                                                     (slow_peripheral_bridge_s1_byteenable),
      .slow_peripheral_bridge_s1_endofpacket                                                    (slow_peripheral_bridge_s1_endofpacket),
      .slow_peripheral_bridge_s1_endofpacket_from_sa                                            (slow_peripheral_bridge_s1_endofpacket_from_sa),
      .slow_peripheral_bridge_s1_nativeaddress                                                  (slow_peripheral_bridge_s1_nativeaddress),
      .slow_peripheral_bridge_s1_read                                                           (slow_peripheral_bridge_s1_read),
      .slow_peripheral_bridge_s1_readdata                                                       (slow_peripheral_bridge_s1_readdata),
      .slow_peripheral_bridge_s1_readdata_from_sa                                               (slow_peripheral_bridge_s1_readdata_from_sa),
      .slow_peripheral_bridge_s1_readdatavalid                                                  (slow_peripheral_bridge_s1_readdatavalid),
      .slow_peripheral_bridge_s1_reset_n                                                        (slow_peripheral_bridge_s1_reset_n),
      .slow_peripheral_bridge_s1_waitrequest                                                    (slow_peripheral_bridge_s1_waitrequest),
      .slow_peripheral_bridge_s1_waitrequest_from_sa                                            (slow_peripheral_bridge_s1_waitrequest_from_sa),
      .slow_peripheral_bridge_s1_write                                                          (slow_peripheral_bridge_s1_write),
      .slow_peripheral_bridge_s1_writedata                                                      (slow_peripheral_bridge_s1_writedata)
    );

  slow_peripheral_bridge_m1_arbitrator the_slow_peripheral_bridge_m1
    (
      .button_pio_s1_readdata_from_sa                                                               (button_pio_s1_readdata_from_sa),
      .clk                                                                                          (pll_c2_out),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_endofpacket_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa                            (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_readdata_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_0_in_waitrequest_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_endofpacket_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa                            (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_readdata_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_1_in_waitrequest_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_endofpacket_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa                            (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_readdata_from_sa),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa                         (cycloneIII_3c120_niosII_standard_sopc_clock_2_in_waitrequest_from_sa),
      .d1_button_pio_s1_end_xfer                                                                    (d1_button_pio_s1_end_xfer),
      .d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer                                 (d1_cycloneIII_3c120_niosII_standard_sopc_clock_0_in_end_xfer),
      .d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer                                 (d1_cycloneIII_3c120_niosII_standard_sopc_clock_1_in_end_xfer),
      .d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer                                 (d1_cycloneIII_3c120_niosII_standard_sopc_clock_2_in_end_xfer),
      .d1_high_res_timer_s1_end_xfer                                                                (d1_high_res_timer_s1_end_xfer),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                                                      (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .d1_led_pio_s1_end_xfer                                                                       (d1_led_pio_s1_end_xfer),
      .d1_performance_counter_control_slave_end_xfer                                                (d1_performance_counter_control_slave_end_xfer),
      .d1_sys_clk_timer_s1_end_xfer                                                                 (d1_sys_clk_timer_s1_end_xfer),
      .d1_sysid_control_slave_end_xfer                                                              (d1_sysid_control_slave_end_xfer),
      .high_res_timer_s1_readdata_from_sa                                                           (high_res_timer_s1_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                                                 (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa                                              (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .led_pio_s1_readdata_from_sa                                                                  (led_pio_s1_readdata_from_sa),
      .performance_counter_control_slave_readdata_from_sa                                           (performance_counter_control_slave_readdata_from_sa),
      .reset_n                                                                                      (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address                                                            (slow_peripheral_bridge_m1_address),
      .slow_peripheral_bridge_m1_address_to_slave                                                   (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_byteenable                                                         (slow_peripheral_bridge_m1_byteenable),
      .slow_peripheral_bridge_m1_endofpacket                                                        (slow_peripheral_bridge_m1_endofpacket),
      .slow_peripheral_bridge_m1_granted_button_pio_s1                                              (slow_peripheral_bridge_m1_granted_button_pio_s1),
      .slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in           (slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_0_in),
      .slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in           (slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_1_in),
      .slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in           (slow_peripheral_bridge_m1_granted_cycloneIII_3c120_niosII_standard_sopc_clock_2_in),
      .slow_peripheral_bridge_m1_granted_high_res_timer_s1                                          (slow_peripheral_bridge_m1_granted_high_res_timer_s1),
      .slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave                                (slow_peripheral_bridge_m1_granted_jtag_uart_avalon_jtag_slave),
      .slow_peripheral_bridge_m1_granted_led_pio_s1                                                 (slow_peripheral_bridge_m1_granted_led_pio_s1),
      .slow_peripheral_bridge_m1_granted_performance_counter_control_slave                          (slow_peripheral_bridge_m1_granted_performance_counter_control_slave),
      .slow_peripheral_bridge_m1_granted_sys_clk_timer_s1                                           (slow_peripheral_bridge_m1_granted_sys_clk_timer_s1),
      .slow_peripheral_bridge_m1_granted_sysid_control_slave                                        (slow_peripheral_bridge_m1_granted_sysid_control_slave),
      .slow_peripheral_bridge_m1_latency_counter                                                    (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_qualified_request_button_pio_s1                                    (slow_peripheral_bridge_m1_qualified_request_button_pio_s1),
      .slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in (slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_0_in),
      .slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in (slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_1_in),
      .slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in (slow_peripheral_bridge_m1_qualified_request_cycloneIII_3c120_niosII_standard_sopc_clock_2_in),
      .slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1                                (slow_peripheral_bridge_m1_qualified_request_high_res_timer_s1),
      .slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave                      (slow_peripheral_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave),
      .slow_peripheral_bridge_m1_qualified_request_led_pio_s1                                       (slow_peripheral_bridge_m1_qualified_request_led_pio_s1),
      .slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave                (slow_peripheral_bridge_m1_qualified_request_performance_counter_control_slave),
      .slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1                                 (slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1),
      .slow_peripheral_bridge_m1_qualified_request_sysid_control_slave                              (slow_peripheral_bridge_m1_qualified_request_sysid_control_slave),
      .slow_peripheral_bridge_m1_read                                                               (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_button_pio_s1                                      (slow_peripheral_bridge_m1_read_data_valid_button_pio_s1),
      .slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in   (slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_0_in),
      .slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in   (slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_1_in),
      .slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in   (slow_peripheral_bridge_m1_read_data_valid_cycloneIII_3c120_niosII_standard_sopc_clock_2_in),
      .slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1                                  (slow_peripheral_bridge_m1_read_data_valid_high_res_timer_s1),
      .slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave                        (slow_peripheral_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave),
      .slow_peripheral_bridge_m1_read_data_valid_led_pio_s1                                         (slow_peripheral_bridge_m1_read_data_valid_led_pio_s1),
      .slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave                  (slow_peripheral_bridge_m1_read_data_valid_performance_counter_control_slave),
      .slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1                                   (slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1),
      .slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave                                (slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave),
      .slow_peripheral_bridge_m1_readdata                                                           (slow_peripheral_bridge_m1_readdata),
      .slow_peripheral_bridge_m1_readdatavalid                                                      (slow_peripheral_bridge_m1_readdatavalid),
      .slow_peripheral_bridge_m1_requests_button_pio_s1                                             (slow_peripheral_bridge_m1_requests_button_pio_s1),
      .slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in          (slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_0_in),
      .slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in          (slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_1_in),
      .slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in          (slow_peripheral_bridge_m1_requests_cycloneIII_3c120_niosII_standard_sopc_clock_2_in),
      .slow_peripheral_bridge_m1_requests_high_res_timer_s1                                         (slow_peripheral_bridge_m1_requests_high_res_timer_s1),
      .slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave                               (slow_peripheral_bridge_m1_requests_jtag_uart_avalon_jtag_slave),
      .slow_peripheral_bridge_m1_requests_led_pio_s1                                                (slow_peripheral_bridge_m1_requests_led_pio_s1),
      .slow_peripheral_bridge_m1_requests_performance_counter_control_slave                         (slow_peripheral_bridge_m1_requests_performance_counter_control_slave),
      .slow_peripheral_bridge_m1_requests_sys_clk_timer_s1                                          (slow_peripheral_bridge_m1_requests_sys_clk_timer_s1),
      .slow_peripheral_bridge_m1_requests_sysid_control_slave                                       (slow_peripheral_bridge_m1_requests_sysid_control_slave),
      .slow_peripheral_bridge_m1_reset_n                                                            (slow_peripheral_bridge_m1_reset_n),
      .slow_peripheral_bridge_m1_waitrequest                                                        (slow_peripheral_bridge_m1_waitrequest),
      .slow_peripheral_bridge_m1_write                                                              (slow_peripheral_bridge_m1_write),
      .slow_peripheral_bridge_m1_writedata                                                          (slow_peripheral_bridge_m1_writedata),
      .sys_clk_timer_s1_readdata_from_sa                                                            (sys_clk_timer_s1_readdata_from_sa),
      .sysid_control_slave_readdata_from_sa                                                         (sysid_control_slave_readdata_from_sa)
    );

  slow_peripheral_bridge the_slow_peripheral_bridge
    (
      .master_address       (slow_peripheral_bridge_m1_address),
      .master_byteenable    (slow_peripheral_bridge_m1_byteenable),
      .master_clk           (pll_c2_out),
      .master_endofpacket   (slow_peripheral_bridge_m1_endofpacket),
      .master_nativeaddress (slow_peripheral_bridge_m1_nativeaddress),
      .master_read          (slow_peripheral_bridge_m1_read),
      .master_readdata      (slow_peripheral_bridge_m1_readdata),
      .master_readdatavalid (slow_peripheral_bridge_m1_readdatavalid),
      .master_reset_n       (slow_peripheral_bridge_m1_reset_n),
      .master_waitrequest   (slow_peripheral_bridge_m1_waitrequest),
      .master_write         (slow_peripheral_bridge_m1_write),
      .master_writedata     (slow_peripheral_bridge_m1_writedata),
      .slave_address        (slow_peripheral_bridge_s1_address),
      .slave_byteenable     (slow_peripheral_bridge_s1_byteenable),
      .slave_clk            (pll_c0_out),
      .slave_endofpacket    (slow_peripheral_bridge_s1_endofpacket),
      .slave_nativeaddress  (slow_peripheral_bridge_s1_nativeaddress),
      .slave_read           (slow_peripheral_bridge_s1_read),
      .slave_readdata       (slow_peripheral_bridge_s1_readdata),
      .slave_readdatavalid  (slow_peripheral_bridge_s1_readdatavalid),
      .slave_reset_n        (slow_peripheral_bridge_s1_reset_n),
      .slave_waitrequest    (slow_peripheral_bridge_s1_waitrequest),
      .slave_write          (slow_peripheral_bridge_s1_write),
      .slave_writedata      (slow_peripheral_bridge_s1_writedata)
    );

  sys_clk_timer_s1_arbitrator the_sys_clk_timer_s1
    (
      .clk                                                          (pll_c2_out),
      .d1_sys_clk_timer_s1_end_xfer                                 (d1_sys_clk_timer_s1_end_xfer),
      .reset_n                                                      (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address_to_slave                   (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_granted_sys_clk_timer_s1           (slow_peripheral_bridge_m1_granted_sys_clk_timer_s1),
      .slow_peripheral_bridge_m1_latency_counter                    (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_nativeaddress                      (slow_peripheral_bridge_m1_nativeaddress),
      .slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1 (slow_peripheral_bridge_m1_qualified_request_sys_clk_timer_s1),
      .slow_peripheral_bridge_m1_read                               (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1   (slow_peripheral_bridge_m1_read_data_valid_sys_clk_timer_s1),
      .slow_peripheral_bridge_m1_requests_sys_clk_timer_s1          (slow_peripheral_bridge_m1_requests_sys_clk_timer_s1),
      .slow_peripheral_bridge_m1_write                              (slow_peripheral_bridge_m1_write),
      .slow_peripheral_bridge_m1_writedata                          (slow_peripheral_bridge_m1_writedata),
      .sys_clk_timer_s1_address                                     (sys_clk_timer_s1_address),
      .sys_clk_timer_s1_chipselect                                  (sys_clk_timer_s1_chipselect),
      .sys_clk_timer_s1_irq                                         (sys_clk_timer_s1_irq),
      .sys_clk_timer_s1_irq_from_sa                                 (sys_clk_timer_s1_irq_from_sa),
      .sys_clk_timer_s1_readdata                                    (sys_clk_timer_s1_readdata),
      .sys_clk_timer_s1_readdata_from_sa                            (sys_clk_timer_s1_readdata_from_sa),
      .sys_clk_timer_s1_reset_n                                     (sys_clk_timer_s1_reset_n),
      .sys_clk_timer_s1_write_n                                     (sys_clk_timer_s1_write_n),
      .sys_clk_timer_s1_writedata                                   (sys_clk_timer_s1_writedata)
    );

  sys_clk_timer the_sys_clk_timer
    (
      .address    (sys_clk_timer_s1_address),
      .chipselect (sys_clk_timer_s1_chipselect),
      .clk        (pll_c2_out),
      .irq        (sys_clk_timer_s1_irq),
      .readdata   (sys_clk_timer_s1_readdata),
      .reset_n    (sys_clk_timer_s1_reset_n),
      .write_n    (sys_clk_timer_s1_write_n),
      .writedata  (sys_clk_timer_s1_writedata)
    );

  sysid_control_slave_arbitrator the_sysid_control_slave
    (
      .clk                                                             (pll_c2_out),
      .d1_sysid_control_slave_end_xfer                                 (d1_sysid_control_slave_end_xfer),
      .reset_n                                                         (pll_c2_out_reset_n),
      .slow_peripheral_bridge_m1_address_to_slave                      (slow_peripheral_bridge_m1_address_to_slave),
      .slow_peripheral_bridge_m1_granted_sysid_control_slave           (slow_peripheral_bridge_m1_granted_sysid_control_slave),
      .slow_peripheral_bridge_m1_latency_counter                       (slow_peripheral_bridge_m1_latency_counter),
      .slow_peripheral_bridge_m1_nativeaddress                         (slow_peripheral_bridge_m1_nativeaddress),
      .slow_peripheral_bridge_m1_qualified_request_sysid_control_slave (slow_peripheral_bridge_m1_qualified_request_sysid_control_slave),
      .slow_peripheral_bridge_m1_read                                  (slow_peripheral_bridge_m1_read),
      .slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave   (slow_peripheral_bridge_m1_read_data_valid_sysid_control_slave),
      .slow_peripheral_bridge_m1_requests_sysid_control_slave          (slow_peripheral_bridge_m1_requests_sysid_control_slave),
      .slow_peripheral_bridge_m1_write                                 (slow_peripheral_bridge_m1_write),
      .sysid_control_slave_address                                     (sysid_control_slave_address),
      .sysid_control_slave_readdata                                    (sysid_control_slave_readdata),
      .sysid_control_slave_readdata_from_sa                            (sysid_control_slave_readdata_from_sa),
      .sysid_control_slave_reset_n                                     (sysid_control_slave_reset_n)
    );

  sysid the_sysid
    (
      .address  (sysid_control_slave_address),
      .clock    (sysid_control_slave_clock),
      .readdata (sysid_control_slave_readdata),
      .reset_n  (sysid_control_slave_reset_n)
    );

  tse_mac_control_port_arbitrator the_tse_mac_control_port
    (
      .clk                                                                                      (pll_c0_out),
      .cpu_data_master_address_to_slave                                                         (cpu_data_master_address_to_slave),
      .cpu_data_master_granted_tse_mac_control_port                                             (cpu_data_master_granted_tse_mac_control_port),
      .cpu_data_master_latency_counter                                                          (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_tse_mac_control_port                                   (cpu_data_master_qualified_request_tse_mac_control_port),
      .cpu_data_master_read                                                                     (cpu_data_master_read),
      .cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register                   (cpu_data_master_read_data_valid_cpu_ddr_clock_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register (cpu_data_master_read_data_valid_pipeline_bridge_before_tristate_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register                 (cpu_data_master_read_data_valid_slow_peripheral_bridge_s1_shift_register),
      .cpu_data_master_read_data_valid_tse_mac_control_port                                     (cpu_data_master_read_data_valid_tse_mac_control_port),
      .cpu_data_master_requests_tse_mac_control_port                                            (cpu_data_master_requests_tse_mac_control_port),
      .cpu_data_master_write                                                                    (cpu_data_master_write),
      .cpu_data_master_writedata                                                                (cpu_data_master_writedata),
      .d1_tse_mac_control_port_end_xfer                                                         (d1_tse_mac_control_port_end_xfer),
      .reset_n                                                                                  (pll_c0_out_reset_n),
      .tse_mac_control_port_address                                                             (tse_mac_control_port_address),
      .tse_mac_control_port_read                                                                (tse_mac_control_port_read),
      .tse_mac_control_port_readdata                                                            (tse_mac_control_port_readdata),
      .tse_mac_control_port_readdata_from_sa                                                    (tse_mac_control_port_readdata_from_sa),
      .tse_mac_control_port_reset                                                               (tse_mac_control_port_reset),
      .tse_mac_control_port_waitrequest                                                         (tse_mac_control_port_waitrequest),
      .tse_mac_control_port_waitrequest_from_sa                                                 (tse_mac_control_port_waitrequest_from_sa),
      .tse_mac_control_port_write                                                               (tse_mac_control_port_write),
      .tse_mac_control_port_writedata                                                           (tse_mac_control_port_writedata)
    );

  tse_mac_transmit_arbitrator the_tse_mac_transmit
    (
      .clk                            (pll_c0_out),
      .reset_n                        (pll_c0_out_reset_n),
      .sgdma_tx_out_data              (sgdma_tx_out_data),
      .sgdma_tx_out_empty             (sgdma_tx_out_empty),
      .sgdma_tx_out_endofpacket       (sgdma_tx_out_endofpacket),
      .sgdma_tx_out_error             (sgdma_tx_out_error),
      .sgdma_tx_out_startofpacket     (sgdma_tx_out_startofpacket),
      .sgdma_tx_out_valid             (sgdma_tx_out_valid),
      .tse_mac_transmit_data          (tse_mac_transmit_data),
      .tse_mac_transmit_empty         (tse_mac_transmit_empty),
      .tse_mac_transmit_endofpacket   (tse_mac_transmit_endofpacket),
      .tse_mac_transmit_error         (tse_mac_transmit_error),
      .tse_mac_transmit_ready         (tse_mac_transmit_ready),
      .tse_mac_transmit_ready_from_sa (tse_mac_transmit_ready_from_sa),
      .tse_mac_transmit_startofpacket (tse_mac_transmit_startofpacket),
      .tse_mac_transmit_valid         (tse_mac_transmit_valid)
    );

  tse_mac_receive_arbitrator the_tse_mac_receive
    (
      .clk                           (pll_c0_out),
      .reset_n                       (pll_c0_out_reset_n),
      .sgdma_rx_in_ready_from_sa     (sgdma_rx_in_ready_from_sa),
      .tse_mac_receive_data          (tse_mac_receive_data),
      .tse_mac_receive_empty         (tse_mac_receive_empty),
      .tse_mac_receive_endofpacket   (tse_mac_receive_endofpacket),
      .tse_mac_receive_error         (tse_mac_receive_error),
      .tse_mac_receive_ready         (tse_mac_receive_ready),
      .tse_mac_receive_startofpacket (tse_mac_receive_startofpacket),
      .tse_mac_receive_valid         (tse_mac_receive_valid)
    );

  tse_mac the_tse_mac
    (
      .address     (tse_mac_control_port_address),
      .clk         (pll_c0_out),
      .ena_10      (ena_10_from_the_tse_mac),
      .eth_mode    (eth_mode_from_the_tse_mac),
      .ff_rx_clk   (pll_c0_out),
      .ff_rx_data  (tse_mac_receive_data),
      .ff_rx_dval  (tse_mac_receive_valid),
      .ff_rx_eop   (tse_mac_receive_endofpacket),
      .ff_rx_mod   (tse_mac_receive_empty),
      .ff_rx_rdy   (tse_mac_receive_ready),
      .ff_rx_sop   (tse_mac_receive_startofpacket),
      .ff_tx_clk   (pll_c0_out),
      .ff_tx_data  (tse_mac_transmit_data),
      .ff_tx_eop   (tse_mac_transmit_endofpacket),
      .ff_tx_err   (tse_mac_transmit_error),
      .ff_tx_mod   (tse_mac_transmit_empty),
      .ff_tx_rdy   (tse_mac_transmit_ready),
      .ff_tx_sop   (tse_mac_transmit_startofpacket),
      .ff_tx_wren  (tse_mac_transmit_valid),
      .mdc         (mdc_from_the_tse_mac),
      .mdio_in     (mdio_in_to_the_tse_mac),
      .mdio_oen    (mdio_oen_from_the_tse_mac),
      .mdio_out    (mdio_out_from_the_tse_mac),
      .read        (tse_mac_control_port_read),
      .readdata    (tse_mac_control_port_readdata),
      .reset       (tse_mac_control_port_reset),
      .rgmii_in    (rgmii_in_to_the_tse_mac),
      .rgmii_out   (rgmii_out_from_the_tse_mac),
      .rx_clk      (rx_clk_to_the_tse_mac),
      .rx_control  (rx_control_to_the_tse_mac),
      .rx_err      (tse_mac_receive_error),
      .set_10      (set_10_to_the_tse_mac),
      .set_1000    (set_1000_to_the_tse_mac),
      .tx_clk      (tx_clk_to_the_tse_mac),
      .tx_control  (tx_control_from_the_tse_mac),
      .waitrequest (tse_mac_control_port_waitrequest),
      .write       (tse_mac_control_port_write),
      .writedata   (tse_mac_control_port_writedata)
    );

  tse_pll_s1_arbitrator the_tse_pll_s1
    (
      .clk                                                                            (clk_to_tse_pll),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave             (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_address_to_slave),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1           (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_granted_tse_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_nativeaddress                (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_nativeaddress),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1 (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_qualified_request_tse_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read                         (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_data_valid_tse_pll_s1   (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_read_data_valid_tse_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1          (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_requests_tse_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write                        (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_write),
      .cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata                    (cycloneIII_3c120_niosII_standard_sopc_clock_1_out_writedata),
      .d1_tse_pll_s1_end_xfer                                                         (d1_tse_pll_s1_end_xfer),
      .reset_n                                                                        (clk_to_tse_pll_reset_n),
      .tse_pll_s1_address                                                             (tse_pll_s1_address),
      .tse_pll_s1_chipselect                                                          (tse_pll_s1_chipselect),
      .tse_pll_s1_read                                                                (tse_pll_s1_read),
      .tse_pll_s1_readdata                                                            (tse_pll_s1_readdata),
      .tse_pll_s1_readdata_from_sa                                                    (tse_pll_s1_readdata_from_sa),
      .tse_pll_s1_reset_n                                                             (tse_pll_s1_reset_n),
      .tse_pll_s1_resetrequest                                                        (tse_pll_s1_resetrequest),
      .tse_pll_s1_resetrequest_from_sa                                                (tse_pll_s1_resetrequest_from_sa),
      .tse_pll_s1_write                                                               (tse_pll_s1_write),
      .tse_pll_s1_writedata                                                           (tse_pll_s1_writedata)
    );

  //tse_pll_c0_out out_clk assignment, which is an e_assign
  assign tse_pll_c0_out = out_clk_tse_pll_c0;

  tse_pll the_tse_pll
    (
      .address      (tse_pll_s1_address),
      .c0           (out_clk_tse_pll_c0),
      .chipselect   (tse_pll_s1_chipselect),
      .clk          (clk_to_tse_pll),
      .locked       (locked_from_the_tse_pll),
      .read         (tse_pll_s1_read),
      .readdata     (tse_pll_s1_readdata),
      .reset_n      (tse_pll_s1_reset_n),
      .resetrequest (tse_pll_s1_resetrequest),
      .write        (tse_pll_s1_write),
      .writedata    (tse_pll_s1_writedata)
    );

  tse_tx_pll_s1_arbitrator the_tse_tx_pll_s1
    (
      .clk                                                                               (clk),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave                (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_address_to_slave),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1           (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_granted_tse_tx_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_nativeaddress                   (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_nativeaddress),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1 (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_qualified_request_tse_tx_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read                            (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_data_valid_tse_tx_pll_s1   (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_read_data_valid_tse_tx_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1          (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_requests_tse_tx_pll_s1),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write                           (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_write),
      .cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata                       (cycloneIII_3c120_niosII_standard_sopc_clock_2_out_writedata),
      .d1_tse_tx_pll_s1_end_xfer                                                         (d1_tse_tx_pll_s1_end_xfer),
      .reset_n                                                                           (clk_reset_n),
      .tse_tx_pll_s1_address                                                             (tse_tx_pll_s1_address),
      .tse_tx_pll_s1_chipselect                                                          (tse_tx_pll_s1_chipselect),
      .tse_tx_pll_s1_read                                                                (tse_tx_pll_s1_read),
      .tse_tx_pll_s1_readdata                                                            (tse_tx_pll_s1_readdata),
      .tse_tx_pll_s1_readdata_from_sa                                                    (tse_tx_pll_s1_readdata_from_sa),
      .tse_tx_pll_s1_reset_n                                                             (tse_tx_pll_s1_reset_n),
      .tse_tx_pll_s1_resetrequest                                                        (tse_tx_pll_s1_resetrequest),
      .tse_tx_pll_s1_resetrequest_from_sa                                                (tse_tx_pll_s1_resetrequest_from_sa),
      .tse_tx_pll_s1_write                                                               (tse_tx_pll_s1_write),
      .tse_tx_pll_s1_writedata                                                           (tse_tx_pll_s1_writedata)
    );

  //tse_tx_pll_c0_out out_clk assignment, which is an e_assign
  assign tse_tx_pll_c0_out = out_clk_tse_tx_pll_c0;

  //tse_tx_pll_c1_out out_clk assignment, which is an e_assign
  assign tse_tx_pll_c1_out = out_clk_tse_tx_pll_c1;

  //tse_tx_pll_c2_out out_clk assignment, which is an e_assign
  assign tse_tx_pll_c2_out = out_clk_tse_tx_pll_c2;

  //tse_tx_pll_c3_out out_clk assignment, which is an e_assign
  assign tse_tx_pll_c3_out = out_clk_tse_tx_pll_c3;

  tse_tx_pll the_tse_tx_pll
    (
      .address      (tse_tx_pll_s1_address),
      .c0           (out_clk_tse_tx_pll_c0),
      .c1           (out_clk_tse_tx_pll_c1),
      .c2           (out_clk_tse_tx_pll_c2),
      .c3           (out_clk_tse_tx_pll_c3),
      .chipselect   (tse_tx_pll_s1_chipselect),
      .clk          (clk),
      .locked       (locked_from_the_tse_tx_pll),
      .read         (tse_tx_pll_s1_read),
      .readdata     (tse_tx_pll_s1_readdata),
      .reset_n      (tse_tx_pll_s1_reset_n),
      .resetrequest (tse_tx_pll_s1_resetrequest),
      .write        (tse_tx_pll_s1_write),
      .writedata    (tse_tx_pll_s1_writedata)
    );

  //reset is asserted asynchronously and deasserted synchronously
  cycloneIII_3c120_niosII_standard_sopc_reset_pll_c2_out_domain_synch_module cycloneIII_3c120_niosII_standard_sopc_reset_pll_c2_out_domain_synch
    (
      .clk      (pll_c2_out),
      .data_in  (1'b1),
      .data_out (pll_c2_out_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  cycloneIII_3c120_niosII_standard_sopc_reset_pll_c0_out_domain_synch_module cycloneIII_3c120_niosII_standard_sopc_reset_pll_c0_out_domain_synch
    (
      .clk      (pll_c0_out),
      .data_in  (1'b1),
      .data_out (pll_c0_out_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  cycloneIII_3c120_niosII_standard_sopc_reset_ddr2_sdram_phy_clk_out_domain_synch_module cycloneIII_3c120_niosII_standard_sopc_reset_ddr2_sdram_phy_clk_out_domain_synch
    (
      .clk      (ddr2_sdram_phy_clk_out),
      .data_in  (1'b1),
      .data_out (ddr2_sdram_phy_clk_out_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  cycloneIII_3c120_niosII_standard_sopc_reset_clk_domain_synch_module cycloneIII_3c120_niosII_standard_sopc_reset_clk_domain_synch
    (
      .clk      (clk),
      .data_in  (1'b1),
      .data_out (clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  cycloneIII_3c120_niosII_standard_sopc_reset_clk_to_tse_pll_domain_synch_module cycloneIII_3c120_niosII_standard_sopc_reset_clk_to_tse_pll_domain_synch
    (
      .clk      (clk_to_tse_pll),
      .data_in  (1'b1),
      .data_out (clk_to_tse_pll_reset_n),
      .reset_n  (reset_n_sources)
    );

  //cpu_ddr_clock_bridge_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign cpu_ddr_clock_bridge_m1_endofpacket = 0;

  //cycloneIII_3c120_niosII_standard_sopc_clock_0_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign cycloneIII_3c120_niosII_standard_sopc_clock_0_out_endofpacket = 0;

  //cycloneIII_3c120_niosII_standard_sopc_clock_1_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign cycloneIII_3c120_niosII_standard_sopc_clock_1_out_endofpacket = 0;

  //cycloneIII_3c120_niosII_standard_sopc_clock_2_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign cycloneIII_3c120_niosII_standard_sopc_clock_2_out_endofpacket = 0;

  //pipeline_bridge_before_tristate_bridge_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign pipeline_bridge_before_tristate_bridge_m1_endofpacket = 0;

  //sysid_control_slave_clock of type clock does not connect to anything so wire it to default (0)
  assign sysid_control_slave_clock = 0;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_lane0_module (
                                // inputs:
                                 data,
                                 rdaddress,
                                 rdclken,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 24: 0] rdaddress;
  input            rdclken;
  input   [ 24: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [33554431: 0];
  wire    [  7: 0] q;
  reg     [ 24: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_flash_lane0.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_flash_lane0.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 25,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash_lane1_module (
                                // inputs:
                                 data,
                                 rdaddress,
                                 rdclken,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 24: 0] rdaddress;
  input            rdclken;
  input   [ 24: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [33554431: 0];
  wire    [  7: 0] q;
  reg     [ 24: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_flash_lane1.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_flash_lane1.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 25,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_flash (
                   // inputs:
                    address,
                    read_n,
                    select_n,
                    write_n,

                   // outputs:
                    data
                 )
;

  inout   [ 15: 0] data;
  input   [ 24: 0] address;
  input            read_n;
  input            select_n;
  input            write_n;

  wire    [ 15: 0] data;
  wire    [  7: 0] data_0;
  wire    [  7: 0] data_1;
  wire    [ 15: 0] logic_vector_gasket;
  wire    [  7: 0] q_0;
  wire    [  7: 0] q_1;
  //s1, which is an e_ptf_slave

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign logic_vector_gasket = data;
  assign data_0 = logic_vector_gasket[7 : 0];
  //ext_flash_lane0, which is an e_ram
  ext_flash_lane0_module ext_flash_lane0
    (
      .data      (data_0),
      .q         (q_0),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data_1 = logic_vector_gasket[15 : 8];
  //ext_flash_lane1, which is an e_ram
  ext_flash_lane1_module ext_flash_lane1
    (
      .data      (data_1),
      .q         (q_1),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data = (~select_n & ~read_n)? {q_1,
    q_0}: {16{1'bz}};


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


//synthesis translate_off



// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE

// AND HERE WILL BE PRESERVED </ALTERA_NOTE>


// If user logic components use Altsync_Ram with convert_hex2ver.dll,
// set USE_convert_hex2ver in the user comments section above

// `ifdef USE_convert_hex2ver
// `else
// `define NO_PLI 1
// `endif

`include "c:/altera/11.0/quartus/eda/sim_lib/altera_mf.v"
`include "c:/altera/11.0/quartus/eda/sim_lib/220model.v"
`include "c:/altera/11.0/quartus/eda/sim_lib/sgate.v"
`include "C:/altera/11.0/quartus/eda/sim_lib/stratixiigx_hssi_atoms.v"
`include "C:/altera/11.0/quartus/eda/sim_lib/stratixiv_hssi_atoms.v"
`include "tse_mac.vo"
`include "tse_mac_loopback.v"
`include "descriptor_memory.v"
`include "pll.v"
`include "altpllpll.v"
`include "sysid.v"
`include "pipeline_bridge_before_tristate_bridge.v"
`include "button_pio.v"
`include "cycloneIII_3c120_niosII_standard_sopc_clock_1.v"
`include "high_res_timer.v"
`include "tse_tx_pll.v"
`include "altplltse_tx_pll.v"
`include "cycloneIII_3c120_niosII_standard_sopc_clock_2.v"
`include "led_pio.v"
`include "jtag_uart.v"
`include "tse_pll.v"
`include "altplltse_pll.v"
`include "sgdma_rx.v"
`include "sys_clk_timer.v"
`include "performance_counter.v"
`include "cpu_test_bench.v"
`include "cpu_mult_cell.v"
`include "cpu_oci_test_bench.v"
`include "cpu_jtag_debug_module_tck.v"
`include "cpu_jtag_debug_module_sysclk.v"
`include "cpu_jtag_debug_module_wrapper.v"
`include "cpu.v"
`include "slow_peripheral_bridge.v"
`include "cpu_ddr_clock_bridge.v"
`include "sgdma_tx.v"
`include "cycloneIII_3c120_niosII_standard_sopc_clock_0.v"

`timescale 1ns / 1ps

module test_bench 
;


  reg              clk;
  reg              clk_125;
  reg              clk_to_tse_pll;
  wire             cpu_ddr_clock_bridge_m1_endofpacket;
  wire    [ 23: 0] cpu_ddr_clock_bridge_m1_nativeaddress;
  wire             cpu_ddr_clock_bridge_s1_endofpacket_from_sa;
  wire             cs_n_to_the_max2;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_0_out_endofpacket;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_1_out_endofpacket;
  wire             cycloneIII_3c120_niosII_standard_sopc_clock_2_out_endofpacket;
  wire             ddr2_sdram_aux_full_rate_clk_out;
  wire             ddr2_sdram_aux_half_rate_clk_out;
  wire             ddr2_sdram_phy_clk_out;
  wire             ena_10_from_the_tse_mac;
  wire             eth_mode_from_the_tse_mac;
  wire    [ 25: 0] flash_tristate_bridge_address;
  wire    [ 31: 0] flash_tristate_bridge_data;
  wire             global_reset_n_to_the_ddr2_sdram;
  wire    [  3: 0] in_port_to_the_button_pio;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             local_init_done_from_the_ddr2_sdram;
  wire             local_refresh_ack_from_the_ddr2_sdram;
  wire             local_wdata_req_from_the_ddr2_sdram;
  wire             locked_from_the_pll;
  wire             locked_from_the_tse_pll;
  wire             locked_from_the_tse_tx_pll;
  wire             mdc_from_the_tse_mac;
  wire             mdio_in_to_the_tse_mac;
  wire             mdio_oen_from_the_tse_mac;
  wire             mdio_out_from_the_tse_mac;
  wire    [ 12: 0] mem_addr_from_the_ddr2_sdram;
  wire    [  1: 0] mem_ba_from_the_ddr2_sdram;
  wire             mem_cas_n_from_the_ddr2_sdram;
  wire             mem_cke_from_the_ddr2_sdram;
  wire             mem_clk_n_to_and_from_the_ddr2_sdram;
  wire             mem_clk_to_and_from_the_ddr2_sdram;
  wire             mem_cs_n_from_the_ddr2_sdram;
  wire    [  1: 0] mem_dm_from_the_ddr2_sdram;
  wire    [ 15: 0] mem_dq_to_and_from_the_ddr2_sdram;
  wire    [  1: 0] mem_dqs_to_and_from_the_ddr2_sdram;
  wire             mem_odt_from_the_ddr2_sdram;
  wire             mem_ras_n_from_the_ddr2_sdram;
  wire             mem_we_n_from_the_ddr2_sdram;
  wire             oe_n_to_the_max2;
  wire    [  7: 0] out_port_from_the_led_pio;
  wire             pipeline_bridge_before_tristate_bridge_m1_debugaccess;
  wire             pipeline_bridge_before_tristate_bridge_m1_endofpacket;
  wire             pipeline_bridge_before_tristate_bridge_s1_endofpacket_from_sa;
  wire             pll_c0_out;
  wire             pll_c2_out;
  wire             pll_c3_out;
  wire             pll_c4_out;
  wire             read_n_to_the_ext_flash;
  reg              reset_n;
  wire             reset_phy_clk_n_from_the_ddr2_sdram;
  wire    [  3: 0] rgmii_in_to_the_tse_mac;
  wire    [  3: 0] rgmii_out_from_the_tse_mac;
  wire             rx_clk_to_the_tse_mac;
  wire             rx_control_to_the_tse_mac;
  wire             select_n_to_the_ext_flash;
  wire             set_1000_to_the_tse_mac;
  wire             set_10_to_the_tse_mac;
  wire             slow_peripheral_bridge_s1_endofpacket_from_sa;
  wire             sysid_control_slave_clock;
  wire             tse_pll_c0_out;
  wire             tse_tx_pll_c0_out;
  wire             tse_tx_pll_c1_out;
  wire             tse_tx_pll_c2_out;
  wire             tse_tx_pll_c3_out;
  wire             tx_clk_to_the_tse_mac;
  wire             tx_control_from_the_tse_mac;
  wire             we_n_to_the_max2;
  wire             write_n_to_the_ext_flash;


// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
//  add your signals and additional architecture here
// AND HERE WILL BE PRESERVED </ALTERA_NOTE>

  //Set us up the Dut
  cycloneIII_3c120_niosII_standard_sopc DUT
    (
      .clk                                   (clk),
      .clk_125                               (clk_125),
      .clk_to_tse_pll                        (clk_to_tse_pll),
      .cs_n_to_the_max2                      (cs_n_to_the_max2),
      .ddr2_sdram_aux_full_rate_clk_out      (ddr2_sdram_aux_full_rate_clk_out),
      .ddr2_sdram_aux_half_rate_clk_out      (ddr2_sdram_aux_half_rate_clk_out),
      .ddr2_sdram_phy_clk_out                (ddr2_sdram_phy_clk_out),
      .ena_10_from_the_tse_mac               (ena_10_from_the_tse_mac),
      .eth_mode_from_the_tse_mac             (eth_mode_from_the_tse_mac),
      .flash_tristate_bridge_address         (flash_tristate_bridge_address),
      .flash_tristate_bridge_data            (flash_tristate_bridge_data),
      .global_reset_n_to_the_ddr2_sdram      (global_reset_n_to_the_ddr2_sdram),
      .in_port_to_the_button_pio             (in_port_to_the_button_pio),
      .local_init_done_from_the_ddr2_sdram   (local_init_done_from_the_ddr2_sdram),
      .local_refresh_ack_from_the_ddr2_sdram (local_refresh_ack_from_the_ddr2_sdram),
      .local_wdata_req_from_the_ddr2_sdram   (local_wdata_req_from_the_ddr2_sdram),
      .locked_from_the_pll                   (locked_from_the_pll),
      .locked_from_the_tse_pll               (locked_from_the_tse_pll),
      .locked_from_the_tse_tx_pll            (locked_from_the_tse_tx_pll),
      .mdc_from_the_tse_mac                  (mdc_from_the_tse_mac),
      .mdio_in_to_the_tse_mac                (mdio_in_to_the_tse_mac),
      .mdio_oen_from_the_tse_mac             (mdio_oen_from_the_tse_mac),
      .mdio_out_from_the_tse_mac             (mdio_out_from_the_tse_mac),
      .mem_addr_from_the_ddr2_sdram          (mem_addr_from_the_ddr2_sdram),
      .mem_ba_from_the_ddr2_sdram            (mem_ba_from_the_ddr2_sdram),
      .mem_cas_n_from_the_ddr2_sdram         (mem_cas_n_from_the_ddr2_sdram),
      .mem_cke_from_the_ddr2_sdram           (mem_cke_from_the_ddr2_sdram),
      .mem_clk_n_to_and_from_the_ddr2_sdram  (mem_clk_n_to_and_from_the_ddr2_sdram),
      .mem_clk_to_and_from_the_ddr2_sdram    (mem_clk_to_and_from_the_ddr2_sdram),
      .mem_cs_n_from_the_ddr2_sdram          (mem_cs_n_from_the_ddr2_sdram),
      .mem_dm_from_the_ddr2_sdram            (mem_dm_from_the_ddr2_sdram),
      .mem_dq_to_and_from_the_ddr2_sdram     (mem_dq_to_and_from_the_ddr2_sdram),
      .mem_dqs_to_and_from_the_ddr2_sdram    (mem_dqs_to_and_from_the_ddr2_sdram),
      .mem_odt_from_the_ddr2_sdram           (mem_odt_from_the_ddr2_sdram),
      .mem_ras_n_from_the_ddr2_sdram         (mem_ras_n_from_the_ddr2_sdram),
      .mem_we_n_from_the_ddr2_sdram          (mem_we_n_from_the_ddr2_sdram),
      .oe_n_to_the_max2                      (oe_n_to_the_max2),
      .out_port_from_the_led_pio             (out_port_from_the_led_pio),
      .pll_c0_out                            (pll_c0_out),
      .pll_c2_out                            (pll_c2_out),
      .pll_c3_out                            (pll_c3_out),
      .pll_c4_out                            (pll_c4_out),
      .read_n_to_the_ext_flash               (read_n_to_the_ext_flash),
      .reset_n                               (reset_n),
      .reset_phy_clk_n_from_the_ddr2_sdram   (reset_phy_clk_n_from_the_ddr2_sdram),
      .rgmii_in_to_the_tse_mac               (rgmii_in_to_the_tse_mac),
      .rgmii_out_from_the_tse_mac            (rgmii_out_from_the_tse_mac),
      .rx_clk_to_the_tse_mac                 (rx_clk_to_the_tse_mac),
      .rx_control_to_the_tse_mac             (rx_control_to_the_tse_mac),
      .select_n_to_the_ext_flash             (select_n_to_the_ext_flash),
      .set_1000_to_the_tse_mac               (set_1000_to_the_tse_mac),
      .set_10_to_the_tse_mac                 (set_10_to_the_tse_mac),
      .tse_pll_c0_out                        (tse_pll_c0_out),
      .tse_tx_pll_c0_out                     (tse_tx_pll_c0_out),
      .tse_tx_pll_c1_out                     (tse_tx_pll_c1_out),
      .tse_tx_pll_c2_out                     (tse_tx_pll_c2_out),
      .tse_tx_pll_c3_out                     (tse_tx_pll_c3_out),
      .tx_clk_to_the_tse_mac                 (tx_clk_to_the_tse_mac),
      .tx_control_from_the_tse_mac           (tx_control_from_the_tse_mac),
      .we_n_to_the_max2                      (we_n_to_the_max2),
      .write_n_to_the_ext_flash              (write_n_to_the_ext_flash)
    );

  //default value specified in MODULE button_pio ptf port section
  assign in_port_to_the_button_pio = 15;

  ext_flash the_ext_flash
    (
      .address  (flash_tristate_bridge_address[25 : 1]),
      .data     (flash_tristate_bridge_data),
      .read_n   (read_n_to_the_ext_flash),
      .select_n (select_n_to_the_ext_flash),
      .write_n  (write_n_to_the_ext_flash)
    );

  tse_mac_loopback the_tse_mac_loopback
    (
      .rgmii_in   (rgmii_in_to_the_tse_mac),
      .rgmii_out  (rgmii_out_from_the_tse_mac),
      .rx_clk     (rx_clk_to_the_tse_mac),
      .rx_control (rx_control_to_the_tse_mac),
      .set_10     (set_10_to_the_tse_mac),
      .set_1000   (set_1000_to_the_tse_mac),
      .tx_clk     (tx_clk_to_the_tse_mac),
      .tx_control (tx_control_from_the_tse_mac)
    );

  initial
    clk = 1'b0;
  always
    #10 clk <= ~clk;
  
  initial
    clk_125 = 1'b0;
  always
    #4 clk_125 <= ~clk_125;
  
  initial
    clk_to_tse_pll = 1'b0;
  always
    #4 clk_to_tse_pll <= ~clk_to_tse_pll;
  
  initial 
    begin
      reset_n <= 0;
      #200 reset_n <= 1;
    end

endmodule


//synthesis translate_on